netcdf PRVI_DOV18 {
types:
  compound ggxfParameterType {
    char parameterName(32) ;
    char parameterSet(32) ;
    char unit(16) ;
    double unitSiRatio ;
    int sourceCrsAxis ;
    float parameterMinimumValue ;
    float parameterMaximumValue ;
    float noDataFlag ;
  }; // ggxfParameterType

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "d2018prvi.gxt" ;
		:content = "deviationsOfTheVertical" ;
		:title = "hybrid defelection of the vertical model" ;
		:summary = "hybrid defelection of the vertical model" ;
		:geospatial_lat_min = 17.67 ;
		:geospatial_lon_min = -65.09 ;
		:geospatial_lat_max = 18.42 ;
		:geospatial_lon_max = -64.6 ;
		:extent_description = "US Puerto Rico and Virgin Islands - onshore." ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		ggxfParameterType :parameters = 
    {{"deviationEast"}, {"deviation"}, {"arc-second"}, 4.84813681109536e-06, -1, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"deviationNorth"}, {"deviation"}, {"arc-second"}, 4.84813681109536e-60, -1, -3.402823e+38, -3.402823e+38, -3.402823e+38} ;
		:organisationName = "National Geodetic Survey, National Oceanic and Atmospheric Administration." ;
		:deliveryPoint = "1315 East West Hwy" ;
		:city = "Silver Spring" ;
		:postalCode = "20910" ;
		:country = "United States of America" ;
		:publisher_url = "https://geodesy.noaa.gov/PC_PROD/GEOID18/Format_ascii/g2018p0.asc.zip" ;

group: Puerto\ Rico\ Virgin\ Islands\ DEFLEC18 {
  dimensions:
  	deviationCount = 2 ;

  // group attributes:
  		:interpolationMethod = "biquadratic" ;

  group: Puerto\ Rico\ Virgin\ Islands\ DEFLEC18 {
    dimensions:
    	iNodeCount = 301 ;
    	jNodeCount = 361 ;
    variables:
    	float deviation(jNodeCount, iNodeCount, deviationCount) ;

    // group attributes:
    		:affineCoeffs = 15., 0., 0.01666666667, -69., 0.01666666667, 0. ;
    		:gridPriority = 1LL ;
    } // group Puerto\ Rico\ Virgin\ Islands\ DEFLEC18
  } // group Puerto\ Rico\ Virgin\ Islands\ DEFLEC18
}

netcdf PRGEOID18c {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "g2018pr.yaml" ;
		:content = "geoidModel" ;
		:title = "hybrid geoid" ;
		:summary = "hybrid geoid" ;
		:geospatial_lat_min = 17.87 ;
		:geospatial_lon_min = -68. ;
		:geospatial_lat_max = 18.53 ;
		:geospatial_lon_max = -65. ;
		:extent_description = "Puerto Rico - onshore." ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,3],\n  AXIS[\"Geodetic latitude (Lat)\",north,\n    ANGLEUNIT[\"degree\",0.0174532925199433]],\n  AXIS[\"Geodetic longitude (Lon)\",east,\n    ANGLEUNIT[\"degree\",0.0174532925199433]],\n  AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1]]]\n" ;
		:targetCrsWkt = "VERTCRS[\"PRVD02 - NOHt\",\n  VDATUM[\"Puerto Rico Vertical Datum of 2002\"],\n  CS[vertical,1],\n  AXIS[\"Gravity-related height (H)\",up],\n  LENGTHUNIT[\"metre\",1]]\n" ;
		:parameters.count = 1LL ;
		:parameters.1.parameterName = "geoidHeight" ;
		:parameters.1.sourceCrsAxis = 2LL ;
		:parameters.1.unit = "metre" ;
		:parameters.1.unitSiRatio = 1. ;
		:operationAccuracy = 0.015 ;
		:organisationName = "National Geodetic Survey, National Oceanic and Atmospheric Administration." ;
		:deliveryPoint = "1315 East West Hwy" ;
		:city = "Silver Spring" ;
		:postalCode = "20910" ;
		:country = "United States of America" ;
		:publisher_url = "https://geodesy.noaa.gov/PC_PROD/GEOID18/Format_ascii/g2018p0.asc.zip" ;

group: puerto_rico_virgin_islands_geoid18 {

  // group attributes:
  		:interpolationMethod = "biquadratic" ;

  group: puerto_rico_virgin_islands_geoid18 {
    dimensions:
    	iNodeCount = 301 ;
    	jNodeCount = 361 ;
    variables:
    	float geoidHeight(jNodeCount, iNodeCount) ;

    // group attributes:
    		:affineCoeffs = 21., 0., -0.01666666667, -69., 0.01666666667, 0. ;
    		:comment = "grid starts in the top left (northwest) corner and works across (east) and down (south)" ;
    data:

     geoidHeight =
  -48.78305, -48.80028, -48.81684, -48.83206, -48.84526, -48.85678, 
        -48.8663, -48.87355, -48.87912, -48.88332, -48.88619, -48.8886, 
        -48.89069, -48.89234, -48.8933, -48.89377, -48.89314, -48.89293, 
        -48.89263, -48.89187, -48.89218, -48.89224, -48.89166, -48.89031, 
        -48.88785, -48.88445, -48.87976, -48.87428, -48.8683, -48.8624, 
        -48.85727, -48.85369, -48.85246, -48.8542, -48.85839, -48.86666, 
        -48.87736, -48.88977, -48.90282, -48.91617, -48.92979, -48.94383, 
        -48.95836, -48.97329, -48.98832, -49.00299, -49.01662, -49.02858, 
        -49.03848, -49.04697, -49.05259, -49.05816, -49.0629, -49.06755, 
        -49.0728, -49.07906, -49.08646, -49.09483, -49.10374, -49.11247, 
        -49.12014, -49.12598, -49.12951, -49.13059, -49.12936, -49.12572, 
        -49.11972, -49.11039, -49.10004, -49.08797, -49.07435, -49.05917, 
        -49.04245, -49.02449, -49.00586, -48.98722, -48.96898, -48.95147, 
        -48.9355, -48.92112, -48.90885, -48.89822, -48.88929, -48.88166, 
        -48.8752, -48.86848, -48.86397, -48.86023, -48.85715, -48.85422, 
        -48.85096, -48.84689, -48.84162, -48.83519, -48.82781, -48.82008, 
        -48.81266, -48.80618, -48.80106, -48.79741, -48.79522, -48.79436, 
        -48.79462, -48.79565, -48.79618, -48.79775, -48.79959, -48.80183, 
        -48.80435, -48.80719, -48.80995, -48.81234, -48.81442, -48.81581, 
        -48.81649, -48.81704, -48.81771, -48.81913, -48.82182, -48.82645, 
        -48.83329, -48.8423, -48.85308, -48.86507, -48.87691, -48.89041, 
        -48.90491, -48.92072, -48.93817, -48.95758, -48.97898, -49.00218, 
        -49.02662, -49.05164, -49.07644, -49.10026, -49.12251, -49.14288, 
        -49.16155, -49.17851, -49.19406, -49.20859, -49.22262, -49.23671, 
        -49.25122, -49.26623, -49.28062, -49.2963, -49.31214, -49.32834, 
        -49.34475, -49.36176, -49.37925, -49.39748, -49.41659, -49.43653, 
        -49.45695, -49.47782, -49.49889, -49.51989, -49.54026, -49.55966, 
        -49.57775, -49.59444, -49.60984, -49.62416, -49.63751, -49.65052, 
        -49.66362, -49.67723, -49.69053, -49.70543, -49.72072, -49.73625, 
        -49.75179, -49.76764, -49.78382, -49.80025, -49.81658, -49.83237, 
        -49.84721, -49.86093, -49.87365, -49.88571, -49.89745, -49.90913, 
        -49.92103, -49.93313, -49.94541, -49.9577, -49.96944, -49.98053, 
        -49.99062, -49.99987, -50.00855, -50.01697, -50.02434, -50.03257, 
        -50.04026, -50.04681, -50.05156, -50.05442, -50.05544, -50.05462, 
        -50.05232, -50.04877, -50.04428, -50.03931, -50.03451, -50.03054, 
        -50.02788, -50.02668, -50.02661, -50.02711, -50.0277, -50.02825, 
        -50.02891, -50.02987, -50.03114, -50.03238, -50.03306, -50.03278, 
        -50.03132, -50.02867, -50.02502, -50.02042, -50.01402, -50.00789, 
        -50.00097, -49.99334, -49.98492, -49.9757, -49.96562, -49.95469, 
        -49.94291, -49.92999, -49.9157, -49.90018, -49.88324, -49.86501, 
        -49.84572, -49.82573, -49.80561, -49.78568, -49.76615, -49.74718, 
        -49.72844, -49.70995, -49.69128, -49.67216, -49.65249, -49.63237, 
        -49.61212, -49.59184, -49.57157, -49.5512, -49.53095, -49.51102, 
        -49.4917, -49.47322, -49.45572, -49.43917, -49.42215, -49.40631, 
        -49.39045, -49.37476, -49.35954, -49.34506, -49.33139, -49.31843, 
        -49.30597, -49.29389, -49.28235, -49.271, -49.25978, -49.24877, 
        -49.23803, -49.22762, -49.21756, -49.20774, -49.19803, -49.1884, 
        -49.17902, -49.17006, -49.16156, -49.15365, -49.14629, -49.13941, 
        -49.13327, -49.12705, -49.12057, -49.11403, -49.10689, -49.09922, 
        -49.09119, -49.08274, -49.07359, -49.06397, -49.05436, -49.04467, 
        -49.0349,
  -48.77826, -48.7972, -48.81584, -48.83282, -48.84852, -48.86188, 
        -48.87299, -48.88194, -48.88895, -48.89429, -48.89832, -48.90161, 
        -48.90447, -48.90558, -48.90684, -48.9073, -48.90725, -48.90718, 
        -48.9072, -48.90772, -48.90806, -48.90825, -48.90792, -48.90695, 
        -48.90519, -48.90242, -48.89851, -48.89352, -48.88675, -48.88072, 
        -48.87512, -48.87073, -48.86853, -48.86912, -48.87296, -48.87985, 
        -48.88933, -48.90055, -48.91275, -48.92563, -48.93908, -48.95332, 
        -48.96848, -48.98429, -48.99942, -49.01521, -49.0298, -49.0425, 
        -49.05298, -49.0612, -49.06752, -49.07245, -49.07655, -49.08053, 
        -49.08506, -49.09067, -49.0975, -49.10551, -49.11434, -49.12339, 
        -49.13187, -49.13797, -49.14322, -49.14639, -49.14732, -49.14598, 
        -49.14218, -49.13591, -49.12749, -49.11721, -49.10534, -49.09181, 
        -49.0767, -49.06021, -49.04321, -49.02615, -49.0093, -48.99311, 
        -48.97797, -48.96328, -48.95122, -48.94062, -48.9318, -48.92413, 
        -48.91755, -48.91194, -48.90766, -48.90468, -48.90239, -48.90055, 
        -48.89879, -48.89631, -48.8927, -48.88785, -48.88208, -48.87584, 
        -48.86987, -48.86377, -48.85978, -48.85689, -48.85512, -48.85429, 
        -48.85399, -48.85427, -48.85487, -48.85551, -48.85638, -48.85754, 
        -48.85899, -48.86065, -48.86223, -48.86342, -48.86429, -48.86451, 
        -48.86436, -48.86405, -48.86407, -48.86397, -48.86632, -48.87069, 
        -48.87716, -48.88597, -48.89672, -48.90891, -48.92208, -48.9361, 
        -48.95102, -48.96719, -48.98489, -49.00462, -49.02645, -49.04998, 
        -49.07475, -49.10016, -49.12541, -49.14962, -49.17221, -49.19302, 
        -49.21099, -49.22835, -49.24408, -49.25874, -49.27266, -49.28642, 
        -49.30035, -49.31454, -49.32909, -49.34408, -49.35919, -49.37477, 
        -49.39087, -49.40763, -49.42527, -49.44406, -49.46407, -49.48512, 
        -49.50681, -49.52883, -49.55084, -49.57249, -49.59332, -49.61171, 
        -49.62936, -49.6453, -49.65972, -49.67294, -49.68539, -49.69756, 
        -49.71017, -49.72351, -49.73784, -49.75312, -49.76914, -49.78571, 
        -49.80264, -49.82008, -49.8378, -49.85561, -49.8731, -49.88974, 
        -49.90501, -49.9188, -49.93132, -49.94309, -49.95443, -49.96596, 
        -49.97686, -49.98917, -50.00189, -50.0145, -50.02696, -50.03865, 
        -50.04947, -50.05938, -50.06858, -50.07735, -50.0859, -50.09419, 
        -50.10185, -50.10829, -50.11286, -50.11543, -50.11604, -50.11508, 
        -50.11273, -50.10921, -50.10465, -50.09953, -50.09442, -50.08997, 
        -50.08666, -50.08459, -50.08336, -50.08237, -50.08017, -50.07876, 
        -50.07744, -50.07655, -50.07623, -50.07617, -50.07599, -50.0752, 
        -50.07354, -50.07093, -50.06736, -50.0629, -50.05733, -50.05082, 
        -50.04326, -50.03475, -50.02532, -50.01507, -50.00407, -49.99237, 
        -49.97981, -49.96645, -49.95189, -49.9365, -49.91981, -49.90236, 
        -49.88407, -49.8652, -49.84607, -49.82691, -49.80781, -49.78882, 
        -49.76983, -49.75075, -49.73023, -49.71069, -49.69061, -49.67023, 
        -49.64968, -49.62918, -49.60841, -49.58744, -49.56649, -49.54588, 
        -49.52594, -49.50678, -49.48864, -49.47144, -49.45462, -49.43809, 
        -49.42158, -49.4054, -49.38937, -49.37421, -49.3599, -49.34614, 
        -49.33283, -49.31975, -49.30689, -49.29419, -49.28167, -49.26945, 
        -49.25773, -49.24656, -49.23599, -49.22588, -49.21599, -49.20626, 
        -49.19674, -49.18761, -49.17883, -49.17044, -49.16244, -49.15519, 
        -49.14848, -49.14202, -49.13586, -49.12834, -49.12151, -49.11411, 
        -49.10621, -49.09772, -49.08901, -49.07997, -49.07088, -49.06176, 
        -49.05282,
  -48.77236, -48.79402, -48.8148, -48.83398, -48.85109, -48.86627, 
        -48.87902, -48.88942, -48.89714, -48.90392, -48.90926, -48.91355, 
        -48.91695, -48.91962, -48.92113, -48.92162, -48.92207, -48.92239, 
        -48.92291, -48.92326, -48.92371, -48.92381, -48.92379, -48.92237, 
        -48.92139, -48.91961, -48.91669, -48.91251, -48.90743, -48.90181, 
        -48.89633, -48.89176, -48.88905, -48.88884, -48.89157, -48.89722, 
        -48.9054, -48.91544, -48.92569, -48.93801, -48.95114, -48.96519, 
        -48.98057, -48.99686, -49.01374, -49.03039, -49.0458, -49.05911, 
        -49.06993, -49.0783, -49.08465, -49.08939, -49.09317, -49.09668, 
        -49.10055, -49.10437, -49.11037, -49.1176, -49.12583, -49.13462, 
        -49.14331, -49.1512, -49.15773, -49.16254, -49.16536, -49.16607, 
        -49.16428, -49.15996, -49.15335, -49.14481, -49.13451, -49.12283, 
        -49.10859, -49.09405, -49.0788, -49.06348, -49.04843, -49.03366, 
        -49.01942, -49.00657, -48.99503, -48.98468, -48.97539, -48.96777, 
        -48.96106, -48.95547, -48.95108, -48.94837, -48.94726, -48.9467, 
        -48.94522, -48.94455, -48.94279, -48.93979, -48.93579, -48.93138, 
        -48.92691, -48.92306, -48.92018, -48.91814, -48.91672, -48.91582, 
        -48.91517, -48.9149, -48.91491, -48.91505, -48.91535, -48.91585, 
        -48.91653, -48.91628, -48.9169, -48.91722, -48.91716, -48.91677, 
        -48.91603, -48.91521, -48.91478, -48.91522, -48.91711, -48.92104, 
        -48.92698, -48.93499, -48.94514, -48.95696, -48.97007, -48.98417, 
        -48.99934, -49.01571, -49.03365, -49.05398, -49.07522, -49.09925, 
        -49.12453, -49.15047, -49.17626, -49.20098, -49.22412, -49.2452, 
        -49.26453, -49.28213, -49.29833, -49.31339, -49.32753, -49.34106, 
        -49.35455, -49.36825, -49.3821, -49.39621, -49.41077, -49.42587, 
        -49.44165, -49.45838, -49.47529, -49.49474, -49.51571, -49.53794, 
        -49.56077, -49.58372, -49.60645, -49.62849, -49.6493, -49.66844, 
        -49.68544, -49.70037, -49.71369, -49.72586, -49.73751, -49.74918, 
        -49.76144, -49.77467, -49.78907, -49.80472, -49.82144, -49.83907, 
        -49.85742, -49.87632, -49.89454, -49.9137, -49.93224, -49.9497, 
        -49.9654, -49.9793, -49.9916, -50.00299, -50.01414, -50.0256, 
        -50.03759, -50.05014, -50.06312, -50.07632, -50.08925, -50.10168, 
        -50.11328, -50.12388, -50.13361, -50.14269, -50.15131, -50.15957, 
        -50.16706, -50.17327, -50.17768, -50.18011, -50.18076, -50.17895, 
        -50.17688, -50.17358, -50.16918, -50.16404, -50.15869, -50.15368, 
        -50.14961, -50.14648, -50.14386, -50.14109, -50.13794, -50.13449, 
        -50.13113, -50.12852, -50.1266, -50.12516, -50.12401, -50.12257, 
        -50.12063, -50.11802, -50.11457, -50.11011, -50.10427, -50.09703, 
        -50.08841, -50.07848, -50.06755, -50.05598, -50.0438, -50.03114, 
        -50.0179, -50.00291, -49.98807, -49.97245, -49.95623, -49.93941, 
        -49.92215, -49.9044, -49.88628, -49.86784, -49.84922, -49.83031, 
        -49.81115, -49.79163, -49.77148, -49.75154, -49.73144, -49.71111, 
        -49.69081, -49.67026, -49.64932, -49.62798, -49.60654, -49.58538, 
        -49.56491, -49.54506, -49.52626, -49.50857, -49.49107, -49.47405, 
        -49.45658, -49.4395, -49.4229, -49.40659, -49.39109, -49.37617, 
        -49.36161, -49.3471, -49.3329, -49.31794, -49.30408, -49.29082, 
        -49.27812, -49.26623, -49.25503, -49.24443, -49.23428, -49.22457, 
        -49.21501, -49.20575, -49.19655, -49.1876, -49.17905, -49.17113, 
        -49.16394, -49.15726, -49.15074, -49.14418, -49.13734, -49.13017, 
        -49.12251, -49.11443, -49.10603, -49.09743, -49.08895, -49.08057, 
        -49.07239,
  -48.76383, -48.78888, -48.81146, -48.83309, -48.85238, -48.86917, 
        -48.88346, -48.89572, -48.90581, -48.914, -48.92066, -48.92598, 
        -48.93024, -48.93346, -48.9355, -48.9365, -48.93698, -48.9363, 
        -48.93664, -48.93692, -48.93712, -48.93737, -48.93761, -48.93785, 
        -48.93791, -48.93748, -48.9358, -48.93277, -48.92872, -48.92393, 
        -48.91916, -48.91495, -48.91216, -48.91052, -48.91246, -48.91706, 
        -48.92408, -48.93304, -48.94341, -48.95507, -48.96764, -48.98152, 
        -48.99661, -49.0128, -49.02995, -49.04691, -49.06269, -49.07641, 
        -49.08759, -49.09558, -49.10239, -49.10751, -49.11141, -49.11485, 
        -49.11835, -49.12249, -49.12764, -49.13388, -49.14119, -49.1493, 
        -49.15769, -49.16583, -49.17306, -49.17895, -49.18317, -49.18543, 
        -49.18435, -49.18177, -49.17678, -49.16981, -49.16123, -49.15119, 
        -49.14019, -49.12801, -49.11507, -49.10198, -49.08882, -49.07574, 
        -49.06298, -49.05088, -49.0397, -49.02954, -49.02026, -49.0113, 
        -49.0044, -48.99863, -48.99451, -48.99196, -48.99134, -48.9918, 
        -48.99287, -48.99369, -48.99389, -48.9928, -48.99065, -48.98796, 
        -48.98504, -48.98244, -48.98056, -48.97929, -48.97824, -48.97745, 
        -48.97572, -48.97528, -48.97512, -48.97519, -48.97537, -48.97562, 
        -48.97586, -48.97599, -48.97598, -48.97575, -48.97531, -48.97459, 
        -48.9736, -48.97256, -48.97194, -48.9721, -48.97333, -48.97628, 
        -48.98116, -48.98821, -48.9962, -49.00717, -49.01977, -49.03374, 
        -49.04895, -49.06573, -49.08406, -49.10488, -49.12767, -49.15265, 
        -49.17873, -49.20538, -49.23183, -49.25713, -49.2805, -49.30204, 
        -49.32167, -49.33955, -49.35623, -49.37179, -49.38625, -49.39901, 
        -49.41226, -49.42532, -49.43858, -49.45203, -49.46598, -49.48067, 
        -49.4963, -49.51318, -49.53164, -49.55191, -49.57387, -49.59711, 
        -49.62082, -49.64443, -49.66749, -49.6896, -49.71024, -49.72868, 
        -49.74477, -49.75883, -49.77111, -49.78246, -49.79358, -49.80405, 
        -49.81628, -49.82964, -49.84434, -49.86042, -49.87771, -49.89621, 
        -49.91569, -49.93585, -49.95632, -49.97661, -49.99616, -50.0142, 
        -50.03031, -50.04438, -50.05635, -50.0675, -50.07849, -50.08986, 
        -50.10198, -50.11479, -50.12812, -50.14174, -50.15533, -50.16853, 
        -50.18093, -50.19128, -50.20156, -50.21085, -50.21948, -50.22749, 
        -50.23459, -50.24063, -50.24495, -50.24747, -50.24829, -50.24796, 
        -50.24637, -50.24342, -50.23915, -50.23395, -50.22835, -50.22293, 
        -50.21809, -50.21371, -50.20939, -50.20469, -50.19946, -50.19408, 
        -50.18899, -50.18467, -50.18131, -50.1787, -50.17639, -50.17427, 
        -50.17098, -50.1682, -50.16468, -50.15999, -50.15367, -50.14557, 
        -50.13533, -50.12364, -50.11086, -50.09761, -50.08404, -50.07032, 
        -50.05626, -50.04162, -50.02632, -50.01049, -49.99443, -49.97824, 
        -49.96185, -49.9451, -49.92792, -49.91026, -49.89206, -49.87331, 
        -49.85429, -49.83481, -49.81477, -49.79453, -49.77439, -49.75442, 
        -49.73436, -49.71399, -49.69305, -49.67152, -49.64972, -49.62813, 
        -49.60592, -49.58553, -49.56607, -49.54759, -49.52958, -49.51167, 
        -49.49406, -49.47607, -49.45839, -49.44105, -49.42429, -49.40775, 
        -49.39163, -49.37566, -49.36007, -49.34468, -49.32962, -49.31536, 
        -49.3018, -49.28907, -49.27712, -49.26598, -49.25549, -49.24553, 
        -49.23592, -49.22651, -49.21719, -49.20768, -49.19851, -49.18996, 
        -49.18216, -49.17501, -49.16825, -49.1616, -49.15482, -49.14777, 
        -49.14033, -49.13254, -49.12451, -49.11631, -49.10815, -49.1002, 
        -49.09243,
  -48.75083, -48.78029, -48.80751, -48.83214, -48.85392, -48.87258, 
        -48.88865, -48.90238, -48.91411, -48.92357, -48.93143, -48.93764, 
        -48.94176, -48.94564, -48.94822, -48.94942, -48.9499, -48.94999, 
        -48.94999, -48.94994, -48.95, -48.95036, -48.95112, -48.95214, 
        -48.95338, -48.95431, -48.95407, -48.95162, -48.949, -48.94554, 
        -48.94173, -48.9383, -48.93586, -48.93518, -48.93671, -48.94062, 
        -48.94682, -48.95499, -48.96474, -48.97572, -48.98775, -49.00109, 
        -49.01577, -49.03067, -49.04716, -49.06382, -49.07939, -49.09322, 
        -49.10485, -49.11457, -49.12229, -49.1284, -49.13302, -49.13687, 
        -49.14047, -49.14427, -49.1487, -49.15396, -49.16015, -49.16638, 
        -49.17413, -49.18189, -49.18924, -49.19556, -49.20053, -49.20377, 
        -49.20486, -49.20354, -49.19988, -49.19432, -49.18742, -49.17948, 
        -49.17054, -49.16098, -49.15071, -49.14006, -49.12918, -49.11713, 
        -49.1061, -49.09524, -49.08478, -49.07495, -49.06586, -49.05765, 
        -49.05048, -49.0446, -49.04039, -49.03804, -49.0376, -49.03854, 
        -49.04097, -49.0433, -49.04499, -49.04547, -49.0451, -49.04298, 
        -49.04158, -49.0403, -49.03924, -49.0386, -49.03818, -49.03783, 
        -49.03746, -49.03733, -49.0374, -49.03777, -49.03826, -49.0385, 
        -49.0386, -49.03846, -49.03818, -49.03782, -49.03738, -49.03682, 
        -49.03485, -49.03376, -49.03294, -49.0327, -49.03347, -49.03524, 
        -49.03872, -49.0442, -49.05188, -49.06169, -49.0735, -49.08725, 
        -49.10266, -49.1199, -49.1391, -49.16074, -49.18448, -49.21003, 
        -49.237, -49.26444, -49.29152, -49.31636, -49.34, -49.36168, 
        -49.38152, -49.39984, -49.41692, -49.43299, -49.44791, -49.46178, 
        -49.47494, -49.48758, -49.5003, -49.51318, -49.52673, -49.54123, 
        -49.55704, -49.57434, -49.5935, -49.61467, -49.63759, -49.66158, 
        -49.68586, -49.70978, -49.73181, -49.75356, -49.77353, -49.79116, 
        -49.8064, -49.81946, -49.83101, -49.8419, -49.85286, -49.86451, 
        -49.87707, -49.89091, -49.90625, -49.92268, -49.94057, -49.95974, 
        -49.98002, -50.0011, -50.02253, -50.04369, -50.06395, -50.08245, 
        -50.09874, -50.11267, -50.12459, -50.1345, -50.14541, -50.15697, 
        -50.16925, -50.18235, -50.19606, -50.21015, -50.22435, -50.23832, 
        -50.25151, -50.26354, -50.27427, -50.28373, -50.29222, -50.29997, 
        -50.30684, -50.31257, -50.31694, -50.3198, -50.3212, -50.32138, 
        -50.32006, -50.3172, -50.31298, -50.3077, -50.30189, -50.29594, 
        -50.2903, -50.28351, -50.27734, -50.27064, -50.26346, -50.25628, 
        -50.24963, -50.24371, -50.23926, -50.23576, -50.23257, -50.22974, 
        -50.22679, -50.2235, -50.21956, -50.21432, -50.20718, -50.19775, 
        -50.186, -50.17241, -50.15772, -50.14256, -50.12728, -50.11245, 
        -50.09745, -50.08208, -50.06628, -50.05022, -50.03423, -50.01845, 
        -50.00277, -49.98679, -49.97038, -49.95335, -49.9347, -49.91643, 
        -49.89767, -49.87843, -49.85878, -49.83889, -49.81907, -49.79922, 
        -49.7793, -49.75904, -49.73812, -49.71642, -49.69427, -49.67208, 
        -49.65039, -49.62946, -49.60946, -49.59027, -49.57161, -49.55329, 
        -49.53499, -49.51651, -49.49794, -49.47942, -49.46112, -49.44308, 
        -49.42525, -49.40772, -49.39054, -49.37387, -49.3578, -49.34235, 
        -49.32801, -49.31455, -49.30187, -49.29001, -49.27913, -49.26888, 
        -49.25907, -49.24943, -49.23978, -49.22903, -49.21933, -49.2103, 
        -49.20185, -49.19423, -49.18716, -49.18046, -49.17354, -49.16649, 
        -49.15923, -49.15171, -49.14401, -49.13589, -49.12788, -49.1201, 
        -49.11286,
  -48.73574, -48.77024, -48.80169, -48.82994, -48.85466, -48.87559, 
        -48.8925, -48.90791, -48.92101, -48.93192, -48.9407, -48.94792, 
        -48.95388, -48.95839, -48.96107, -48.96264, -48.96298, -48.96255, 
        -48.96202, -48.96156, -48.96146, -48.961, -48.9623, -48.96437, 
        -48.96696, -48.96909, -48.97049, -48.9708, -48.96976, -48.96789, 
        -48.96542, -48.96298, -48.96123, -48.96087, -48.96244, -48.9662, 
        -48.9721, -48.97884, -48.98811, -48.99864, -49.01031, -49.02326, 
        -49.03735, -49.0524, -49.06802, -49.08342, -49.09825, -49.11187, 
        -49.12407, -49.1348, -49.14368, -49.15091, -49.15672, -49.16049, 
        -49.16462, -49.16854, -49.17262, -49.17713, -49.18238, -49.18845, 
        -49.19529, -49.20226, -49.20913, -49.21515, -49.22011, -49.22362, 
        -49.22517, -49.2246, -49.22197, -49.21771, -49.21143, -49.20546, 
        -49.19909, -49.19218, -49.18472, -49.1768, -49.16855, -49.16, 
        -49.15122, -49.14215, -49.13259, -49.12329, -49.11443, -49.10625, 
        -49.09904, -49.09313, -49.08885, -49.08647, -49.08512, -49.08649, 
        -49.08934, -49.09233, -49.09525, -49.09719, -49.0981, -49.0984, 
        -49.09827, -49.09802, -49.09793, -49.09813, -49.0985, -49.09898, 
        -49.09946, -49.10008, -49.10073, -49.1016, -49.10251, -49.10212, 
        -49.10233, -49.10225, -49.10206, -49.10196, -49.10188, -49.10162, 
        -49.10096, -49.10008, -49.09924, -49.09856, -49.09845, -49.09925, 
        -49.10122, -49.10512, -49.11129, -49.11989, -49.13105, -49.14452, 
        -49.16022, -49.17713, -49.1973, -49.21991, -49.24466, -49.27117, 
        -49.29884, -49.32697, -49.35453, -49.38064, -49.40461, -49.42646, 
        -49.44648, -49.4651, -49.4825, -49.49905, -49.51436, -49.52849, 
        -49.54147, -49.5539, -49.56624, -49.57898, -49.59226, -49.60596, 
        -49.62209, -49.64008, -49.66012, -49.68217, -49.70581, -49.7303, 
        -49.75482, -49.77867, -49.80124, -49.82222, -49.84118, -49.85779, 
        -49.87211, -49.88445, -49.89559, -49.9064, -49.91766, -49.92983, 
        -49.9431, -49.95759, -49.97349, -49.99075, -50.00914, -50.0279, 
        -50.04864, -50.07029, -50.09236, -50.11407, -50.13473, -50.15348, 
        -50.16977, -50.18359, -50.19552, -50.20654, -50.21761, -50.22934, 
        -50.24198, -50.25543, -50.2696, -50.2841, -50.29887, -50.31345, 
        -50.32727, -50.33983, -50.35089, -50.3604, -50.36872, -50.37612, 
        -50.38278, -50.38838, -50.39201, -50.39535, -50.3973, -50.39777, 
        -50.3966, -50.39373, -50.38939, -50.38386, -50.37761, -50.37112, 
        -50.36421, -50.35703, -50.34915, -50.34065, -50.33182, -50.32313, 
        -50.31528, -50.30854, -50.30314, -50.29862, -50.29467, -50.29093, 
        -50.28714, -50.28299, -50.27807, -50.27188, -50.26362, -50.2528, 
        -50.23949, -50.22417, -50.20766, -50.18974, -50.17292, -50.1567, 
        -50.14062, -50.12446, -50.10815, -50.09188, -50.07589, -50.06031, 
        -50.04493, -50.0294, -50.01345, -49.99695, -49.97968, -49.96184, 
        -49.94353, -49.92481, -49.90573, -49.88639, -49.86702, -49.84738, 
        -49.8276, -49.80704, -49.78579, -49.76379, -49.74129, -49.71874, 
        -49.69667, -49.67533, -49.65486, -49.63516, -49.61608, -49.59726, 
        -49.57844, -49.5594, -49.54007, -49.52061, -49.50087, -49.48024, 
        -49.46078, -49.44149, -49.42279, -49.4049, -49.38786, -49.37147, 
        -49.35618, -49.34196, -49.32867, -49.31621, -49.30475, -49.29393, 
        -49.28368, -49.2737, -49.26362, -49.25354, -49.24361, -49.23413, 
        -49.22533, -49.21728, -49.20987, -49.20302, -49.19621, -49.18879, 
        -49.18149, -49.174, -49.16634, -49.15828, -49.15029, -49.14257, 
        -49.13534,
  -48.71621, -48.75557, -48.79247, -48.82492, -48.85335, -48.87735, 
        -48.89738, -48.91454, -48.92908, -48.94116, -48.95101, -48.9591, 
        -48.9654, -48.97024, -48.97351, -48.9749, -48.97417, -48.9734, 
        -48.97226, -48.97146, -48.97133, -48.97232, -48.97416, -48.97715, 
        -48.98086, -48.98422, -48.98708, -48.98905, -48.98979, -48.98957, 
        -48.98866, -48.98645, -48.98558, -48.98586, -48.98788, -48.99195, 
        -48.998, -49.00574, -49.01496, -49.0253, -49.03686, -49.04947, 
        -49.06293, -49.07702, -49.09135, -49.10556, -49.11934, -49.1313, 
        -49.14389, -49.15522, -49.16515, -49.17371, -49.18089, -49.18694, 
        -49.19211, -49.19667, -49.20089, -49.2051, -49.20959, -49.21474, 
        -49.22049, -49.22638, -49.23227, -49.23735, -49.24068, -49.24361, 
        -49.24487, -49.24457, -49.2426, -49.23944, -49.23566, -49.23171, 
        -49.22773, -49.22353, -49.21903, -49.21412, -49.20886, -49.20319, 
        -49.19691, -49.18999, -49.18209, -49.17253, -49.16418, -49.15636, 
        -49.14945, -49.14382, -49.13956, -49.1372, -49.13677, -49.13811, 
        -49.14077, -49.14399, -49.14706, -49.14991, -49.15199, -49.15339, 
        -49.15444, -49.15522, -49.15606, -49.1572, -49.15762, -49.15929, 
        -49.16095, -49.16257, -49.1642, -49.16573, -49.16714, -49.16817, 
        -49.16875, -49.16897, -49.16919, -49.16957, -49.17007, -49.17039, 
        -49.17028, -49.16972, -49.16889, -49.16784, -49.16704, -49.16674, 
        -49.16652, -49.16906, -49.17394, -49.18149, -49.19208, -49.20543, 
        -49.22159, -49.24029, -49.26147, -49.28506, -49.31074, -49.33806, 
        -49.36637, -49.39486, -49.42274, -49.44901, -49.47318, -49.4952, 
        -49.51537, -49.53436, -49.55223, -49.56809, -49.58378, -49.59819, 
        -49.61139, -49.62367, -49.63594, -49.64846, -49.66193, -49.67687, 
        -49.69355, -49.71248, -49.73348, -49.75632, -49.78048, -49.80515, 
        -49.82954, -49.85282, -49.8746, -49.8944, -49.91209, -49.92751, 
        -49.94101, -49.95287, -49.96304, -49.97423, -49.98614, -49.99916, 
        -50.01339, -50.02877, -50.04542, -50.06326, -50.08226, -50.10229, 
        -50.12341, -50.14538, -50.16778, -50.18981, -50.21061, -50.22931, 
        -50.24548, -50.2593, -50.27147, -50.28289, -50.29438, -50.30654, 
        -50.31965, -50.33348, -50.34819, -50.36316, -50.37738, -50.39237, 
        -50.40657, -50.41938, -50.43049, -50.43998, -50.44809, -50.4553, 
        -50.46175, -50.46746, -50.47235, -50.47612, -50.47843, -50.479, 
        -50.47776, -50.47475, -50.47017, -50.46424, -50.4574, -50.4499, 
        -50.44186, -50.4332, -50.42375, -50.41392, -50.40392, -50.39428, 
        -50.38561, -50.37803, -50.37165, -50.36527, -50.3605, -50.35585, 
        -50.351, -50.34563, -50.33939, -50.33179, -50.32208, -50.30984, 
        -50.29525, -50.2785, -50.26052, -50.24215, -50.22395, -50.20628, 
        -50.18909, -50.17211, -50.15533, -50.1388, -50.12272, -50.10723, 
        -50.09177, -50.07613, -50.06015, -50.0438, -50.02685, -50.00931, 
        -49.99146, -49.97334, -49.95488, -49.93619, -49.917, -49.89725, 
        -49.87719, -49.8564, -49.83373, -49.81131, -49.78844, -49.76575, 
        -49.74349, -49.72192, -49.70116, -49.68105, -49.66138, -49.64211, 
        -49.62291, -49.60345, -49.58354, -49.56316, -49.54234, -49.52139, 
        -49.50048, -49.47982, -49.45973, -49.44039, -49.4221, -49.40501, 
        -49.38886, -49.37363, -49.35978, -49.3469, -49.3348, -49.32342, 
        -49.31249, -49.30181, -49.29112, -49.28076, -49.27052, -49.26071, 
        -49.25152, -49.24316, -49.23524, -49.22788, -49.22077, -49.2133, 
        -49.20593, -49.19823, -49.19028, -49.18225, -49.17426, -49.16552, 
        -49.15826,
  -48.694, -48.74025, -48.78254, -48.82038, -48.85283, -48.8799, 
        -48.90248, -48.92153, -48.93739, -48.95059, -48.96041, -48.96906, 
        -48.97598, -48.98117, -48.98441, -48.98604, -48.98603, -48.98497, 
        -48.98337, -48.98268, -48.98254, -48.98399, -48.98651, -48.99035, 
        -48.99489, -48.99828, -49.00232, -49.00574, -49.00822, -49.00969, 
        -49.01031, -49.01038, -49.01058, -49.0118, -49.01456, -49.01931, 
        -49.026, -49.03422, -49.04367, -49.05421, -49.06576, -49.07713, 
        -49.09004, -49.10311, -49.11608, -49.1289, -49.14147, -49.15396, 
        -49.16626, -49.17799, -49.18881, -49.19844, -49.20692, -49.21438, 
        -49.22091, -49.22661, -49.23164, -49.23522, -49.23952, -49.24401, 
        -49.24866, -49.25332, -49.25784, -49.26171, -49.26464, -49.26652, 
        -49.26692, -49.26626, -49.26464, -49.26227, -49.25976, -49.25756, 
        -49.25581, -49.25432, -49.25282, -49.25008, -49.24809, -49.24567, 
        -49.24227, -49.23752, -49.23134, -49.22413, -49.21656, -49.20963, 
        -49.20351, -49.19854, -49.19477, -49.19264, -49.19199, -49.19291, 
        -49.19482, -49.19741, -49.20041, -49.20231, -49.20509, -49.20754, 
        -49.20962, -49.21144, -49.21328, -49.21547, -49.21818, -49.2212, 
        -49.22424, -49.22713, -49.22976, -49.23215, -49.23415, -49.23568, 
        -49.23671, -49.23744, -49.23827, -49.23935, -49.23959, -49.24066, 
        -49.2412, -49.24103, -49.24024, -49.23903, -49.23769, -49.23669, 
        -49.23664, -49.23827, -49.24224, -49.24917, -49.25927, -49.27274, 
        -49.28947, -49.30892, -49.33108, -49.35557, -49.38197, -49.40977, 
        -49.43837, -49.46598, -49.4938, -49.52007, -49.54435, -49.56665, 
        -49.58736, -49.60664, -49.62488, -49.64223, -49.65836, -49.67313, 
        -49.68662, -49.69917, -49.71126, -49.72385, -49.73761, -49.75314, 
        -49.77077, -49.7906, -49.81252, -49.83596, -49.8603, -49.88375, 
        -49.90759, -49.93006, -49.95063, -49.9691, -49.98543, -49.99979, 
        -50.01256, -50.02434, -50.03587, -50.04783, -50.06072, -50.07485, 
        -50.09014, -50.10654, -50.12397, -50.14239, -50.16175, -50.18208, 
        -50.20341, -50.22555, -50.24804, -50.27005, -50.29069, -50.30908, 
        -50.32411, -50.33807, -50.35065, -50.36264, -50.37475, -50.38746, 
        -50.40107, -50.41555, -50.43082, -50.44645, -50.46205, -50.47714, 
        -50.49132, -50.504, -50.51498, -50.52434, -50.53235, -50.5394, 
        -50.54581, -50.55167, -50.55678, -50.56086, -50.56323, -50.56368, 
        -50.56219, -50.55892, -50.55399, -50.54774, -50.53924, -50.5306, 
        -50.52134, -50.51134, -50.50076, -50.48987, -50.47916, -50.46889, 
        -50.45938, -50.45091, -50.4437, -50.43746, -50.43177, -50.42623, 
        -50.42021, -50.41345, -50.40566, -50.39646, -50.38521, -50.37176, 
        -50.35568, -50.33789, -50.31899, -50.29961, -50.28025, -50.26125, 
        -50.24282, -50.22498, -50.20775, -50.19093, -50.17454, -50.15855, 
        -50.14155, -50.12548, -50.10918, -50.09262, -50.0757, -50.05845, 
        -50.04083, -50.02331, -50.00528, -49.98655, -49.96772, -49.94788, 
        -49.92739, -49.90591, -49.88357, -49.86064, -49.83757, -49.81483, 
        -49.79266, -49.77119, -49.75025, -49.72979, -49.70964, -49.68987, 
        -49.67044, -49.65051, -49.63008, -49.60909, -49.58751, -49.56553, 
        -49.5435, -49.52161, -49.50027, -49.47969, -49.46013, -49.44183, 
        -49.4247, -49.4091, -49.3947, -49.38132, -49.36767, -49.35562, 
        -49.34389, -49.33241, -49.32124, -49.31009, -49.29937, -49.28907, 
        -49.27938, -49.27039, -49.2621, -49.25438, -49.24671, -49.23886, 
        -49.23103, -49.22296, -49.21478, -49.2066, -49.19848, -49.19068, 
        -49.18333,
  -48.6722, -48.72416, -48.77217, -48.81497, -48.8519, -48.88167, 
        -48.90704, -48.92806, -48.94542, -48.96, -48.97165, -48.98077, 
        -48.98791, -48.99332, -48.99657, -48.99791, -48.99764, -48.99636, 
        -48.99503, -48.99417, -48.99338, -48.99503, -48.99837, -49.00309, 
        -49.00839, -49.01358, -49.01872, -49.02338, -49.02727, -49.03019, 
        -49.03224, -49.03369, -49.0352, -49.03748, -49.0414, -49.04622, 
        -49.05381, -49.06276, -49.07275, -49.0836, -49.0952, -49.10732, 
        -49.1197, -49.13192, -49.14382, -49.15543, -49.16701, -49.17871, 
        -49.19054, -49.20223, -49.21342, -49.22282, -49.23242, -49.24116, 
        -49.24928, -49.25655, -49.26296, -49.26854, -49.27338, -49.27773, 
        -49.28173, -49.28528, -49.28841, -49.29067, -49.29187, -49.29214, 
        -49.29144, -49.29002, -49.28714, -49.28519, -49.28369, -49.28294, 
        -49.28313, -49.28405, -49.28531, -49.28661, -49.2877, -49.28839, 
        -49.28761, -49.28511, -49.28093, -49.27545, -49.26947, -49.26382, 
        -49.259, -49.25519, -49.25147, -49.24995, -49.24913, -49.24955, 
        -49.25063, -49.25229, -49.25466, -49.25743, -49.26039, -49.26354, 
        -49.26651, -49.26936, -49.27235, -49.27577, -49.27973, -49.28403, 
        -49.28844, -49.29257, -49.29629, -49.29856, -49.3013, -49.30352, 
        -49.30522, -49.30667, -49.30824, -49.31003, -49.31207, -49.31394, 
        -49.31522, -49.31565, -49.3153, -49.3143, -49.31281, -49.31148, 
        -49.31126, -49.3126, -49.31613, -49.32259, -49.33254, -49.34519, 
        -49.36221, -49.38233, -49.40524, -49.43037, -49.45724, -49.4853, 
        -49.51389, -49.5423, -49.56988, -49.59602, -49.62036, -49.64286, 
        -49.66402, -49.68393, -49.7029, -49.72076, -49.73742, -49.7527, 
        -49.76663, -49.77952, -49.79202, -49.80394, -49.81812, -49.83421, 
        -49.8525, -49.87304, -49.89561, -49.91921, -49.94355, -49.96775, 
        -49.99073, -50.01213, -50.03152, -50.0488, -50.06408, -50.07765, 
        -50.09001, -50.10181, -50.11377, -50.12653, -50.14046, -50.15572, 
        -50.17221, -50.18968, -50.20798, -50.22606, -50.24585, -50.26647, 
        -50.28787, -50.31007, -50.3324, -50.35416, -50.37443, -50.39248, 
        -50.40854, -50.42262, -50.43547, -50.44805, -50.46074, -50.47406, 
        -50.48828, -50.50333, -50.5192, -50.53526, -50.55109, -50.56623, 
        -50.58013, -50.59249, -50.60315, -50.61228, -50.6201, -50.62609, 
        -50.63255, -50.63856, -50.64397, -50.64799, -50.65023, -50.65047, 
        -50.64866, -50.64497, -50.63972, -50.6329, -50.62467, -50.61525, 
        -50.60493, -50.59393, -50.58253, -50.57107, -50.55986, -50.54905, 
        -50.53885, -50.52959, -50.52134, -50.51398, -50.50745, -50.50079, 
        -50.49357, -50.48545, -50.47622, -50.46552, -50.45291, -50.43712, 
        -50.42011, -50.40168, -50.38208, -50.36193, -50.34162, -50.32148, 
        -50.30201, -50.28328, -50.2652, -50.2477, -50.23063, -50.21377, 
        -50.19697, -50.18005, -50.16298, -50.14586, -50.12861, -50.11124, 
        -50.09375, -50.07611, -50.05812, -50.03959, -50.02038, -50.00028, 
        -49.97922, -49.95717, -49.93436, -49.91112, -49.88797, -49.86531, 
        -49.84331, -49.82203, -49.80111, -49.7804, -49.76005, -49.73981, 
        -49.71896, -49.6988, -49.67798, -49.65646, -49.63431, -49.61169, 
        -49.58884, -49.566, -49.5435, -49.52183, -49.50109, -49.48167, 
        -49.46384, -49.44758, -49.43277, -49.41905, -49.40606, -49.39352, 
        -49.38112, -49.36879, -49.35659, -49.34464, -49.33297, -49.32186, 
        -49.31133, -49.30157, -49.29259, -49.28412, -49.2758, -49.26739, 
        -49.25885, -49.25015, -49.24152, -49.233, -49.22466, -49.21672, 
        -49.20923,
  -48.65121, -48.70842, -48.76182, -48.80944, -48.85052, -48.88491, 
        -48.91314, -48.93649, -48.95575, -48.97151, -48.984, -48.99383, 
        -49.00123, -49.00642, -49.00846, -49.00958, -49.0092, -49.00794, 
        -49.00658, -49.00584, -49.0064, -49.00867, -49.01262, -49.01786, 
        -49.02372, -49.02974, -49.03564, -49.0412, -49.04615, -49.04931, 
        -49.05267, -49.05546, -49.05828, -49.06191, -49.0671, -49.07415, 
        -49.08286, -49.09277, -49.10347, -49.11477, -49.12655, -49.13861, 
        -49.15061, -49.16223, -49.17331, -49.18296, -49.19354, -49.20435, 
        -49.21551, -49.22683, -49.23801, -49.24883, -49.25919, -49.26911, 
        -49.27863, -49.28762, -49.29586, -49.3031, -49.30917, -49.31406, 
        -49.31786, -49.32061, -49.32137, -49.32203, -49.32158, -49.32013, 
        -49.31794, -49.31546, -49.31308, -49.31121, -49.31028, -49.31063, 
        -49.3124, -49.31534, -49.31901, -49.32299, -49.32686, -49.3301, 
        -49.33202, -49.33104, -49.32906, -49.32556, -49.32144, -49.31758, 
        -49.31451, -49.31235, -49.31095, -49.31007, -49.30951, -49.30928, 
        -49.30944, -49.31018, -49.31172, -49.31409, -49.3172, -49.3208, 
        -49.32462, -49.32856, -49.33178, -49.33642, -49.34158, -49.34708, 
        -49.35259, -49.35783, -49.36258, -49.36679, -49.37043, -49.37347, 
        -49.37602, -49.37831, -49.38069, -49.38336, -49.38624, -49.38898, 
        -49.39116, -49.39249, -49.39289, -49.39245, -49.39049, -49.38959, 
        -49.38946, -49.39084, -49.39444, -49.40098, -49.41095, -49.42462, 
        -49.44192, -49.46254, -49.48599, -49.51162, -49.53873, -49.56671, 
        -49.5949, -49.62275, -49.64972, -49.67542, -49.69964, -49.72243, 
        -49.74407, -49.76373, -49.78345, -49.80207, -49.81937, -49.83522, 
        -49.84972, -49.8632, -49.87628, -49.88977, -49.90455, -49.92126, 
        -49.9402, -49.9613, -49.98409, -50.00792, -50.03202, -50.05557, 
        -50.0778, -50.0982, -50.11656, -50.13289, -50.14743, -50.16054, 
        -50.17176, -50.18375, -50.19622, -50.20973, -50.22465, -50.24101, 
        -50.25864, -50.27726, -50.29659, -50.31647, -50.33681, -50.3577, 
        -50.37918, -50.40116, -50.42319, -50.44448, -50.46426, -50.482, 
        -50.49773, -50.51189, -50.5251, -50.53802, -50.5512, -50.56508, 
        -50.57991, -50.59465, -50.611, -50.62742, -50.64337, -50.65833, 
        -50.67186, -50.68373, -50.69391, -50.70264, -50.71029, -50.71723, 
        -50.72374, -50.72986, -50.73522, -50.73919, -50.74121, -50.74108, 
        -50.73893, -50.73499, -50.72942, -50.72221, -50.71344, -50.70329, 
        -50.69213, -50.68036, -50.66835, -50.65644, -50.64481, -50.63351, 
        -50.62167, -50.6115, -50.60226, -50.59396, -50.58629, -50.5786, 
        -50.57032, -50.56104, -50.55051, -50.53848, -50.52465, -50.50885, 
        -50.49122, -50.47217, -50.4521, -50.43138, -50.41031, -50.38923, 
        -50.3686, -50.34871, -50.32964, -50.31124, -50.29325, -50.27537, 
        -50.25741, -50.23932, -50.22124, -50.20324, -50.18536, -50.16753, 
        -50.14965, -50.13161, -50.11322, -50.09329, -50.07359, -50.05289, 
        -50.03115, -50.00841, -49.98501, -49.96144, -49.93826, -49.91582, 
        -49.89418, -49.87315, -49.85238, -49.83167, -49.81109, -49.79071, 
        -49.77053, -49.75018, -49.72924, -49.70747, -49.68489, -49.66177, 
        -49.63835, -49.61488, -49.59161, -49.56888, -49.5471, -49.5267, 
        -49.50803, -49.49123, -49.47611, -49.46223, -49.44907, -49.43616, 
        -49.42321, -49.41011, -49.39695, -49.38388, -49.37109, -49.35881, 
        -49.34725, -49.33657, -49.32668, -49.31732, -49.3081, -49.29774, 
        -49.28821, -49.27861, -49.26913, -49.25994, -49.25117, -49.24288, 
        -49.23512,
  -48.63464, -48.69619, -48.75407, -48.80608, -48.85109, -48.88881, 
        -48.91992, -48.94566, -48.96579, -48.98306, -48.99672, -49.00712, 
        -49.01469, -49.01965, -49.02252, -49.02351, -49.02312, -49.02202, 
        -49.02083, -49.02032, -49.02118, -49.02385, -49.02828, -49.03399, 
        -49.03932, -49.04578, -49.05211, -49.05819, -49.06389, -49.06904, 
        -49.07357, -49.0777, -49.08192, -49.08698, -49.09355, -49.10191, 
        -49.11185, -49.12283, -49.1344, -49.14529, -49.15736, -49.16948, 
        -49.18134, -49.19265, -49.20326, -49.21329, -49.22308, -49.23302, 
        -49.24335, -49.25403, -49.26489, -49.27574, -49.28652, -49.29726, 
        -49.30804, -49.31871, -49.32795, -49.33727, -49.34512, -49.3512, 
        -49.35542, -49.35787, -49.35868, -49.35802, -49.35601, -49.35289, 
        -49.34914, -49.34539, -49.34223, -49.34013, -49.33947, -49.34052, 
        -49.34337, -49.3468, -49.35236, -49.35848, -49.36461, -49.37015, 
        -49.37442, -49.37684, -49.37722, -49.37602, -49.3741, -49.37236, 
        -49.3713, -49.37097, -49.37106, -49.37116, -49.37098, -49.37052, 
        -49.37003, -49.36893, -49.36973, -49.37169, -49.37481, -49.37884, 
        -49.38349, -49.38857, -49.39405, -49.39988, -49.40613, -49.41251, 
        -49.41884, -49.4249, -49.43053, -49.43563, -49.44016, -49.44415, 
        -49.44767, -49.45094, -49.45326, -49.45683, -49.46064, -49.46443, 
        -49.46779, -49.47038, -49.47198, -49.47263, -49.47262, -49.47255, 
        -49.47319, -49.47527, -49.47947, -49.4864, -49.49659, -49.51036, 
        -49.5278, -49.54866, -49.5724, -49.5983, -49.62547, -49.65214, 
        -49.67965, -49.70657, -49.73259, -49.75755, -49.78141, -49.80429, 
        -49.82638, -49.84775, -49.86827, -49.88768, -49.90569, -49.92224, 
        -49.93744, -49.95169, -49.9656, -49.97995, -49.99551, -50.01288, 
        -50.03236, -50.05383, -50.0768, -50.09958, -50.12338, -50.14636, 
        -50.16788, -50.18751, -50.20515, -50.22093, -50.23512, -50.24811, 
        -50.26042, -50.27271, -50.28563, -50.29977, -50.31548, -50.33281, 
        -50.35152, -50.37128, -50.39172, -50.41254, -50.43357, -50.45486, 
        -50.47643, -50.4982, -50.51978, -50.53948, -50.55862, -50.57581, 
        -50.59122, -50.6053, -50.61864, -50.63177, -50.64523, -50.65947, 
        -50.67473, -50.69092, -50.70765, -50.72435, -50.74032, -50.75503, 
        -50.76809, -50.77935, -50.78896, -50.79726, -50.80467, -50.81154, 
        -50.8181, -50.82428, -50.82962, -50.83344, -50.83516, -50.83468, 
        -50.83125, -50.82712, -50.8214, -50.814, -50.80483, -50.79412, 
        -50.78234, -50.76997, -50.75747, -50.74514, -50.7331, -50.72135, 
        -50.70991, -50.69897, -50.6888, -50.67947, -50.67074, -50.66207, 
        -50.65284, -50.64258, -50.63099, -50.61788, -50.6031, -50.58655, 
        -50.56837, -50.54886, -50.52833, -50.50704, -50.48523, -50.46324, 
        -50.44152, -50.42048, -50.39927, -50.37977, -50.36065, -50.34153, 
        -50.3222, -50.30274, -50.28336, -50.26425, -50.24543, -50.22676, 
        -50.20805, -50.18914, -50.16985, -50.15, -50.12939, -50.10782, 
        -50.08522, -50.06174, -50.03777, -50.01393, -49.99075, -49.96853, 
        -49.94724, -49.9265, -49.90594, -49.88536, -49.86481, -49.84445, 
        -49.82421, -49.80379, -49.78276, -49.76085, -49.7381, -49.71481, 
        -49.69118, -49.66735, -49.64351, -49.61998, -49.59729, -49.57504, 
        -49.55566, -49.53835, -49.52291, -49.50889, -49.49563, -49.48253, 
        -49.46918, -49.45543, -49.44133, -49.42713, -49.41312, -49.39964, 
        -49.38696, -49.37519, -49.36421, -49.35367, -49.34321, -49.33258, 
        -49.32175, -49.31092, -49.30034, -49.29019, -49.28065, -49.27182, 
        -49.26374,
  -48.62285, -48.68734, -48.74835, -48.80273, -48.85112, -48.89201, 
        -48.92604, -48.95414, -48.97756, -48.99635, -49.01124, -49.02217, 
        -49.0301, -49.03519, -49.03797, -49.03889, -49.03847, -49.03754, 
        -49.03553, -49.03524, -49.03639, -49.03938, -49.0442, -49.05026, 
        -49.05677, -49.06348, -49.07003, -49.07628, -49.08258, -49.08852, 
        -49.09406, -49.09952, -49.10525, -49.11073, -49.1187, -49.1284, 
        -49.13961, -49.15178, -49.16437, -49.17706, -49.18963, -49.20206, 
        -49.21399, -49.22517, -49.2356, -49.24534, -49.25461, -49.26384, 
        -49.27336, -49.2823, -49.29259, -49.30311, -49.31393, -49.32519, 
        -49.33695, -49.34914, -49.36132, -49.3728, -49.38275, -49.39047, 
        -49.39573, -49.39861, -49.39905, -49.39753, -49.39437, -49.38965, 
        -49.38338, -49.37831, -49.37423, -49.37167, -49.37098, -49.37234, 
        -49.37583, -49.38116, -49.38809, -49.39578, -49.40359, -49.41095, 
        -49.41724, -49.42188, -49.42467, -49.42596, -49.42644, -49.42694, 
        -49.42692, -49.42838, -49.42996, -49.43122, -49.43176, -49.43159, 
        -49.4311, -49.43067, -49.43103, -49.43276, -49.43589, -49.44035, 
        -49.44581, -49.45205, -49.45884, -49.46591, -49.47303, -49.48003, 
        -49.48681, -49.4923, -49.49845, -49.50419, -49.50939, -49.51424, 
        -49.51873, -49.52292, -49.52719, -49.53176, -49.53672, -49.54197, 
        -49.5469, -49.55123, -49.55464, -49.55698, -49.55851, -49.5598, 
        -49.56177, -49.56513, -49.57036, -49.57703, -49.58763, -49.60156, 
        -49.61901, -49.63985, -49.66361, -49.68951, -49.71649, -49.74368, 
        -49.77025, -49.79604, -49.82086, -49.84491, -49.86821, -49.89098, 
        -49.91334, -49.93525, -49.95643, -49.97651, -49.99527, -50.01245, 
        -50.02741, -50.04263, -50.05751, -50.07291, -50.08962, -50.10741, 
        -50.1273, -50.14902, -50.17211, -50.19587, -50.21944, -50.24199, 
        -50.26319, -50.28243, -50.29976, -50.31539, -50.32956, -50.34264, 
        -50.35518, -50.36782, -50.38121, -50.39592, -50.41236, -50.43055, 
        -50.44924, -50.46981, -50.49149, -50.51345, -50.53529, -50.55706, 
        -50.57874, -50.60024, -50.62123, -50.64121, -50.65962, -50.6762, 
        -50.69123, -50.70518, -50.71849, -50.73159, -50.74513, -50.7594, 
        -50.77489, -50.79102, -50.80791, -50.82488, -50.84074, -50.85509, 
        -50.8676, -50.87821, -50.88624, -50.89413, -50.90128, -50.90808, 
        -50.9146, -50.92083, -50.92622, -50.92999, -50.93157, -50.93094, 
        -50.92837, -50.92409, -50.91828, -50.91079, -50.90132, -50.89012, 
        -50.87791, -50.86506, -50.85208, -50.83933, -50.82692, -50.81477, 
        -50.80294, -50.79145, -50.78048, -50.77018, -50.7604, -50.75073, 
        -50.74058, -50.72956, -50.71596, -50.70203, -50.68652, -50.66949, 
        -50.65083, -50.63081, -50.60963, -50.58768, -50.56515, -50.54225, 
        -50.51955, -50.49746, -50.4761, -50.45543, -50.43517, -50.41468, 
        -50.39382, -50.37278, -50.35177, -50.3313, -50.31123, -50.29136, 
        -50.27147, -50.25124, -50.23053, -50.20922, -50.18723, -50.16443, 
        -50.14082, -50.11653, -50.09187, -50.06794, -50.04488, -50.02287, 
        -50.00189, -49.98143, -49.9601, -49.93972, -49.91957, -49.89945, 
        -49.8793, -49.85891, -49.83785, -49.81583, -49.79296, -49.76966, 
        -49.74603, -49.72205, -49.6979, -49.67383, -49.65054, -49.62867, 
        -49.60886, -49.59097, -49.57509, -49.56082, -49.54739, -49.5341, 
        -49.52041, -49.50605, -49.49114, -49.47597, -49.46094, -49.44644, 
        -49.43277, -49.41991, -49.4076, -49.39562, -49.38361, -49.37143, 
        -49.35912, -49.34693, -49.33509, -49.32383, -49.31333, -49.30377, 
        -49.29525,
  -48.61504, -48.68104, -48.74378, -48.80117, -48.85208, -48.89595, 
        -48.9329, -48.96383, -48.98943, -49.01009, -49.02621, -49.03809, 
        -49.04527, -49.05064, -49.05349, -49.05456, -49.05435, -49.05341, 
        -49.05238, -49.05217, -49.05366, -49.05703, -49.06215, -49.06848, 
        -49.07522, -49.08192, -49.08841, -49.09478, -49.10035, -49.1069, 
        -49.11367, -49.12041, -49.12741, -49.13528, -49.1446, -49.15569, 
        -49.16818, -49.18165, -49.19548, -49.20926, -49.22271, -49.23564, 
        -49.24779, -49.25808, -49.26847, -49.27794, -49.28703, -49.29593, 
        -49.30487, -49.31403, -49.32353, -49.33343, -49.34402, -49.35552, 
        -49.368, -49.38141, -49.39528, -49.40872, -49.4207, -49.43032, 
        -49.43613, -49.43998, -49.44095, -49.4392, -49.43524, -49.4295, 
        -49.42296, -49.41677, -49.41179, -49.40865, -49.40769, -49.40908, 
        -49.41294, -49.41873, -49.42644, -49.43522, -49.44405, -49.45174, 
        -49.45961, -49.46614, -49.47113, -49.47477, -49.47754, -49.4802, 
        -49.4831, -49.48621, -49.48926, -49.49185, -49.49358, -49.49439, 
        -49.49455, -49.49467, -49.49518, -49.49717, -49.50043, -49.5053, 
        -49.51057, -49.51787, -49.52606, -49.53432, -49.54218, -49.54947, 
        -49.55636, -49.5628, -49.56891, -49.57488, -49.58054, -49.58589, 
        -49.59084, -49.59577, -49.60096, -49.6067, -49.6131, -49.62001, 
        -49.62716, -49.63297, -49.63881, -49.64352, -49.64729, -49.6507, 
        -49.65456, -49.65952, -49.66605, -49.67467, -49.68584, -49.70004, 
        -49.71744, -49.73817, -49.76175, -49.78739, -49.81392, -49.84027, 
        -49.86589, -49.89053, -49.91418, -49.93719, -49.95884, -49.98136, 
        -50.0038, -50.02604, -50.04761, -50.06803, -50.08729, -50.10508, 
        -50.1217, -50.13783, -50.15386, -50.17038, -50.18779, -50.20645, 
        -50.22667, -50.24854, -50.27177, -50.29572, -50.31936, -50.34196, 
        -50.36317, -50.38247, -50.39994, -50.41471, -50.42905, -50.44231, 
        -50.45516, -50.46824, -50.48221, -50.49761, -50.51474, -50.53365, 
        -50.55415, -50.57589, -50.5985, -50.62127, -50.64383, -50.6661, 
        -50.68785, -50.70892, -50.72916, -50.74826, -50.76587, -50.78198, 
        -50.79683, -50.81075, -50.82405, -50.83706, -50.84941, -50.86364, 
        -50.87887, -50.89513, -50.91175, -50.92822, -50.94375, -50.95757, 
        -50.96954, -50.9796, -50.98811, -50.99557, -51.00248, -51.00906, 
        -51.01552, -51.02178, -51.02728, -51.03127, -51.03315, -51.03276, 
        -51.03025, -51.02597, -51.02007, -51.01218, -51.00225, -50.99071, 
        -50.97808, -50.96476, -50.95038, -50.93725, -50.92451, -50.91215, 
        -50.90007, -50.88829, -50.87666, -50.86554, -50.85475, -50.84402, 
        -50.83286, -50.82079, -50.80753, -50.79296, -50.7768, -50.75918, 
        -50.74, -50.7194, -50.69757, -50.67476, -50.65131, -50.6276, 
        -50.60416, -50.58123, -50.55902, -50.53736, -50.51585, -50.49398, 
        -50.4715, -50.44862, -50.42585, -50.40357, -50.38191, -50.35957, 
        -50.33814, -50.31622, -50.29359, -50.27034, -50.24649, -50.22213, 
        -50.19754, -50.17236, -50.14745, -50.12327, -50.10032, -50.07864, 
        -50.05791, -50.03773, -50.01775, -49.9978, -49.97801, -49.9583, 
        -49.93846, -49.91813, -49.89691, -49.87468, -49.85171, -49.82823, 
        -49.80451, -49.78046, -49.7562, -49.73204, -49.70855, -49.68639, 
        -49.66605, -49.64774, -49.63137, -49.61658, -49.60275, -49.58909, 
        -49.57485, -49.55994, -49.54442, -49.52866, -49.51294, -49.49678, 
        -49.48229, -49.46834, -49.45475, -49.44116, -49.42739, -49.41351, 
        -49.39969, -49.38618, -49.37323, -49.3609, -49.3494, -49.33896, 
        -49.32983,
  -48.61321, -48.67939, -48.74238, -48.80071, -48.85317, -48.89936, 
        -48.93907, -48.9717, -48.99971, -49.0225, -49.04023, -49.05335, 
        -49.06244, -49.06829, -49.07133, -49.07244, -49.07213, -49.07105, 
        -49.07002, -49.0702, -49.07203, -49.07585, -49.0803, -49.08691, 
        -49.09378, -49.10037, -49.10691, -49.11329, -49.11996, -49.127, 
        -49.13466, -49.14254, -49.15087, -49.16012, -49.17081, -49.18319, 
        -49.19707, -49.21189, -49.22603, -49.24097, -49.25539, -49.26913, 
        -49.28164, -49.29308, -49.30358, -49.31323, -49.32241, -49.33122, 
        -49.3397, -49.34826, -49.35699, -49.36604, -49.37612, -49.38751, 
        -49.39939, -49.41369, -49.42887, -49.44396, -49.45781, -49.46928, 
        -49.47786, -49.48321, -49.48524, -49.48416, -49.48022, -49.47416, 
        -49.46712, -49.46029, -49.45479, -49.45127, -49.45008, -49.4504, 
        -49.45424, -49.46034, -49.46828, -49.47752, -49.48714, -49.49658, 
        -49.50543, -49.51315, -49.51957, -49.52488, -49.52952, -49.53401, 
        -49.53864, -49.54343, -49.54813, -49.55231, -49.55563, -49.55701, 
        -49.55864, -49.56002, -49.56176, -49.56457, -49.56844, -49.57399, 
        -49.58109, -49.58958, -49.5989, -49.60805, -49.61647, -49.62392, 
        -49.63051, -49.63654, -49.64229, -49.64783, -49.65308, -49.65826, 
        -49.66224, -49.66766, -49.67366, -49.68062, -49.68872, -49.6978, 
        -49.7074, -49.7169, -49.72571, -49.73349, -49.74037, -49.74651, 
        -49.75289, -49.76007, -49.76817, -49.77793, -49.78986, -49.80434, 
        -49.82182, -49.84237, -49.86466, -49.88971, -49.91548, -49.94101, 
        -49.96564, -49.98927, -50.01194, -50.03403, -50.05604, -50.0782, 
        -50.10032, -50.12244, -50.14414, -50.16472, -50.18416, -50.20241, 
        -50.21966, -50.23655, -50.25353, -50.27102, -50.28932, -50.30879, 
        -50.32862, -50.35098, -50.37476, -50.39902, -50.42295, -50.44599, 
        -50.46749, -50.4872, -50.50499, -50.52108, -50.53572, -50.54939, 
        -50.56272, -50.57646, -50.59124, -50.60749, -50.62545, -50.6451, 
        -50.66634, -50.68877, -50.71189, -50.73518, -50.75818, -50.78056, 
        -50.80107, -50.82164, -50.84116, -50.85944, -50.87648, -50.89233, 
        -50.9071, -50.92106, -50.93434, -50.9473, -50.96048, -50.97445, 
        -50.98946, -51.00525, -51.0214, -51.03728, -51.0521, -51.06535, 
        -51.07664, -51.0861, -51.09409, -51.10109, -51.10757, -51.11392, 
        -51.1203, -51.12656, -51.1323, -51.13577, -51.13828, -51.13855, 
        -51.13624, -51.13206, -51.12591, -51.11768, -51.10739, -51.09537, 
        -51.08232, -51.06866, -51.0549, -51.04144, -51.02837, -51.01574, 
        -51.00335, -50.99117, -50.97912, -50.96721, -50.95544, -50.94364, 
        -50.93145, -50.91848, -50.90443, -50.88908, -50.8723, -50.85387, 
        -50.83394, -50.81258, -50.7899, -50.76622, -50.74089, -50.7164, 
        -50.69222, -50.66864, -50.64581, -50.62323, -50.60065, -50.5776, 
        -50.55361, -50.52899, -50.50421, -50.47996, -50.45636, -50.43313, 
        -50.40973, -50.38578, -50.36114, -50.3359, -50.31024, -50.28432, 
        -50.25828, -50.23246, -50.20714, -50.18292, -50.16006, -50.1386, 
        -50.11815, -50.09813, -50.07849, -50.05883, -50.03954, -50.01993, 
        -50.00029, -49.98003, -49.95876, -49.93638, -49.91315, -49.88942, 
        -49.86446, -49.84035, -49.81602, -49.79193, -49.76842, -49.74616, 
        -49.72557, -49.70687, -49.69, -49.67462, -49.66018, -49.64595, 
        -49.63132, -49.61589, -49.60016, -49.58401, -49.56786, -49.55225, 
        -49.53698, -49.52203, -49.50707, -49.49186, -49.47641, -49.46088, 
        -49.44555, -49.43071, -49.41665, -49.40329, -49.39083, -49.37956, 
        -49.36992,
  -48.61456, -48.68003, -48.74151, -48.79993, -48.85313, -48.90097, 
        -48.94301, -48.97934, -49.01008, -49.03487, -49.0545, -49.06915, 
        -49.07948, -49.08617, -49.08979, -49.09131, -49.08982, -49.08855, 
        -49.08759, -49.08789, -49.09005, -49.09444, -49.10043, -49.10728, 
        -49.11423, -49.12069, -49.12711, -49.13349, -49.14032, -49.14793, 
        -49.15628, -49.16523, -49.17391, -49.18461, -49.19671, -49.21049, 
        -49.22568, -49.24178, -49.2582, -49.2743, -49.28965, -49.30393, 
        -49.31698, -49.32883, -49.33971, -49.34985, -49.35945, -49.3685, 
        -49.37605, -49.384, -49.39198, -49.40021, -49.40966, -49.42083, 
        -49.43391, -49.44868, -49.46475, -49.48107, -49.49647, -49.50977, 
        -49.52029, -49.52757, -49.53136, -49.53162, -49.52857, -49.52208, 
        -49.5153, -49.50861, -49.50309, -49.49948, -49.49813, -49.49924, 
        -49.50285, -49.50882, -49.51671, -49.52588, -49.53562, -49.54528, 
        -49.55438, -49.56253, -49.56964, -49.57593, -49.58085, -49.58677, 
        -49.59296, -49.59942, -49.60589, -49.61195, -49.61731, -49.62201, 
        -49.62605, -49.62955, -49.63304, -49.63739, -49.64237, -49.649, 
        -49.65705, -49.66651, -49.67663, -49.68643, -49.69516, -49.70149, 
        -49.70763, -49.71284, -49.71767, -49.72224, -49.72659, -49.73101, 
        -49.7357, -49.74115, -49.74785, -49.75606, -49.76605, -49.77758, 
        -49.78996, -49.80257, -49.81477, -49.82613, -49.83643, -49.84605, 
        -49.85548, -49.86426, -49.8744, -49.88536, -49.89813, -49.9133, 
        -49.9308, -49.95123, -49.97396, -49.99833, -50.02322, -50.04786, 
        -50.07166, -50.09441, -50.11632, -50.13778, -50.15927, -50.18077, 
        -50.20271, -50.22455, -50.24599, -50.26631, -50.2849, -50.30355, 
        -50.32143, -50.33896, -50.35667, -50.37494, -50.39388, -50.41422, 
        -50.43597, -50.45897, -50.48339, -50.50828, -50.53283, -50.5565, 
        -50.57858, -50.59882, -50.61719, -50.63381, -50.64899, -50.66327, 
        -50.67732, -50.69195, -50.70774, -50.72388, -50.74271, -50.76281, 
        -50.78441, -50.80717, -50.83046, -50.8539, -50.87693, -50.89916, 
        -50.92032, -50.94038, -50.95932, -50.97718, -50.99396, -51.00976, 
        -51.0247, -51.03889, -51.05216, -51.0648, -51.07762, -51.09111, 
        -51.10561, -51.12069, -51.13611, -51.15125, -51.1654, -51.17694, 
        -51.18761, -51.19647, -51.20388, -51.21034, -51.21637, -51.22234, 
        -51.2285, -51.23481, -51.24086, -51.24606, -51.24941, -51.25036, 
        -51.24872, -51.24463, -51.23816, -51.22935, -51.2184, -51.2059, 
        -51.19233, -51.17833, -51.1643, -51.15052, -51.13725, -51.12426, 
        -51.11174, -51.09949, -51.08712, -51.07455, -51.06079, -51.04795, 
        -51.03467, -51.02068, -51.00572, -50.98955, -50.97187, -50.95256, 
        -50.93162, -50.90912, -50.88528, -50.8605, -50.83522, -50.80996, 
        -50.78513, -50.76098, -50.73765, -50.71442, -50.69075, -50.66654, 
        -50.64111, -50.61506, -50.58825, -50.56187, -50.53603, -50.51057, 
        -50.48499, -50.45888, -50.43214, -50.40494, -50.37756, -50.35027, 
        -50.32318, -50.29665, -50.27099, -50.24553, -50.22263, -50.20121, 
        -50.18087, -50.16126, -50.14161, -50.12205, -50.10275, -50.08349, 
        -50.06404, -50.04363, -50.02217, -49.9995, -49.97591, -49.95182, 
        -49.92759, -49.90335, -49.87909, -49.85526, -49.83202, -49.80991, 
        -49.78926, -49.77034, -49.75283, -49.73663, -49.72143, -49.70654, 
        -49.69144, -49.67585, -49.65983, -49.6436, -49.6273, -49.61128, 
        -49.59526, -49.5793, -49.56309, -49.54636, -49.5293, -49.51221, 
        -49.49549, -49.47947, -49.46426, -49.45004, -49.43659, -49.42461, 
        -49.41443,
  -48.61562, -48.68038, -48.74215, -48.79999, -48.8536, -48.90276, 
        -48.94687, -48.98577, -49.019, -49.04635, -49.06805, -49.08347, 
        -49.09497, -49.10286, -49.10731, -49.10934, -49.10904, -49.1079, 
        -49.10703, -49.10762, -49.11024, -49.11504, -49.12146, -49.12861, 
        -49.13563, -49.14226, -49.14759, -49.15397, -49.16111, -49.16922, 
        -49.17833, -49.18837, -49.19937, -49.2115, -49.22499, -49.23997, 
        -49.25637, -49.27368, -49.29122, -49.3083, -49.32442, -49.33925, 
        -49.35186, -49.36432, -49.37583, -49.3867, -49.39705, -49.4066, 
        -49.41521, -49.42291, -49.43018, -49.43781, -49.44664, -49.45754, 
        -49.47071, -49.48584, -49.50257, -49.51975, -49.53535, -49.55038, 
        -49.563, -49.57256, -49.57858, -49.58083, -49.57949, -49.57535, 
        -49.56968, -49.56382, -49.55886, -49.55553, -49.55424, -49.55505, 
        -49.55835, -49.56383, -49.57119, -49.57986, -49.58822, -49.59755, 
        -49.60629, -49.61416, -49.62121, -49.62782, -49.6344, -49.64134, 
        -49.64884, -49.65688, -49.66517, -49.67324, -49.68101, -49.68829, 
        -49.69503, -49.70133, -49.70777, -49.71421, -49.72, -49.72792, 
        -49.73726, -49.74747, -49.75827, -49.76843, -49.77734, -49.78449, 
        -49.79004, -49.79442, -49.79807, -49.80128, -49.80431, -49.80748, 
        -49.81134, -49.81663, -49.82367, -49.83333, -49.84515, -49.85814, 
        -49.87351, -49.88947, -49.9053, -49.92046, -49.93467, -49.94794, 
        -49.96075, -49.97329, -49.98592, -49.99862, -50.01237, -50.02839, 
        -50.04614, -50.06634, -50.08831, -50.1118, -50.1358, -50.15958, 
        -50.18267, -50.20492, -50.2254, -50.2464, -50.26718, -50.28816, 
        -50.30974, -50.33115, -50.3522, -50.3725, -50.39242, -50.41149, 
        -50.4299, -50.44791, -50.46614, -50.48494, -50.50473, -50.52575, 
        -50.54836, -50.57239, -50.59756, -50.6232, -50.6485, -50.67272, 
        -50.6954, -50.71529, -50.73439, -50.75177, -50.76776, -50.78296, 
        -50.7981, -50.81393, -50.8309, -50.84906, -50.86866, -50.88906, 
        -50.9108, -50.93322, -50.9561, -50.97917, -51.00187, -51.02371, 
        -51.04451, -51.06433, -51.08308, -51.10091, -51.11787, -51.13383, 
        -51.14918, -51.16232, -51.17534, -51.18767, -51.19994, -51.21276, 
        -51.22644, -51.24085, -51.2556, -51.27007, -51.28355, -51.29549, 
        -51.30557, -51.31382, -51.32055, -51.32631, -51.33165, -51.33703, 
        -51.34289, -51.34911, -51.35553, -51.36152, -51.36593, -51.36782, 
        -51.36686, -51.36283, -51.35588, -51.34623, -51.33443, -51.32011, 
        -51.30597, -51.29158, -51.27729, -51.26334, -51.24981, -51.23659, 
        -51.22422, -51.21165, -51.19913, -51.1859, -51.17258, -51.1587, 
        -51.14431, -51.12929, -51.11334, -51.09615, -51.07737, -51.05685, 
        -51.03452, -51.01062, -50.98543, -50.95939, -50.93304, -50.90689, 
        -50.88134, -50.85652, -50.83233, -50.80837, -50.78405, -50.75886, 
        -50.73243, -50.70479, -50.67535, -50.64668, -50.6184, -50.59049, 
        -50.56255, -50.53432, -50.50574, -50.47699, -50.44831, -50.41982, 
        -50.392, -50.36481, -50.33868, -50.31388, -50.29082, -50.2693, 
        -50.24873, -50.22872, -50.20891, -50.18932, -50.1699, -50.15062, 
        -50.13087, -50.11024, -50.08838, -50.06538, -50.0414, -50.01691, 
        -49.99236, -49.96801, -49.94398, -49.9205, -49.89765, -49.87586, 
        -49.85526, -49.83607, -49.81817, -49.80144, -49.78556, -49.77013, 
        -49.75364, -49.73778, -49.72174, -49.70556, -49.68919, -49.67258, 
        -49.65575, -49.63875, -49.62117, -49.60299, -49.58458, -49.56625, 
        -49.54836, -49.53125, -49.51507, -49.49986, -49.4857, -49.4732, 
        -49.46253,
  -48.61656, -48.68063, -48.74174, -48.79948, -48.85351, -48.90277, 
        -48.94859, -48.98956, -49.02503, -49.05474, -49.0786, -49.09687, 
        -49.11038, -49.11968, -49.12535, -49.12814, -49.12862, -49.12813, 
        -49.12795, -49.12893, -49.13106, -49.13611, -49.14274, -49.14996, 
        -49.15707, -49.16375, -49.17022, -49.17698, -49.18456, -49.19331, 
        -49.20317, -49.21431, -49.22656, -49.24, -49.25476, -49.27092, 
        -49.28733, -49.30556, -49.32394, -49.34176, -49.35854, -49.3741, 
        -49.38847, -49.40186, -49.41426, -49.42598, -49.437, -49.44708, 
        -49.45594, -49.46363, -49.47062, -49.47776, -49.4854, -49.49607, 
        -49.50916, -49.52449, -49.54152, -49.55941, -49.57719, -49.59389, 
        -49.60865, -49.62069, -49.62931, -49.63407, -49.63503, -49.6329, 
        -49.62891, -49.62438, -49.6204, -49.61665, -49.61551, -49.61627, 
        -49.61908, -49.62392, -49.63052, -49.63839, -49.64692, -49.65543, 
        -49.66339, -49.67059, -49.67715, -49.68354, -49.69027, -49.69775, 
        -49.70618, -49.71554, -49.72552, -49.73472, -49.74482, -49.75467, 
        -49.76431, -49.77378, -49.78311, -49.79235, -49.80171, -49.81161, 
        -49.8223, -49.83359, -49.84491, -49.85538, -49.86424, -49.87114, 
        -49.87616, -49.87979, -49.88241, -49.88445, -49.88529, -49.88741, 
        -49.89051, -49.89536, -49.90279, -49.91333, -49.927, -49.94336, 
        -49.96159, -49.98075, -50.00008, -50.01884, -50.03674, -50.05369, 
        -50.06985, -50.08536, -50.1004, -50.11532, -50.13076, -50.14742, 
        -50.16464, -50.1846, -50.20612, -50.22875, -50.25188, -50.2749, 
        -50.29739, -50.31914, -50.3402, -50.36079, -50.38126, -50.4019, 
        -50.42284, -50.44389, -50.46476, -50.48529, -50.50541, -50.52504, 
        -50.54416, -50.56293, -50.58173, -50.60112, -50.62064, -50.64262, 
        -50.66618, -50.69117, -50.71716, -50.74348, -50.76933, -50.79401, 
        -50.81714, -50.83858, -50.85837, -50.87664, -50.89373, -50.91018, 
        -50.92663, -50.94377, -50.96194, -50.98113, -51.00117, -51.02183, 
        -51.0431, -51.06492, -51.08718, -51.10961, -51.13078, -51.15231, 
        -51.17301, -51.19285, -51.21182, -51.22994, -51.24721, -51.26355, 
        -51.27882, -51.2928, -51.30549, -51.31732, -51.32897, -51.34113, 
        -51.35415, -51.36795, -51.38214, -51.39605, -51.40895, -51.4203, 
        -51.42975, -51.43734, -51.4434, -51.44849, -51.45321, -51.45802, 
        -51.4624, -51.46857, -51.47532, -51.48182, -51.48691, -51.48949, 
        -51.48888, -51.48486, -51.4775, -51.46711, -51.45433, -51.44003, 
        -51.42505, -51.41, -51.39526, -51.38103, -51.36737, -51.35434, 
        -51.3418, -51.32935, -51.31659, -51.30323, -51.28925, -51.27467, 
        -51.25946, -51.24353, -51.22655, -51.20818, -51.18808, -51.16603, 
        -51.1421, -51.11553, -51.08872, -51.06118, -51.03349, -51.00619, 
        -50.97961, -50.95384, -50.92877, -50.90397, -50.87888, -50.85286, 
        -50.82544, -50.79652, -50.76642, -50.73576, -50.70512, -50.67474, 
        -50.6445, -50.6143, -50.58409, -50.55405, -50.52438, -50.49516, 
        -50.46656, -50.43876, -50.41212, -50.38699, -50.36344, -50.34129, 
        -50.32013, -50.29953, -50.27923, -50.25916, -50.23924, -50.2193, 
        -50.19897, -50.17783, -50.15461, -50.13126, -50.10707, -50.08248, 
        -50.05792, -50.03365, -50.0098, -49.98649, -49.96391, -49.94228, 
        -49.92177, -49.90247, -49.88445, -49.86757, -49.85155, -49.83595, 
        -49.82033, -49.80449, -49.78838, -49.77197, -49.75519, -49.73798, 
        -49.72031, -49.70212, -49.68336, -49.66409, -49.64454, -49.62507, 
        -49.60607, -49.58785, -49.57061, -49.55449, -49.53973, -49.5267, 
        -49.51575,
  -48.61311, -48.67715, -48.73832, -48.79646, -48.85137, -48.90292, 
        -48.95053, -48.99351, -49.03135, -49.06343, -49.08945, -49.10977, 
        -49.12523, -49.13618, -49.14329, -49.14635, -49.14819, -49.14869, 
        -49.14927, -49.15094, -49.15441, -49.15974, -49.16646, -49.17376, 
        -49.1811, -49.18816, -49.19508, -49.20249, -49.21079, -49.22025, 
        -49.22972, -49.24193, -49.25519, -49.26982, -49.28564, -49.30273, 
        -49.32101, -49.34004, -49.35915, -49.37764, -49.39505, -49.41138, 
        -49.42672, -49.4412, -49.45476, -49.46726, -49.47779, -49.48836, 
        -49.49743, -49.50523, -49.51246, -49.51958, -49.52819, -49.53893, 
        -49.5521, -49.56749, -49.58475, -49.60313, -49.62192, -49.64014, 
        -49.65696, -49.67151, -49.68291, -49.68949, -49.69309, -49.69335, 
        -49.69144, -49.68863, -49.68596, -49.68402, -49.68323, -49.6841, 
        -49.68655, -49.69067, -49.69631, -49.70312, -49.71061, -49.71812, 
        -49.7251, -49.7314, -49.73616, -49.74197, -49.74845, -49.75611, 
        -49.76505, -49.77536, -49.7868, -49.79878, -49.81111, -49.82351, 
        -49.83602, -49.84867, -49.8613, -49.87373, -49.88596, -49.8982, 
        -49.91054, -49.92298, -49.935, -49.94479, -49.95385, -49.96086, 
        -49.96569, -49.96915, -49.97112, -49.97209, -49.9728, -49.97417, 
        -49.97647, -49.98074, -49.98821, -49.99943, -50.01477, -50.03337, 
        -50.05437, -50.07666, -50.09912, -50.12121, -50.14248, -50.16179, 
        -50.18109, -50.19937, -50.21701, -50.23404, -50.2513, -50.26926, 
        -50.28801, -50.30782, -50.32874, -50.35054, -50.37286, -50.39516, 
        -50.41719, -50.43863, -50.45951, -50.48001, -50.50033, -50.52074, 
        -50.54138, -50.56217, -50.58192, -50.60252, -50.62303, -50.64347, 
        -50.66365, -50.68339, -50.70285, -50.72269, -50.74372, -50.76651, 
        -50.79112, -50.81715, -50.8441, -50.87098, -50.89749, -50.92245, 
        -50.94574, -50.96758, -50.98798, -51.00706, -51.02532, -51.04338, 
        -51.06127, -51.07898, -51.09853, -51.1187, -51.13932, -51.15993, 
        -51.18057, -51.2014, -51.22251, -51.24415, -51.26577, -51.28711, 
        -51.30801, -51.32821, -51.34762, -51.3662, -51.38391, -51.40055, 
        -51.41587, -51.42964, -51.44194, -51.45325, -51.46432, -51.47591, 
        -51.48846, -51.50196, -51.51483, -51.52872, -51.54094, -51.55191, 
        -51.5607, -51.56756, -51.57279, -51.57704, -51.58101, -51.58511, 
        -51.5899, -51.59571, -51.60252, -51.60923, -51.6147, -51.61777, 
        -51.61744, -51.6133, -51.60549, -51.59415, -51.58012, -51.5646, 
        -51.54858, -51.53281, -51.51767, -51.50328, -51.48962, -51.47671, 
        -51.46432, -51.45097, -51.43817, -51.42458, -51.41008, -51.39476, 
        -51.37867, -51.36182, -51.34365, -51.32402, -51.30249, -51.27885, 
        -51.25318, -51.22579, -51.19721, -51.16808, -51.13897, -51.11042, 
        -51.0827, -51.0558, -51.02966, -51.00385, -50.97787, -50.95107, 
        -50.92285, -50.89283, -50.86118, -50.82844, -50.79544, -50.76268, 
        -50.73014, -50.6982, -50.66679, -50.63588, -50.60572, -50.57498, 
        -50.54582, -50.51747, -50.49013, -50.46442, -50.43993, -50.41669, 
        -50.39442, -50.3728, -50.35156, -50.33068, -50.30994, -50.28909, 
        -50.2678, -50.24578, -50.22292, -50.19921, -50.1749, -50.1503, 
        -50.1258, -50.10163, -50.07792, -50.05478, -50.03234, -50.0108, 
        -49.99035, -49.9711, -49.95334, -49.93674, -49.92102, -49.90563, 
        -49.89012, -49.87423, -49.85793, -49.84115, -49.82377, -49.80574, 
        -49.78705, -49.76782, -49.74796, -49.72793, -49.70761, -49.68748, 
        -49.66771, -49.64857, -49.62945, -49.61254, -49.59719, -49.58393, 
        -49.573,
  -48.6062, -48.67093, -48.73301, -48.79227, -48.84852, -48.90183, 
        -48.95143, -48.99656, -49.03656, -49.06994, -49.09827, -49.12099, 
        -49.13849, -49.15136, -49.16048, -49.16645, -49.16998, -49.17208, 
        -49.1737, -49.17607, -49.17977, -49.18501, -49.19156, -49.19888, 
        -49.20533, -49.21276, -49.22049, -49.22863, -49.23767, -49.24815, 
        -49.25974, -49.27267, -49.28716, -49.30291, -49.31981, -49.33787, 
        -49.35703, -49.37682, -49.3966, -49.41573, -49.43284, -49.44998, 
        -49.46626, -49.48173, -49.49625, -49.50954, -49.52181, -49.53283, 
        -49.54238, -49.55072, -49.5584, -49.56627, -49.57518, -49.58602, 
        -49.59911, -49.61428, -49.63145, -49.64909, -49.66858, -49.68812, 
        -49.70682, -49.72389, -49.73813, -49.74866, -49.75513, -49.75804, 
        -49.75844, -49.75755, -49.75629, -49.75531, -49.75507, -49.75586, 
        -49.75804, -49.76153, -49.76526, -49.771, -49.7774, -49.78386, 
        -49.7899, -49.79525, -49.80019, -49.80531, -49.81126, -49.8186, 
        -49.82769, -49.83854, -49.85094, -49.86446, -49.87866, -49.8934, 
        -49.90864, -49.9243, -49.93913, -49.95472, -49.96989, -49.9847, 
        -49.99916, -50.01303, -50.02588, -50.03725, -50.04675, -50.05421, 
        -50.05937, -50.06289, -50.06477, -50.06567, -50.06607, -50.06696, 
        -50.06892, -50.07322, -50.08094, -50.09205, -50.10869, -50.12919, 
        -50.1524, -50.17715, -50.20219, -50.22697, -50.25101, -50.27401, 
        -50.29586, -50.31661, -50.33635, -50.35541, -50.37424, -50.39337, 
        -50.41302, -50.43323, -50.45412, -50.47564, -50.49746, -50.51923, 
        -50.53971, -50.56089, -50.58162, -50.60211, -50.62253, -50.64299, 
        -50.66365, -50.68438, -50.70519, -50.72593, -50.74689, -50.76822, 
        -50.78961, -50.81046, -50.83087, -50.85146, -50.87311, -50.89668, 
        -50.92213, -50.9492, -50.97693, -51.00448, -51.03014, -51.05536, 
        -51.07897, -51.10126, -51.12236, -51.14244, -51.16194, -51.18135, 
        -51.20086, -51.22085, -51.24143, -51.26226, -51.28296, -51.30324, 
        -51.32319, -51.34312, -51.36345, -51.38453, -51.40592, -51.42736, 
        -51.44867, -51.46936, -51.48919, -51.50822, -51.52629, -51.54216, 
        -51.55751, -51.57121, -51.58323, -51.59422, -51.60493, -51.61614, 
        -51.6283, -51.64156, -51.65526, -51.66901, -51.68135, -51.69171, 
        -51.6998, -51.70591, -51.71052, -51.71427, -51.7177, -51.72131, 
        -51.7256, -51.73096, -51.73737, -51.74384, -51.74909, -51.75196, 
        -51.75146, -51.74699, -51.73745, -51.72515, -51.71, -51.69321, 
        -51.67608, -51.65946, -51.64381, -51.62923, -51.61544, -51.60264, 
        -51.5905, -51.57835, -51.56569, -51.5521, -51.53729, -51.52141, 
        -51.50455, -51.48644, -51.46717, -51.44605, -51.42299, -51.39773, 
        -51.37023, -51.34097, -51.31057, -51.27971, -51.2491, -51.21918, 
        -51.19018, -51.16215, -51.1348, -51.10791, -51.0799, -51.05214, 
        -51.02295, -50.99176, -50.95864, -50.92414, -50.88903, -50.85403, 
        -50.81957, -50.78598, -50.75326, -50.72149, -50.69052, -50.66021, 
        -50.63059, -50.60181, -50.5741, -50.54755, -50.52214, -50.49764, 
        -50.47398, -50.45108, -50.42902, -50.40669, -50.38473, -50.36263, 
        -50.34007, -50.31691, -50.29315, -50.26888, -50.24434, -50.21962, 
        -50.19508, -50.17096, -50.14721, -50.12399, -50.10142, -50.07973, 
        -50.05921, -50.03912, -50.02161, -50.00542, -49.99031, -49.97543, 
        -49.96021, -49.94411, -49.92781, -49.91082, -49.89294, -49.87427, 
        -49.85489, -49.83493, -49.81449, -49.79383, -49.77321, -49.7527, 
        -49.73256, -49.71288, -49.69418, -49.67684, -49.66135, -49.64814, 
        -49.63739,
  -48.59428, -48.66057, -48.7243, -48.78547, -48.84299, -48.89844, 
        -48.95031, -48.99789, -49.04039, -49.07726, -49.10797, -49.13305, 
        -49.15285, -49.16807, -49.17954, -49.18783, -49.19344, -49.19724, 
        -49.20019, -49.20226, -49.20612, -49.2112, -49.21736, -49.2245, 
        -49.23216, -49.24018, -49.24865, -49.25778, -49.26787, -49.27919, 
        -49.29179, -49.30598, -49.32167, -49.33871, -49.35591, -49.37512, 
        -49.39509, -49.41567, -49.43615, -49.45594, -49.47472, -49.49254, 
        -49.50953, -49.52571, -49.54094, -49.55507, -49.56802, -49.5797, 
        -49.59013, -49.59949, -49.6072, -49.61593, -49.62548, -49.6365, 
        -49.64936, -49.66421, -49.68103, -49.6996, -49.71948, -49.74004, 
        -49.76046, -49.77972, -49.79664, -49.8101, -49.8195, -49.82512, 
        -49.82792, -49.82795, -49.82816, -49.82814, -49.8284, -49.82933, 
        -49.83121, -49.83418, -49.83817, -49.84304, -49.8485, -49.85403, 
        -49.85918, -49.86372, -49.86788, -49.87226, -49.87755, -49.88441, 
        -49.8933, -49.90337, -49.91646, -49.93117, -49.94707, -49.96389, 
        -49.98156, -49.9999, -50.01856, -50.03708, -50.05512, -50.07252, 
        -50.08914, -50.10472, -50.11888, -50.13123, -50.14156, -50.14971, 
        -50.15567, -50.15966, -50.16107, -50.16251, -50.16358, -50.16492, 
        -50.16743, -50.17228, -50.18079, -50.19389, -50.21173, -50.23366, 
        -50.25848, -50.28495, -50.31198, -50.33876, -50.36479, -50.38972, 
        -50.41343, -50.43589, -50.45724, -50.47782, -50.49714, -50.51764, 
        -50.53848, -50.55965, -50.581, -50.60257, -50.62419, -50.64561, 
        -50.66672, -50.68755, -50.70823, -50.7289, -50.74966, -50.7705, 
        -50.79145, -50.8124, -50.83337, -50.85447, -50.87605, -50.89819, 
        -50.92055, -50.94254, -50.96298, -50.98447, -51.00698, -51.03123, 
        -51.05737, -51.08495, -51.11316, -51.14113, -51.16817, -51.19388, 
        -51.21822, -51.24134, -51.26345, -51.28481, -51.30569, -51.32644, 
        -51.34726, -51.36834, -51.38956, -51.41061, -51.43114, -51.45094, 
        -51.47025, -51.48855, -51.5084, -51.52907, -51.55047, -51.57226, 
        -51.59398, -51.61522, -51.63564, -51.65507, -51.6734, -51.69041, 
        -51.70583, -51.71947, -51.73148, -51.74236, -51.75289, -51.76384, 
        -51.77572, -51.78864, -51.80219, -51.81552, -51.82759, -51.83763, 
        -51.84544, -51.8513, -51.85569, -51.85827, -51.8615, -51.8648, 
        -51.86868, -51.87344, -51.87904, -51.88472, -51.88929, -51.89146, 
        -51.89022, -51.88499, -51.8756, -51.86233, -51.84611, -51.82825, 
        -51.81015, -51.79282, -51.77668, -51.76178, -51.74802, -51.73532, 
        -51.72332, -51.7114, -51.69889, -51.68525, -51.6702, -51.65371, 
        -51.63582, -51.61653, -51.5957, -51.57204, -51.54727, -51.5202, 
        -51.49095, -51.45992, -51.4278, -51.39536, -51.36327, -51.33202, 
        -51.30177, -51.27247, -51.24392, -51.2158, -51.18763, -51.15874, 
        -51.12839, -51.09598, -51.06149, -51.02541, -50.98855, -50.95172, 
        -50.91546, -50.88018, -50.84609, -50.81317, -50.78129, -50.75032, 
        -50.7202, -50.69104, -50.66291, -50.63578, -50.6095, -50.5839, 
        -50.55896, -50.53461, -50.5108, -50.48724, -50.46275, -50.43902, 
        -50.41489, -50.39029, -50.3653, -50.34007, -50.3148, -50.28963, 
        -50.26471, -50.2402, -50.21611, -50.19255, -50.16968, -50.14777, 
        -50.12717, -50.10819, -50.09096, -50.07528, -50.06063, -50.04625, 
        -50.03141, -50.01576, -49.99926, -49.9819, -49.96371, -49.94473, 
        -49.92505, -49.90483, -49.88428, -49.86362, -49.84304, -49.82267, 
        -49.80264, -49.78317, -49.76463, -49.74748, -49.73223, -49.71926, 
        -49.7087,
  -48.57708, -48.64562, -48.71181, -48.77557, -48.83683, -48.89499, 
        -48.9493, -48.99936, -49.04453, -49.08412, -49.11756, -49.1452, 
        -49.16751, -49.18436, -49.19838, -49.2092, -49.21713, -49.22295, 
        -49.22732, -49.23102, -49.235, -49.23978, -49.24557, -49.25267, 
        -49.26075, -49.26943, -49.27902, -49.2893, -49.30054, -49.312, 
        -49.32587, -49.34131, -49.35828, -49.3767, -49.39628, -49.41663, 
        -49.4375, -49.45883, -49.47992, -49.50042, -49.51995, -49.5385, 
        -49.55609, -49.57282, -49.58754, -49.60223, -49.61579, -49.6283, 
        -49.63971, -49.65034, -49.66048, -49.67046, -49.68079, -49.69208, 
        -49.70474, -49.71911, -49.73542, -49.75359, -49.77366, -49.79505, 
        -49.81685, -49.83707, -49.85636, -49.87246, -49.88456, -49.89278, 
        -49.8979, -49.90093, -49.90261, -49.90363, -49.9045, -49.90564, 
        -49.90739, -49.91002, -49.91335, -49.91737, -49.92193, -49.9267, 
        -49.9311, -49.934, -49.93757, -49.94134, -49.94601, -49.95235, 
        -49.96096, -49.97205, -49.98568, -50.00148, -50.01871, -50.03732, 
        -50.05686, -50.07744, -50.09846, -50.11942, -50.14023, -50.16022, 
        -50.17917, -50.19571, -50.21146, -50.22517, -50.23674, -50.2462, 
        -50.25347, -50.25874, -50.26242, -50.26515, -50.26758, -50.27033, 
        -50.27412, -50.28028, -50.28987, -50.30402, -50.32286, -50.34568, 
        -50.37153, -50.39912, -50.4274, -50.45433, -50.48164, -50.5079, 
        -50.53268, -50.55627, -50.57866, -50.60025, -50.62194, -50.6441, 
        -50.66642, -50.68884, -50.71108, -50.7331, -50.75474, -50.77589, 
        -50.79663, -50.81719, -50.83778, -50.85887, -50.88034, -50.90193, 
        -50.92249, -50.94399, -50.96535, -50.98687, -51.00891, -51.03174, 
        -51.05503, -51.07816, -51.10069, -51.12319, -51.14669, -51.17153, 
        -51.19828, -51.22628, -51.25474, -51.28304, -51.31057, -51.33698, 
        -51.36227, -51.38654, -51.41001, -51.43277, -51.45413, -51.47625, 
        -51.4982, -51.51995, -51.54155, -51.56251, -51.58296, -51.60225, 
        -51.62122, -51.64015, -51.65982, -51.68051, -51.70215, -51.72438, 
        -51.7466, -51.76831, -51.78912, -51.80885, -51.82724, -51.84424, 
        -51.8596, -51.87305, -51.88523, -51.89622, -51.90683, -51.91673, 
        -51.9284, -51.94095, -51.95406, -51.96697, -51.97871, -51.98838, 
        -51.99616, -52.00228, -52.00671, -52.01059, -52.01393, -52.01716, 
        -52.02069, -52.02481, -52.02947, -52.03389, -52.03712, -52.03807, 
        -52.03564, -52.0295, -52.01925, -52.00518, -51.98816, -51.96951, 
        -51.95066, -51.93275, -51.91627, -51.9011, -51.88631, -51.87369, 
        -51.86173, -51.84982, -51.83719, -51.82324, -51.8076, -51.79021, 
        -51.77118, -51.75037, -51.72787, -51.70345, -51.67688, -51.64814, 
        -51.61724, -51.58464, -51.55103, -51.51725, -51.48392, -51.45153, 
        -51.41999, -51.3894, -51.35951, -51.33, -51.30044, -51.27012, 
        -51.23847, -51.20475, -51.16896, -51.13155, -51.09327, -51.05488, 
        -51.01702, -50.97913, -50.94353, -50.90946, -50.87646, -50.84481, 
        -50.81405, -50.7846, -50.75607, -50.7284, -50.7013, -50.6745, 
        -50.64824, -50.6223, -50.59674, -50.57143, -50.54611, -50.52041, 
        -50.49455, -50.46825, -50.44174, -50.41523, -50.38896, -50.36294, 
        -50.33718, -50.31187, -50.28704, -50.2628, -50.23943, -50.21724, 
        -50.19654, -50.17763, -50.16071, -50.14544, -50.13126, -50.11737, 
        -50.10284, -50.08727, -50.07071, -50.05308, -50.03475, -50.01561, 
        -49.996, -49.97601, -49.95487, -49.93464, -49.91455, -49.89491, 
        -49.87565, -49.85719, -49.83959, -49.82329, -49.80876, -49.79636, 
        -49.78615,
  -48.55737, -48.62886, -48.69833, -48.76539, -48.82982, -48.89106, 
        -48.94836, -49.00098, -49.04763, -49.08976, -49.12578, -49.15612, 
        -49.18121, -49.20188, -49.21864, -49.23214, -49.24248, -49.25018, 
        -49.25595, -49.26062, -49.26485, -49.26968, -49.27553, -49.28178, 
        -49.29021, -49.29989, -49.31056, -49.32214, -49.33479, -49.3487, 
        -49.36399, -49.38093, -49.39941, -49.4192, -49.43997, -49.46113, 
        -49.48301, -49.50498, -49.52682, -49.547, -49.5673, -49.58646, 
        -49.60451, -49.62149, -49.63758, -49.65276, -49.66696, -49.68036, 
        -49.69299, -49.7051, -49.71678, -49.72825, -49.73958, -49.75124, 
        -49.7638, -49.77672, -49.79247, -49.81034, -49.83033, -49.85208, 
        -49.87486, -49.89759, -49.91883, -49.93718, -49.95171, -49.96239, 
        -49.9698, -49.97474, -49.97793, -49.97997, -49.98144, -49.98286, 
        -49.98344, -49.98564, -49.98853, -49.99205, -49.99601, -50.00006, 
        -50.00387, -50.00734, -50.01057, -50.014, -50.01834, -50.02422, 
        -50.03284, -50.04435, -50.05856, -50.07515, -50.09361, -50.1135, 
        -50.13357, -50.15549, -50.17834, -50.20158, -50.22441, -50.24686, 
        -50.26804, -50.28779, -50.30547, -50.32088, -50.33417, -50.3453, 
        -50.35436, -50.36153, -50.36718, -50.37193, -50.37661, -50.38157, 
        -50.38764, -50.39474, -50.40594, -50.4215, -50.44098, -50.4645, 
        -50.49087, -50.51875, -50.54736, -50.57581, -50.60365, -50.63038, 
        -50.6559, -50.68002, -50.70298, -50.72581, -50.7487, -50.77209, 
        -50.79589, -50.81971, -50.84309, -50.86579, -50.88674, -50.90795, 
        -50.92857, -50.94905, -50.9699, -50.99141, -51.01347, -51.0361, 
        -51.05872, -51.08105, -51.1031, -51.12535, -51.14805, -51.17145, 
        -51.19522, -51.21901, -51.24242, -51.26596, -51.29022, -51.31582, 
        -51.3429, -51.37106, -51.39877, -51.42739, -51.4556, -51.48307, 
        -51.50966, -51.5355, -51.56054, -51.58503, -51.60896, -51.63242, 
        -51.65536, -51.67772, -51.69966, -51.72064, -51.74047, -51.75974, 
        -51.77845, -51.79737, -51.81715, -51.83815, -51.86011, -51.88278, 
        -51.90538, -51.92735, -51.94737, -51.96718, -51.98561, -52.00247, 
        -52.01772, -52.03127, -52.04334, -52.05457, -52.06541, -52.07644, 
        -52.08799, -52.1001, -52.11248, -52.12497, -52.13633, -52.14585, 
        -52.15401, -52.16032, -52.16531, -52.16943, -52.17318, -52.17659, 
        -52.17991, -52.18335, -52.18685, -52.18987, -52.19149, -52.1898, 
        -52.186, -52.17856, -52.16745, -52.15283, -52.13533, -52.11628, 
        -52.09696, -52.07866, -52.06185, -52.04662, -52.03285, -52.02026, 
        -52.0083, -51.99617, -51.98301, -51.96833, -51.95182, -51.93325, 
        -51.91263, -51.8901, -51.86562, -51.83929, -51.81096, -51.7805, 
        -51.74806, -51.7141, -51.67932, -51.64452, -51.6102, -51.57667, 
        -51.54297, -51.51102, -51.47965, -51.4486, -51.41747, -51.38562, 
        -51.3524, -51.31716, -51.28029, -51.24179, -51.20236, -51.16277, 
        -51.1236, -51.08536, -51.04841, -51.01279, -50.97872, -50.94617, 
        -50.91471, -50.88482, -50.85582, -50.82777, -50.80001, -50.77234, 
        -50.74469, -50.71716, -50.68972, -50.6624, -50.63498, -50.60727, 
        -50.5791, -50.55092, -50.52261, -50.49447, -50.46667, -50.4392, 
        -50.41212, -50.38551, -50.35952, -50.33331, -50.30942, -50.28691, 
        -50.26613, -50.24727, -50.23043, -50.21522, -50.20107, -50.18714, 
        -50.17264, -50.15708, -50.14037, -50.1227, -50.10427, -50.08545, 
        -50.06617, -50.0468, -50.02741, -50.00819, -49.98924, -49.97086, 
        -49.95327, -49.93661, -49.92077, -49.90609, -49.89273, -49.88123, 
        -49.87127,
  -48.53508, -48.6101, -48.68322, -48.75311, -48.82104, -48.88544, 
        -48.94583, -49.00122, -49.05142, -49.096, -49.13472, -49.16762, 
        -49.19531, -49.21854, -49.23814, -49.25431, -49.26732, -49.27615, 
        -49.2834, -49.28902, -49.29409, -49.29941, -49.30568, -49.31347, 
        -49.32278, -49.33361, -49.3456, -49.3588, -49.37305, -49.38843, 
        -49.40549, -49.42391, -49.44379, -49.46368, -49.48524, -49.50736, 
        -49.52989, -49.55248, -49.57511, -49.59718, -49.61829, -49.63799, 
        -49.65644, -49.67369, -49.68998, -49.70546, -49.72022, -49.7346, 
        -49.74857, -49.76128, -49.77457, -49.78746, -49.7999, -49.81219, 
        -49.82481, -49.83846, -49.85378, -49.87119, -49.89101, -49.91299, 
        -49.93637, -49.96008, -49.98279, -50.00297, -50.01964, -50.03261, 
        -50.04127, -50.0481, -50.05273, -50.05572, -50.0577, -50.05927, 
        -50.06086, -50.06287, -50.06549, -50.06866, -50.07216, -50.07569, 
        -50.07897, -50.08232, -50.08552, -50.08883, -50.09349, -50.09867, 
        -50.10754, -50.11939, -50.13422, -50.1517, -50.17117, -50.19214, 
        -50.21432, -50.23753, -50.26153, -50.28597, -50.3107, -50.33501, 
        -50.35831, -50.38025, -50.40006, -50.41755, -50.4327, -50.44572, 
        -50.45612, -50.4657, -50.47397, -50.48162, -50.48924, -50.49726, 
        -50.50631, -50.51692, -50.53009, -50.54683, -50.56725, -50.59111, 
        -50.61731, -50.64501, -50.67319, -50.70142, -50.72929, -50.75607, 
        -50.78152, -50.8061, -50.82888, -50.85237, -50.87622, -50.90069, 
        -50.92599, -50.95116, -50.97573, -50.99941, -51.02203, -51.04367, 
        -51.06463, -51.08543, -51.10666, -51.12868, -51.15161, -51.17519, 
        -51.19904, -51.2225, -51.24573, -51.26885, -51.29221, -51.31506, 
        -51.33916, -51.36343, -51.38748, -51.41172, -51.43674, -51.46291, 
        -51.49019, -51.51849, -51.54736, -51.57632, -51.60548, -51.63406, 
        -51.6622, -51.68965, -51.71657, -51.74286, -51.76846, -51.79332, 
        -51.81725, -51.84032, -51.86255, -51.88358, -51.90322, -51.92147, 
        -51.94046, -51.95969, -51.97984, -52.00119, -52.02346, -52.04624, 
        -52.06894, -52.09101, -52.11206, -52.13182, -52.15017, -52.16692, 
        -52.182, -52.19553, -52.20773, -52.21921, -52.23035, -52.24158, 
        -52.2531, -52.26495, -52.27687, -52.2888, -52.29959, -52.30944, 
        -52.31732, -52.32312, -52.32825, -52.33332, -52.33744, -52.34092, 
        -52.34422, -52.34704, -52.34948, -52.35113, -52.35096, -52.34852, 
        -52.34317, -52.33449, -52.3226, -52.30736, -52.2897, -52.27051, 
        -52.2512, -52.2328, -52.2159, -52.20066, -52.18702, -52.1745, 
        -52.16231, -52.14955, -52.13552, -52.11964, -52.10171, -52.08154, 
        -52.05819, -52.03362, -52.00705, -51.97866, -51.94848, -51.91642, 
        -51.88265, -51.84762, -51.81196, -51.77639, -51.74134, -51.70673, 
        -51.67276, -51.63929, -51.60628, -51.57355, -51.54071, -51.50721, 
        -51.4724, -51.43578, -51.39772, -51.35829, -51.31799, -51.27746, 
        -51.23723, -51.19783, -51.15966, -51.12292, -51.08773, -51.05396, 
        -51.02187, -50.99139, -50.96198, -50.93337, -50.90508, -50.8756, 
        -50.84679, -50.81765, -50.78831, -50.7588, -50.72905, -50.69897, 
        -50.66859, -50.63813, -50.60776, -50.57766, -50.54794, -50.51852, 
        -50.48958, -50.4613, -50.4339, -50.40772, -50.38301, -50.3601, 
        -50.33921, -50.3202, -50.30302, -50.28724, -50.27245, -50.25804, 
        -50.24307, -50.2272, -50.2103, -50.19254, -50.17425, -50.15572, 
        -50.13715, -50.11876, -50.10052, -50.08262, -50.06542, -50.04909, 
        -50.03377, -50.01957, -50.00614, -49.99357, -49.982, -49.97147, 
        -49.96194,
  -48.50956, -48.58907, -48.66609, -48.74084, -48.81234, -48.88008, 
        -48.94317, -49.00134, -49.05405, -49.10101, -49.14215, -49.17767, 
        -49.2071, -49.23302, -49.25526, -49.27404, -49.28935, -49.30146, 
        -49.31061, -49.31768, -49.3241, -49.33053, -49.33796, -49.34697, 
        -49.35756, -49.36982, -49.38343, -49.39729, -49.41341, -49.43065, 
        -49.44909, -49.46865, -49.48951, -49.51115, -49.53352, -49.5563, 
        -49.57932, -49.60278, -49.62617, -49.64917, -49.67113, -49.69163, 
        -49.7105, -49.72678, -49.74328, -49.75916, -49.77442, -49.7897, 
        -49.8049, -49.82006, -49.83501, -49.84938, -49.86298, -49.87605, 
        -49.88903, -49.90269, -49.9178, -49.93503, -49.95465, -49.97556, 
        -49.99918, -50.02348, -50.04711, -50.06871, -50.08728, -50.10235, 
        -50.11415, -50.12283, -50.12884, -50.13271, -50.13517, -50.13702, 
        -50.13873, -50.14076, -50.14333, -50.14632, -50.14951, -50.1517, 
        -50.15483, -50.15797, -50.16151, -50.16546, -50.17049, -50.17731, 
        -50.18681, -50.19935, -50.21505, -50.23341, -50.25381, -50.27572, 
        -50.29878, -50.32274, -50.34751, -50.37294, -50.39875, -50.42351, 
        -50.44877, -50.47267, -50.49463, -50.51426, -50.53176, -50.54705, 
        -50.56062, -50.5732, -50.5846, -50.59563, -50.60674, -50.61833, 
        -50.63065, -50.6442, -50.65976, -50.67807, -50.69889, -50.72259, 
        -50.74738, -50.77443, -50.80205, -50.82966, -50.85708, -50.8836, 
        -50.90912, -50.93371, -50.95778, -50.98193, -51.00663, -51.03204, 
        -51.05841, -51.08492, -51.1107, -51.13549, -51.15925, -51.18195, 
        -51.20388, -51.22554, -51.24753, -51.26936, -51.29316, -51.31774, 
        -51.34265, -51.36741, -51.39183, -51.41597, -51.44006, -51.46431, 
        -51.48875, -51.51329, -51.5378, -51.56258, -51.58836, -51.61504, 
        -51.64254, -51.67091, -51.70002, -51.7297, -51.75952, -51.78933, 
        -51.81886, -51.84791, -51.87546, -51.9036, -51.93103, -51.95747, 
        -51.98272, -52.00671, -52.0294, -52.05092, -52.07114, -52.09053, 
        -52.10982, -52.12963, -52.15033, -52.17199, -52.19436, -52.21698, 
        -52.23944, -52.26125, -52.28198, -52.30161, -52.31985, -52.33644, 
        -52.35146, -52.36501, -52.37739, -52.38816, -52.39965, -52.41107, 
        -52.42257, -52.43432, -52.44615, -52.4577, -52.4685, -52.47807, 
        -52.48617, -52.49281, -52.49863, -52.50345, -52.50786, -52.51142, 
        -52.51464, -52.51708, -52.51868, -52.51896, -52.51729, -52.51329, 
        -52.50644, -52.49664, -52.48373, -52.4681, -52.45036, -52.43131, 
        -52.41221, -52.39286, -52.37602, -52.36088, -52.34725, -52.33471, 
        -52.32225, -52.30874, -52.2935, -52.27597, -52.25622, -52.23409, 
        -52.20966, -52.18295, -52.15424, -52.12382, -52.09184, -52.05834, 
        -52.02346, -51.98757, -51.95131, -51.91515, -51.87922, -51.8437, 
        -51.80844, -51.77347, -51.73867, -51.70417, -51.66952, -51.63419, 
        -51.59774, -51.55981, -51.52056, -51.48021, -51.43819, -51.39697, 
        -51.35595, -51.31569, -51.27654, -51.23882, -51.20261, -51.1682, 
        -51.13535, -51.10402, -51.0739, -51.04475, -51.0158, -50.9867, 
        -50.9568, -50.92596, -50.89467, -50.86286, -50.83067, -50.798, 
        -50.7652, -50.73245, -50.69992, -50.66758, -50.63551, -50.60387, 
        -50.57287, -50.54275, -50.51386, -50.48656, -50.46112, -50.43769, 
        -50.41618, -50.39661, -50.37859, -50.36179, -50.34576, -50.32978, 
        -50.31371, -50.29725, -50.27993, -50.26106, -50.24292, -50.22491, 
        -50.20692, -50.1895, -50.17274, -50.15663, -50.1416, -50.12776, 
        -50.11526, -50.10387, -50.09329, -50.08322, -50.07354, -50.06426, 
        -50.05532,
  -48.48346, -48.56753, -48.64923, -48.72787, -48.80294, -48.87368, 
        -48.93848, -48.99907, -49.05403, -49.10311, -49.14638, -49.18445, 
        -49.21756, -49.24635, -49.27149, -49.29285, -49.31068, -49.32489, 
        -49.3359, -49.34502, -49.35316, -49.3605, -49.36987, -49.38066, 
        -49.3932, -49.40724, -49.42281, -49.43955, -49.45753, -49.47633, 
        -49.49611, -49.51672, -49.53821, -49.56041, -49.58307, -49.60628, 
        -49.63008, -49.65337, -49.6778, -49.70176, -49.7245, -49.74577, 
        -49.76511, -49.78297, -49.79969, -49.81558, -49.83133, -49.84733, 
        -49.86357, -49.87998, -49.89633, -49.91215, -49.92705, -49.94013, 
        -49.95377, -49.96782, -49.98308, -50.00027, -50.0198, -50.04163, 
        -50.06523, -50.08968, -50.11373, -50.13641, -50.15658, -50.17366, 
        -50.18751, -50.19788, -50.20518, -50.20999, -50.21213, -50.2145, 
        -50.21654, -50.21893, -50.22169, -50.22468, -50.22765, -50.2306, 
        -50.23365, -50.23707, -50.24087, -50.2455, -50.25135, -50.25919, 
        -50.26968, -50.28327, -50.29995, -50.31932, -50.33969, -50.3625, 
        -50.38632, -50.41087, -50.43611, -50.4621, -50.4887, -50.51561, 
        -50.54222, -50.5678, -50.59174, -50.61354, -50.63331, -50.65119, 
        -50.66769, -50.68299, -50.69789, -50.71252, -50.72742, -50.74171, 
        -50.7575, -50.77407, -50.792, -50.81139, -50.8327, -50.85602, 
        -50.88118, -50.90755, -50.93445, -50.96141, -50.98817, -51.01411, 
        -51.03938, -51.06402, -51.08844, -51.11329, -51.1389, -51.16512, 
        -51.19231, -51.21979, -51.24585, -51.27182, -51.29718, -51.32157, 
        -51.34514, -51.36846, -51.39175, -51.41552, -51.44021, -51.46562, 
        -51.4916, -51.51765, -51.5432, -51.56839, -51.59337, -51.61824, 
        -51.64293, -51.66784, -51.69284, -51.71832, -51.74466, -51.77071, 
        -51.79849, -51.82708, -51.85647, -51.88659, -51.91718, -51.94798, 
        -51.97853, -52.00891, -52.03903, -52.06896, -52.09838, -52.12677, 
        -52.15373, -52.17904, -52.2027, -52.22489, -52.24581, -52.26597, 
        -52.28602, -52.30646, -52.32766, -52.34959, -52.37182, -52.39315, 
        -52.41516, -52.43635, -52.45662, -52.47577, -52.49363, -52.51002, 
        -52.52501, -52.5387, -52.5513, -52.56356, -52.57523, -52.58673, 
        -52.59822, -52.60991, -52.62178, -52.63345, -52.64436, -52.65398, 
        -52.66216, -52.66898, -52.67454, -52.6793, -52.68351, -52.68696, 
        -52.69006, -52.69234, -52.69234, -52.69167, -52.68876, -52.68337, 
        -52.67519, -52.66418, -52.65043, -52.63429, -52.61636, -52.59755, 
        -52.57866, -52.56059, -52.54386, -52.5288, -52.51512, -52.50234, 
        -52.48924, -52.4747, -52.45797, -52.43867, -52.41689, -52.39266, 
        -52.36603, -52.33723, -52.30649, -52.27418, -52.24054, -52.20577, 
        -52.16999, -52.13348, -52.09666, -52.05876, -52.02208, -51.98559, 
        -51.94906, -51.91255, -51.87601, -51.8396, -51.80298, -51.76579, 
        -51.72767, -51.68837, -51.64797, -51.60678, -51.56514, -51.52345, 
        -51.48198, -51.44114, -51.40139, -51.363, -51.32622, -51.2911, 
        -51.25748, -51.22538, -51.19447, -51.16446, -51.13464, -51.10444, 
        -51.07331, -51.04083, -51.00773, -50.97356, -50.93876, -50.90358, 
        -50.86841, -50.83339, -50.79853, -50.7638, -50.72833, -50.69432, 
        -50.6612, -50.62928, -50.59895, -50.57047, -50.54405, -50.51973, 
        -50.49731, -50.47656, -50.45729, -50.43866, -50.42081, -50.40329, 
        -50.38536, -50.36742, -50.3494, -50.33115, -50.31301, -50.29519, 
        -50.27798, -50.2617, -50.24643, -50.23238, -50.21973, -50.20859, 
        -50.19889, -50.19043, -50.18276, -50.17524, -50.16755, -50.15962, 
        -50.15166,
  -48.4557, -48.54394, -48.63021, -48.71289, -48.79132, -48.86483, 
        -48.93289, -48.99561, -49.05246, -49.10366, -49.14924, -49.18938, 
        -49.2252, -49.25694, -49.285, -49.30922, -49.3286, -49.34515, 
        -49.35852, -49.3697, -49.37997, -49.39058, -49.40236, -49.41572, 
        -49.43078, -49.4472, -49.46507, -49.48409, -49.50386, -49.52439, 
        -49.5453, -49.56577, -49.58757, -49.60984, -49.6327, -49.6564, 
        -49.68099, -49.70625, -49.73162, -49.7566, -49.78055, -49.80275, 
        -49.82272, -49.84119, -49.85815, -49.87433, -49.89021, -49.90556, 
        -49.92247, -49.93984, -49.95736, -49.97451, -49.9908, -50.00617, 
        -50.02097, -50.03587, -50.0517, -50.06912, -50.08865, -50.11033, 
        -50.1337, -50.15799, -50.18225, -50.20555, -50.22604, -50.24493, 
        -50.26062, -50.27278, -50.28157, -50.2877, -50.2917, -50.29486, 
        -50.2978, -50.3007, -50.30381, -50.3068, -50.30968, -50.31246, 
        -50.31557, -50.31911, -50.32335, -50.32863, -50.33442, -50.3434, 
        -50.35516, -50.36996, -50.38791, -50.4084, -50.43086, -50.45459, 
        -50.47908, -50.50418, -50.52988, -50.55631, -50.58351, -50.6111, 
        -50.63867, -50.66552, -50.69106, -50.7149, -50.73598, -50.75653, 
        -50.77594, -50.79466, -50.81302, -50.8312, -50.84956, -50.86818, 
        -50.88701, -50.90615, -50.92573, -50.94619, -50.96798, -50.99139, 
        -51.01637, -51.04242, -51.06901, -51.09565, -51.12197, -51.14767, 
        -51.17174, -51.19651, -51.2212, -51.24627, -51.27234, -51.29939, 
        -51.32726, -51.35544, -51.38354, -51.41099, -51.43804, -51.46439, 
        -51.49014, -51.51542, -51.54054, -51.56588, -51.59175, -51.61822, 
        -51.64513, -51.67224, -51.69922, -51.72466, -51.7506, -51.77606, 
        -51.80139, -51.82686, -51.85231, -51.87833, -51.90503, -51.93246, 
        -51.96057, -51.9894, -52.01915, -52.04965, -52.08069, -52.11198, 
        -52.14344, -52.17482, -52.20635, -52.23814, -52.26965, -52.30022, 
        -52.32916, -52.35602, -52.38012, -52.40342, -52.42544, -52.44672, 
        -52.46781, -52.48914, -52.51088, -52.53291, -52.55503, -52.57701, 
        -52.59825, -52.61896, -52.6382, -52.65656, -52.67377, -52.68977, 
        -52.70459, -52.7184, -52.7314, -52.74381, -52.75563, -52.76727, 
        -52.77885, -52.79071, -52.80285, -52.81493, -52.82529, -52.83536, 
        -52.84383, -52.85077, -52.85629, -52.86061, -52.8643, -52.86744, 
        -52.87024, -52.87221, -52.87267, -52.87121, -52.86727, -52.86092, 
        -52.85172, -52.83965, -52.825, -52.80828, -52.79016, -52.77148, 
        -52.75264, -52.73473, -52.7181, -52.70295, -52.6889, -52.67538, 
        -52.6612, -52.64534, -52.62706, -52.60501, -52.58128, -52.55502, 
        -52.52635, -52.49559, -52.46306, -52.42908, -52.39406, -52.35822, 
        -52.32166, -52.28451, -52.247, -52.20937, -52.17176, -52.13419, 
        -52.09647, -52.05849, -52.02024, -51.98195, -51.94329, -51.90421, 
        -51.86444, -51.82375, -51.78228, -51.74033, -51.69827, -51.6563, 
        -51.61466, -51.57378, -51.53389, -51.49532, -51.45807, -51.42236, 
        -51.38801, -51.3549, -51.32182, -51.29037, -51.25904, -51.22723, 
        -51.19441, -51.16033, -51.12485, -51.08876, -51.05184, -51.01463, 
        -50.97736, -50.94014, -50.90297, -50.86589, -50.82911, -50.79293, 
        -50.75777, -50.72411, -50.69221, -50.66239, -50.63471, -50.60913, 
        -50.58541, -50.56325, -50.54213, -50.52184, -50.50192, -50.48214, 
        -50.46207, -50.44214, -50.42252, -50.40337, -50.38471, -50.36691, 
        -50.35023, -50.33495, -50.32128, -50.30933, -50.29914, -50.29065, 
        -50.28366, -50.2778, -50.27265, -50.26736, -50.26153, -50.25412, 
        -50.24755,
  -48.42575, -48.5201, -48.61108, -48.6978, -48.77954, -48.85552, 
        -48.92594, -48.99042, -49.04891, -49.10193, -49.14848, -49.19104, 
        -49.22922, -49.26376, -49.29454, -49.32153, -49.34457, -49.36372, 
        -49.37956, -49.3933, -49.40621, -49.41942, -49.43409, -49.45041, 
        -49.46844, -49.48783, -49.50754, -49.52905, -49.55119, -49.57347, 
        -49.59558, -49.6176, -49.63962, -49.66188, -49.685, -49.70922, 
        -49.73447, -49.76069, -49.78717, -49.81329, -49.83813, -49.86021, 
        -49.88123, -49.90025, -49.91768, -49.93409, -49.95012, -49.96649, 
        -49.98376, -50.00187, -50.02044, -50.03883, -50.05655, -50.07341, 
        -50.08957, -50.10572, -50.12249, -50.14043, -50.15902, -50.18059, 
        -50.20367, -50.22774, -50.25209, -50.27591, -50.29848, -50.3189, 
        -50.33638, -50.35039, -50.36093, -50.36854, -50.37408, -50.3785, 
        -50.38244, -50.38621, -50.38963, -50.39172, -50.39447, -50.39704, 
        -50.40017, -50.4038, -50.40824, -50.41413, -50.42184, -50.4321, 
        -50.44522, -50.46146, -50.48082, -50.50262, -50.52621, -50.55088, 
        -50.57607, -50.60171, -50.62783, -50.65355, -50.68114, -50.70925, 
        -50.73737, -50.76507, -50.79196, -50.81763, -50.84184, -50.86504, 
        -50.88744, -50.90943, -50.93113, -50.95261, -50.97402, -50.99545, 
        -51.0168, -51.03793, -51.059, -51.08052, -51.103, -51.12592, 
        -51.15123, -51.17755, -51.20439, -51.23109, -51.25763, -51.28342, 
        -51.3086, -51.33348, -51.35844, -51.38397, -51.41043, -51.43788, 
        -51.4662, -51.49507, -51.52393, -51.55267, -51.58131, -51.60971, 
        -51.63773, -51.66431, -51.69148, -51.71865, -51.74635, -51.77422, 
        -51.80247, -51.83087, -51.85898, -51.88669, -51.91384, -51.94032, 
        -51.96636, -51.99236, -52.01844, -52.04486, -52.07179, -52.09929, 
        -52.12758, -52.15676, -52.18676, -52.21752, -52.24877, -52.28033, 
        -52.3112, -52.34355, -52.37661, -52.41027, -52.44386, -52.47658, 
        -52.50758, -52.53636, -52.56277, -52.58769, -52.61121, -52.63401, 
        -52.65656, -52.67904, -52.70148, -52.72382, -52.7458, -52.76723, 
        -52.78782, -52.80742, -52.82592, -52.84332, -52.85966, -52.87501, 
        -52.88858, -52.90224, -52.91534, -52.92794, -52.94001, -52.95173, 
        -52.96348, -52.97562, -52.98824, -53.00092, -53.01297, -53.02377, 
        -53.03289, -53.04016, -53.04563, -53.04962, -53.05276, -53.05547, 
        -53.05781, -53.05929, -53.05926, -53.05704, -53.05244, -53.04499, 
        -53.03505, -53.02208, -53.00663, -52.98933, -52.96995, -52.95112, 
        -52.93245, -52.91457, -52.89789, -52.88219, -52.86744, -52.85258, 
        -52.83702, -52.81958, -52.79949, -52.77678, -52.7513, -52.72327, 
        -52.69289, -52.66051, -52.62647, -52.59114, -52.55499, -52.51817, 
        -52.48085, -52.44295, -52.40454, -52.36588, -52.32713, -52.28837, 
        -52.2494, -52.21, -52.17017, -52.12996, -52.08941, -52.04856, 
        -52.00613, -51.96416, -51.92177, -51.87932, -51.83704, -51.79507, 
        -51.75362, -51.71284, -51.67314, -51.63469, -51.59729, -51.56097, 
        -51.52554, -51.49126, -51.45755, -51.42416, -51.39073, -51.35677, 
        -51.32191, -51.28579, -51.24854, -51.21056, -51.17177, -51.13293, 
        -51.09375, -51.05465, -51.01539, -50.97615, -50.93732, -50.89917, 
        -50.86214, -50.82671, -50.79316, -50.76173, -50.73249, -50.70549, 
        -50.68016, -50.65604, -50.6332, -50.61095, -50.58778, -50.56542, 
        -50.5429, -50.52058, -50.4989, -50.47819, -50.45861, -50.44046, 
        -50.42403, -50.40957, -50.3973, -50.38724, -50.37933, -50.37317, 
        -50.36852, -50.36475, -50.36167, -50.3581, -50.35387, -50.34916, 
        -50.34438,
  -48.39558, -48.49541, -48.59116, -48.68172, -48.76666, -48.84443, 
        -48.91685, -48.98288, -49.04295, -49.0974, -49.14676, -49.1914, 
        -49.23187, -49.26875, -49.30193, -49.33139, -49.35691, -49.37876, 
        -49.39734, -49.41412, -49.42924, -49.44582, -49.46383, -49.48351, 
        -49.5048, -49.52766, -49.5515, -49.5761, -49.60085, -49.62516, 
        -49.64866, -49.67154, -49.694, -49.71661, -49.73986, -49.76344, 
        -49.78925, -49.8162, -49.84359, -49.87072, -49.89661, -49.92071, 
        -49.94257, -49.96247, -49.9804, -49.99696, -50.01319, -50.02979, 
        -50.04734, -50.06587, -50.08525, -50.10479, -50.12287, -50.14122, 
        -50.15892, -50.17638, -50.19412, -50.2127, -50.23264, -50.25416, 
        -50.27711, -50.30111, -50.3256, -50.34998, -50.37353, -50.39537, 
        -50.41461, -50.4306, -50.44321, -50.45185, -50.45928, -50.46534, 
        -50.47055, -50.47516, -50.47908, -50.48226, -50.48488, -50.48732, 
        -50.49009, -50.49365, -50.49836, -50.5047, -50.51323, -50.52457, 
        -50.53912, -50.55695, -50.57678, -50.59995, -50.6247, -50.65028, 
        -50.67619, -50.70236, -50.72888, -50.75599, -50.78375, -50.81199, 
        -50.84048, -50.86886, -50.89679, -50.92395, -50.95024, -50.97592, 
        -51.00116, -51.02617, -51.0509, -51.07427, -51.09834, -51.12203, 
        -51.14537, -51.16824, -51.19074, -51.21344, -51.23693, -51.26175, 
        -51.28791, -51.31503, -51.34262, -51.37011, -51.39718, -51.42358, 
        -51.4493, -51.47472, -51.50018, -51.52612, -51.55286, -51.57955, 
        -51.60812, -51.63727, -51.66681, -51.69663, -51.7267, -51.75691, 
        -51.78704, -51.81693, -51.84653, -51.87597, -51.90547, -51.93516, 
        -51.96505, -51.995, -52.02465, -52.05376, -52.08211, -52.10972, 
        -52.13672, -52.16339, -52.18999, -52.21571, -52.24276, -52.27036, 
        -52.29873, -52.32798, -52.35814, -52.38902, -52.42043, -52.45226, 
        -52.48466, -52.51797, -52.55237, -52.58765, -52.62308, -52.65767, 
        -52.69052, -52.72113, -52.74949, -52.77607, -52.80146, -52.8262, 
        -52.85052, -52.87452, -52.89805, -52.91998, -52.94207, -52.96319, 
        -52.98317, -53.0019, -53.01942, -53.03576, -53.05109, -53.06561, 
        -53.07949, -53.09295, -53.10601, -53.11866, -53.13086, -53.14273, 
        -53.15474, -53.16725, -53.18034, -53.1936, -53.20633, -53.21787, 
        -53.22766, -53.23545, -53.2412, -53.24522, -53.24818, -53.24955, 
        -53.25145, -53.25236, -53.25159, -53.24869, -53.2433, -53.23522, 
        -53.22429, -53.21054, -53.19444, -53.17669, -53.15807, -53.13917, 
        -53.12047, -53.10246, -53.08526, -53.06886, -53.05284, -53.03648, 
        -53.01906, -52.99973, -52.97802, -52.95366, -52.92662, -52.89714, 
        -52.86537, -52.83171, -52.79651, -52.76015, -52.72303, -52.68529, 
        -52.64602, -52.60709, -52.56752, -52.52758, -52.48745, -52.44722, 
        -52.40674, -52.3658, -52.32433, -52.28239, -52.24018, -52.19769, 
        -52.15487, -52.11184, -52.06876, -52.026, -51.98373, -51.94201, 
        -51.90096, -51.86063, -51.82122, -51.78273, -51.74504, -51.70802, 
        -51.67154, -51.63551, -51.59978, -51.56408, -51.52821, -51.49184, 
        -51.45471, -51.41665, -51.37763, -51.33791, -51.29771, -51.25728, 
        -51.21562, -51.17474, -51.13371, -51.0927, -51.05209, -51.01223, 
        -50.97351, -50.93638, -50.9011, -50.86789, -50.83682, -50.80779, 
        -50.78055, -50.75471, -50.72987, -50.70541, -50.6808, -50.65581, 
        -50.6306, -50.60572, -50.58177, -50.55923, -50.53846, -50.51968, 
        -50.50323, -50.48935, -50.4781, -50.46941, -50.46301, -50.45851, 
        -50.4555, -50.4534, -50.45156, -50.44936, -50.44664, -50.44372, 
        -50.44102,
  -48.36154, -48.46762, -48.56858, -48.66368, -48.75213, -48.83358, 
        -48.9082, -48.97605, -49.03753, -49.09324, -49.14383, -49.18992, 
        -49.23211, -49.27063, -49.30461, -49.33608, -49.36389, -49.38829, 
        -49.41005, -49.43031, -49.45028, -49.47099, -49.49327, -49.51689, 
        -49.54229, -49.56865, -49.59608, -49.62392, -49.65139, -49.67807, 
        -49.70234, -49.72639, -49.74968, -49.77296, -49.79681, -49.82182, 
        -49.84831, -49.87586, -49.90406, -49.93188, -49.95881, -49.98372, 
        -50.00663, -50.02721, -50.0456, -50.06252, -50.07777, -50.09454, 
        -50.11242, -50.13162, -50.15166, -50.1723, -50.19265, -50.21231, 
        -50.23148, -50.25032, -50.26909, -50.28835, -50.30862, -50.3302, 
        -50.3532, -50.37727, -50.40105, -50.426, -50.45045, -50.47359, 
        -50.49452, -50.51255, -50.52745, -50.53947, -50.5492, -50.5573, 
        -50.56416, -50.56997, -50.57468, -50.57827, -50.58084, -50.58338, 
        -50.58579, -50.58915, -50.59293, -50.59937, -50.60851, -50.62071, 
        -50.63643, -50.65569, -50.67793, -50.70236, -50.72812, -50.75455, 
        -50.78121, -50.80804, -50.83514, -50.86259, -50.89053, -50.91886, 
        -50.94741, -50.97625, -51.00385, -51.03227, -51.06028, -51.08826, 
        -51.11613, -51.14395, -51.17141, -51.19831, -51.22448, -51.2499, 
        -51.27472, -51.29917, -51.32316, -51.34727, -51.37218, -51.39847, 
        -51.42612, -51.45476, -51.48367, -51.51242, -51.53971, -51.56725, 
        -51.59398, -51.62056, -51.64679, -51.67313, -51.70005, -51.72773, 
        -51.75621, -51.78532, -51.8151, -51.8456, -51.87679, -51.90859, 
        -51.94067, -51.97272, -52.00461, -52.03632, -52.06794, -52.09966, 
        -52.1314, -52.1621, -52.19345, -52.22419, -52.25404, -52.28305, 
        -52.31117, -52.33858, -52.36576, -52.39272, -52.41978, -52.44733, 
        -52.47566, -52.50494, -52.53518, -52.56613, -52.59761, -52.62959, 
        -52.66255, -52.69695, -52.73286, -52.76984, -52.80679, -52.84301, 
        -52.87651, -52.9088, -52.93899, -52.9675, -52.99509, -53.02201, 
        -53.04843, -53.07421, -53.09902, -53.12271, -53.14501, -53.1659, 
        -53.18549, -53.2036, -53.22029, -53.23569, -53.25009, -53.26386, 
        -53.27726, -53.29046, -53.30339, -53.31582, -53.32789, -53.33991, 
        -53.35224, -53.36413, -53.37764, -53.39145, -53.4049, -53.41729, 
        -53.4279, -53.43655, -53.4428, -53.44728, -53.45028, -53.45237, 
        -53.45367, -53.4539, -53.4524, -53.44882, -53.44272, -53.43388, 
        -53.4221, -53.40768, -53.39084, -53.37258, -53.35355, -53.33448, 
        -53.31572, -53.29738, -53.2795, -53.26194, -53.24438, -53.22619, 
        -53.2058, -53.18456, -53.16114, -53.13538, -53.10707, -53.07654, 
        -53.04371, -53.00905, -52.97298, -52.9358, -52.89779, -52.85896, 
        -52.81945, -52.77914, -52.738, -52.69633, -52.65455, -52.61235, 
        -52.57025, -52.52783, -52.48493, -52.44156, -52.39793, -52.35415, 
        -52.31029, -52.26646, -52.2229, -52.18006, -52.13803, -52.09679, 
        -52.0563, -52.01639, -51.97723, -51.93871, -51.89948, -51.86154, 
        -51.82367, -51.78564, -51.74751, -51.7092, -51.67059, -51.63163, 
        -51.59207, -51.552, -51.51137, -51.47025, -51.42874, -51.38697, 
        -51.34492, -51.30249, -51.25986, -51.21725, -51.17514, -51.13388, 
        -51.09373, -51.055, -51.01791, -50.98273, -50.9496, -50.91843, 
        -50.88905, -50.8611, -50.8341, -50.8074, -50.78041, -50.75291, 
        -50.72512, -50.6977, -50.67149, -50.64713, -50.62508, -50.60557, 
        -50.58881, -50.57511, -50.56436, -50.55641, -50.55085, -50.54619, 
        -50.54388, -50.54235, -50.541, -50.53944, -50.53786, -50.53659, 
        -50.53623,
  -48.3257, -48.43881, -48.546, -48.64597, -48.73829, -48.82272, 
        -48.89963, -48.96913, -49.03165, -49.08727, -49.13844, -49.18509, 
        -49.22787, -49.26706, -49.30301, -49.33582, -49.36583, -49.39308, 
        -49.4184, -49.44284, -49.46743, -49.4932, -49.52044, -49.54903, 
        -49.57785, -49.60863, -49.63978, -49.6711, -49.70166, -49.73088, 
        -49.75847, -49.78432, -49.80915, -49.83346, -49.85813, -49.88377, 
        -49.91072, -49.93878, -49.96739, -49.99598, -50.02268, -50.04871, 
        -50.07257, -50.09387, -50.11287, -50.13027, -50.14694, -50.16381, 
        -50.18198, -50.20157, -50.22232, -50.2436, -50.26488, -50.28576, 
        -50.30616, -50.32604, -50.3448, -50.36491, -50.38579, -50.40784, 
        -50.43116, -50.45561, -50.48086, -50.50657, -50.53176, -50.5561, 
        -50.57872, -50.59863, -50.61583, -50.63041, -50.64265, -50.65304, 
        -50.66187, -50.66817, -50.674, -50.67834, -50.68137, -50.68377, 
        -50.68614, -50.68929, -50.69388, -50.70039, -50.70989, -50.72281, 
        -50.73963, -50.76009, -50.78346, -50.80888, -50.83546, -50.86261, 
        -50.8899, -50.91619, -50.94363, -50.97134, -50.99957, -51.02826, 
        -51.05708, -51.08629, -51.11566, -51.14526, -51.17495, -51.20486, 
        -51.23508, -51.26527, -51.29511, -51.32408, -51.35201, -51.37894, 
        -51.40536, -51.43127, -51.45687, -51.48172, -51.50851, -51.53667, 
        -51.56618, -51.59657, -51.62725, -51.65759, -51.68719, -51.71625, 
        -51.7445, -51.7721, -51.79942, -51.82603, -51.85315, -51.8807, 
        -51.90908, -51.93783, -51.96778, -51.99865, -52.03074, -52.06277, 
        -52.09646, -52.13041, -52.1644, -52.19831, -52.23212, -52.26606, 
        -52.29994, -52.33376, -52.36701, -52.39961, -52.43106, -52.46169, 
        -52.49081, -52.5192, -52.54691, -52.57423, -52.60151, -52.62911, 
        -52.65746, -52.68681, -52.71714, -52.7472, -52.7789, -52.81145, 
        -52.84513, -52.88058, -52.91787, -52.95626, -52.99422, -53.03153, 
        -53.0673, -53.10113, -53.13317, -53.1638, -53.19358, -53.22282, 
        -53.25146, -53.27929, -53.30579, -53.33071, -53.3537, -53.37488, 
        -53.39441, -53.41222, -53.42837, -53.44313, -53.45589, -53.46914, 
        -53.48216, -53.49502, -53.50762, -53.51989, -53.53197, -53.54403, 
        -53.55642, -53.56944, -53.58311, -53.59715, -53.61092, -53.62379, 
        -53.63517, -53.64456, -53.65174, -53.6568, -53.66011, -53.66229, 
        -53.6632, -53.66286, -53.66065, -53.65617, -53.64924, -53.63965, 
        -53.62729, -53.61119, -53.5939, -53.57524, -53.55593, -53.5367, 
        -53.51758, -53.49865, -53.47979, -53.46083, -53.44159, -53.42149, 
        -53.40009, -53.37694, -53.35174, -53.32473, -53.29514, -53.26359, 
        -53.2297, -53.19424, -53.15763, -53.11975, -53.08083, -53.04103, 
        -53.00021, -52.95839, -52.9155, -52.87186, -52.82794, -52.78385, 
        -52.73989, -52.69599, -52.65157, -52.60583, -52.561, -52.51633, 
        -52.47165, -52.42717, -52.38319, -52.34042, -52.29882, -52.25804, 
        -52.21788, -52.17823, -52.13905, -52.1002, -52.06127, -52.02199, 
        -51.98227, -51.94206, -51.90146, -51.86066, -51.81931, -51.778, 
        -51.73625, -51.69421, -51.65203, -51.60942, -51.56657, -51.5235, 
        -51.48019, -51.4365, -51.39253, -51.34859, -51.30531, -51.26289, 
        -51.22146, -51.18134, -51.14268, -51.10571, -51.07061, -51.03727, 
        -51.00458, -50.97417, -50.94458, -50.91535, -50.88569, -50.85559, 
        -50.82537, -50.79573, -50.76763, -50.74178, -50.71869, -50.69851, 
        -50.68128, -50.6673, -50.65638, -50.64824, -50.64247, -50.63857, 
        -50.63583, -50.63394, -50.63248, -50.63124, -50.63057, -50.63097, 
        -50.63281,
  -48.28697, -48.4079, -48.52179, -48.62751, -48.72338, -48.81132, 
        -48.89043, -48.96143, -49.02479, -49.08157, -49.13232, -49.17812, 
        -49.22003, -49.2586, -49.29455, -49.32803, -49.35978, -49.3901, 
        -49.41975, -49.44833, -49.47873, -49.51059, -49.54392, -49.57836, 
        -49.61341, -49.64886, -49.6845, -49.71951, -49.7534, -49.78556, 
        -49.81578, -49.84406, -49.8709, -49.89683, -49.92181, -49.94827, 
        -49.97565, -50.00423, -50.03333, -50.06279, -50.09139, -50.11843, 
        -50.14326, -50.16555, -50.1851, -50.20297, -50.22016, -50.2375, 
        -50.25598, -50.27579, -50.29582, -50.31761, -50.3395, -50.36125, 
        -50.38259, -50.40345, -50.42417, -50.44525, -50.46691, -50.48959, 
        -50.51356, -50.5386, -50.56444, -50.59068, -50.61676, -50.64208, 
        -50.66596, -50.6866, -50.70598, -50.72305, -50.73795, -50.75089, 
        -50.76198, -50.77119, -50.77867, -50.78429, -50.78832, -50.79129, 
        -50.79386, -50.79692, -50.80128, -50.80773, -50.81737, -50.8308, 
        -50.84836, -50.86857, -50.89267, -50.91867, -50.9457, -50.97328, 
        -51.00094, -51.02866, -51.05651, -51.08463, -51.11325, -51.14226, 
        -51.17175, -51.20147, -51.23169, -51.26248, -51.29368, -51.32547, 
        -51.35776, -51.38902, -51.42083, -51.45155, -51.48096, -51.50937, 
        -51.53721, -51.56482, -51.59224, -51.62017, -51.64925, -51.67971, 
        -51.71157, -51.74414, -51.77659, -51.80875, -51.84034, -51.87123, 
        -51.90111, -51.93011, -51.95827, -51.98471, -52.01216, -52.03913, 
        -52.06672, -52.09515, -52.12489, -52.15592, -52.18866, -52.22254, 
        -52.25746, -52.29289, -52.32864, -52.36448, -52.40047, -52.43661, 
        -52.4728, -52.50874, -52.54412, -52.57874, -52.6119, -52.64387, 
        -52.67463, -52.70311, -52.73137, -52.75926, -52.78686, -52.81463, 
        -52.84309, -52.87258, -52.90311, -52.93441, -52.96655, -52.99982, 
        -53.03446, -53.07121, -53.10946, -53.14868, -53.18777, -53.22575, 
        -53.26245, -53.29762, -53.33138, -53.36405, -53.39605, -53.42756, 
        -53.45755, -53.48755, -53.51601, -53.54243, -53.56665, -53.5886, 
        -53.60847, -53.62634, -53.64243, -53.65686, -53.67025, -53.68332, 
        -53.69614, -53.70898, -53.72137, -53.73342, -53.74539, -53.75743, 
        -53.76984, -53.78284, -53.79642, -53.8104, -53.82421, -53.83737, 
        -53.84937, -53.85955, -53.86768, -53.87255, -53.87648, -53.87874, 
        -53.87937, -53.87826, -53.87519, -53.8698, -53.86205, -53.85174, 
        -53.83889, -53.82346, -53.80603, -53.78704, -53.76755, -53.74811, 
        -53.72839, -53.70859, -53.68855, -53.66796, -53.64682, -53.62469, 
        -53.60124, -53.5763, -53.54963, -53.52119, -53.49059, -53.45787, 
        -53.42319, -53.38689, -53.34846, -53.3099, -53.27028, -53.22942, 
        -53.18722, -53.14376, -53.09898, -53.0533, -53.00726, -52.96121, 
        -52.91539, -52.86951, -52.82376, -52.77792, -52.73215, -52.68658, 
        -52.64134, -52.59631, -52.55238, -52.50955, -52.46796, -52.42759, 
        -52.38787, -52.34827, -52.30883, -52.26928, -52.22911, -52.18809, 
        -52.1462, -52.10359, -52.06055, -52.01715, -51.97355, -51.9299, 
        -51.88607, -51.84261, -51.79782, -51.7538, -51.70955, -51.66515, 
        -51.62066, -51.57576, -51.53052, -51.48553, -51.44114, -51.39775, 
        -51.35538, -51.31414, -51.27418, -51.23565, -51.19865, -51.1632, 
        -51.1291, -51.09621, -51.06377, -51.03173, -50.99958, -50.96699, 
        -50.93475, -50.90317, -50.87355, -50.8465, -50.82251, -50.80165, 
        -50.78398, -50.76937, -50.75767, -50.74856, -50.74165, -50.73642, 
        -50.73241, -50.72934, -50.72701, -50.72555, -50.72545, -50.72725, 
        -50.73109,
  -48.24429, -48.37439, -48.49574, -48.60764, -48.70931, -48.80083, 
        -48.88244, -48.95459, -49.01793, -49.07368, -49.12246, -49.16607, 
        -49.20554, -49.24116, -49.27587, -49.30954, -49.34276, -49.37651, 
        -49.41117, -49.44721, -49.48491, -49.52425, -49.5651, -49.60633, 
        -49.64768, -49.68881, -49.72893, -49.76793, -49.80434, -49.83981, 
        -49.87309, -49.90422, -49.93354, -49.96165, -49.98933, -50.01713, 
        -50.04533, -50.07458, -50.1043, -50.13449, -50.16403, -50.19201, 
        -50.21796, -50.2411, -50.2607, -50.27917, -50.29682, -50.31496, 
        -50.33381, -50.35385, -50.37489, -50.39682, -50.41916, -50.44152, 
        -50.46354, -50.48546, -50.50721, -50.52917, -50.55181, -50.57539, 
        -50.60004, -50.62471, -50.65105, -50.6778, -50.7043, -50.73045, 
        -50.75515, -50.77817, -50.79944, -50.81887, -50.83646, -50.85205, 
        -50.86577, -50.8773, -50.88687, -50.89444, -50.90018, -50.90441, 
        -50.90675, -50.91005, -50.91436, -50.92089, -50.93064, -50.94436, 
        -50.9622, -50.98371, -51.008, -51.03402, -51.06096, -51.08841, 
        -51.11614, -51.14408, -51.17231, -51.201, -51.2302, -51.25991, 
        -51.28922, -51.31994, -51.35142, -51.3834, -51.4161, -51.44981, 
        -51.48404, -51.51816, -51.55161, -51.58393, -51.61504, -51.64513, 
        -51.67453, -51.70366, -51.73307, -51.76336, -51.79496, -51.82806, 
        -51.86234, -51.89718, -51.93087, -51.96516, -51.99874, -52.03149, 
        -52.06325, -52.09372, -52.12305, -52.15107, -52.1779, -52.20503, 
        -52.23186, -52.25969, -52.28884, -52.31985, -52.35288, -52.3876, 
        -52.42348, -52.4601, -52.4972, -52.53474, -52.57268, -52.60991, 
        -52.64832, -52.68642, -52.72377, -52.76035, -52.79538, -52.82885, 
        -52.86079, -52.89128, -52.92078, -52.94941, -52.97761, -53.00583, 
        -53.03456, -53.06421, -53.09499, -53.12679, -53.15965, -53.19373, 
        -53.22958, -53.26735, -53.30686, -53.34679, -53.38527, -53.42381, 
        -53.46119, -53.49754, -53.53292, -53.56751, -53.60162, -53.63535, 
        -53.66855, -53.70074, -53.73121, -53.75973, -53.78557, -53.80864, 
        -53.82882, -53.84736, -53.86354, -53.878, -53.89139, -53.90461, 
        -53.91781, -53.93081, -53.94342, -53.95559, -53.96761, -53.97878, 
        -53.99114, -54.00402, -54.01739, -54.03091, -54.04457, -54.05791, 
        -54.07033, -54.08125, -54.09022, -54.09698, -54.10149, -54.10375, 
        -54.10383, -54.1017, -54.09744, -54.0912, -54.08262, -54.07179, 
        -54.05871, -54.04334, -54.02601, -54.00726, -53.9877, -53.96766, 
        -53.94737, -53.92657, -53.9051, -53.88179, -53.85858, -53.8343, 
        -53.80889, -53.7822, -53.75412, -53.7244, -53.69279, -53.65907, 
        -53.6233, -53.58582, -53.54738, -53.50799, -53.46762, -53.42587, 
        -53.38248, -53.33741, -53.29087, -53.24324, -53.19516, -53.14708, 
        -53.09918, -53.05162, -53.00436, -52.95745, -52.91083, -52.86462, 
        -52.81886, -52.77368, -52.72943, -52.68647, -52.64499, -52.60492, 
        -52.56432, -52.52441, -52.48433, -52.44352, -52.4017, -52.3585, 
        -52.31421, -52.26909, -52.2235, -52.17777, -52.13219, -52.08697, 
        -52.04161, -51.99658, -51.95126, -51.90588, -51.86019, -51.81442, 
        -51.7685, -51.72232, -51.67599, -51.62988, -51.5845, -51.54025, 
        -51.49723, -51.45528, -51.41438, -51.37459, -51.33599, -51.29861, 
        -51.26217, -51.22644, -51.19117, -51.15615, -51.1212, -51.08626, 
        -51.05225, -51.01934, -50.98869, -50.96077, -50.93601, -50.9146, 
        -50.89531, -50.87976, -50.86688, -50.85633, -50.8477, -50.84055, 
        -50.83454, -50.82958, -50.82579, -50.82364, -50.82372, -50.82646, 
        -50.83178,
  -48.20109, -48.3407, -48.47003, -48.58858, -48.69539, -48.7904, 
        -48.87419, -48.94704, -49.00829, -49.06166, -49.10696, -49.14619, 
        -49.18142, -49.21432, -49.24661, -49.27968, -49.3146, -49.35227, 
        -49.39316, -49.43726, -49.48418, -49.53312, -49.58274, -49.63166, 
        -49.68019, -49.72733, -49.77249, -49.81568, -49.85675, -49.89555, 
        -49.93192, -49.96621, -49.99858, -50.0295, -50.05944, -50.08917, 
        -50.11896, -50.14911, -50.1786, -50.20934, -50.23947, -50.2683, 
        -50.29493, -50.31925, -50.34119, -50.36076, -50.37957, -50.39847, 
        -50.41793, -50.43817, -50.45938, -50.48146, -50.50395, -50.52673, 
        -50.54944, -50.57115, -50.59393, -50.61699, -50.64058, -50.6649, 
        -50.69004, -50.71597, -50.74251, -50.76936, -50.79608, -50.82238, 
        -50.84781, -50.87211, -50.89518, -50.91692, -50.93714, -50.95557, 
        -50.97116, -50.98544, -50.99763, -51.00749, -51.01526, -51.02122, 
        -51.02586, -51.03008, -51.03505, -51.04206, -51.05225, -51.0661, 
        -51.08386, -51.10505, -51.12883, -51.15416, -51.18037, -51.20712, 
        -51.23336, -51.26116, -51.28962, -51.3188, -51.34884, -51.37973, 
        -51.4114, -51.4437, -51.47658, -51.51016, -51.54467, -51.58025, 
        -51.61627, -51.65231, -51.68748, -51.7216, -51.75459, -51.78658, 
        -51.81778, -51.84776, -51.87912, -51.91158, -51.94561, -51.98119, 
        -52.01796, -52.05525, -52.09244, -52.12907, -52.16479, -52.19938, 
        -52.23264, -52.26434, -52.29435, -52.32265, -52.3497, -52.37622, 
        -52.40271, -52.42995, -52.45882, -52.48887, -52.52226, -52.55767, 
        -52.59449, -52.63219, -52.67051, -52.70938, -52.7488, -52.78863, 
        -52.82866, -52.8683, -52.9074, -52.9456, -52.98225, -53.01724, 
        -53.0507, -53.08279, -53.11362, -53.14341, -53.17258, -53.20161, 
        -53.23084, -53.25996, -53.29121, -53.32363, -53.35727, -53.39223, 
        -53.42898, -53.46774, -53.50795, -53.54856, -53.58866, -53.62782, 
        -53.66626, -53.70377, -53.74069, -53.77696, -53.81285, -53.84843, 
        -53.88362, -53.91774, -53.95012, -53.98024, -54.0077, -54.03185, 
        -54.05339, -54.07114, -54.08803, -54.10305, -54.11724, -54.13114, 
        -54.14504, -54.15882, -54.17216, -54.18501, -54.19746, -54.20982, 
        -54.22233, -54.2351, -54.24823, -54.26137, -54.27486, -54.2883, 
        -54.30118, -54.31277, -54.32243, -54.32972, -54.33447, -54.33644, 
        -54.33574, -54.33245, -54.32693, -54.31941, -54.3089, -54.29764, 
        -54.28459, -54.26932, -54.25233, -54.23392, -54.21451, -54.19418, 
        -54.17319, -54.15137, -54.12859, -54.10455, -54.07928, -54.05277, 
        -54.02513, -53.99648, -53.9667, -53.93546, -53.90263, -53.86792, 
        -53.83128, -53.79303, -53.75356, -53.71331, -53.67212, -53.62947, 
        -53.585, -53.53851, -53.49033, -53.44089, -53.391, -53.33991, 
        -53.29004, -53.24079, -53.19217, -53.1442, -53.09701, -53.05044, 
        -53.00452, -52.95932, -52.91505, -52.87196, -52.83013, -52.7896, 
        -52.7494, -52.70887, -52.66768, -52.62524, -52.58129, -52.53611, 
        -52.48967, -52.44236, -52.39453, -52.34675, -52.29947, -52.25265, 
        -52.20597, -52.15923, -52.11235, -52.06527, -52.01806, -51.97078, 
        -51.9234, -51.87606, -51.8287, -51.78174, -51.73559, -51.69061, 
        -51.64676, -51.60318, -51.56147, -51.5206, -51.48029, -51.44071, 
        -51.40189, -51.36332, -51.32493, -51.287, -51.24951, -51.2127, 
        -51.17709, -51.14326, -51.11193, -51.08355, -51.05841, -51.03649, 
        -51.01756, -51.00111, -50.98692, -50.97466, -50.96396, -50.95441, 
        -50.94603, -50.93881, -50.93327, -50.92999, -50.92964, -50.93258, 
        -50.93859,
  -48.15976, -48.30864, -48.44465, -48.56899, -48.68033, -48.77814, 
        -48.86285, -48.93507, -48.99521, -49.04447, -49.08459, -49.11775, 
        -49.14682, -49.17454, -49.20329, -49.23537, -49.27237, -49.31401, 
        -49.36269, -49.4168, -49.47504, -49.53539, -49.59618, -49.65589, 
        -49.7129, -49.76671, -49.81726, -49.86475, -49.90936, -49.95145, 
        -49.99107, -50.02869, -50.06355, -50.09784, -50.1309, -50.16309, 
        -50.19483, -50.22639, -50.25786, -50.28914, -50.31974, -50.34924, 
        -50.37677, -50.40228, -50.42555, -50.44687, -50.4672, -50.48738, 
        -50.50657, -50.52716, -50.54853, -50.57064, -50.59328, -50.61646, 
        -50.63983, -50.66331, -50.6869, -50.71095, -50.73539, -50.76032, 
        -50.78574, -50.81166, -50.838, -50.86462, -50.89122, -50.9166, 
        -50.94255, -50.96795, -50.99267, -51.01657, -51.03933, -51.0606, 
        -51.08006, -51.09738, -51.11232, -51.12477, -51.13508, -51.14328, 
        -51.14992, -51.15578, -51.16208, -51.1701, -51.18092, -51.19399, 
        -51.21149, -51.23187, -51.25446, -51.27846, -51.30337, -51.32896, 
        -51.35531, -51.38264, -51.41112, -51.44084, -51.47195, -51.50423, 
        -51.53758, -51.57178, -51.60677, -51.64233, -51.67864, -51.71605, 
        -51.75304, -51.79097, -51.82814, -51.86422, -51.89924, -51.93325, 
        -51.9665, -51.9994, -52.03276, -52.06736, -52.10389, -52.14208, 
        -52.1814, -52.22126, -52.26102, -52.3001, -52.33807, -52.37443, 
        -52.40896, -52.44047, -52.47089, -52.49924, -52.52631, -52.55275, 
        -52.57899, -52.60617, -52.63514, -52.66643, -52.70022, -52.7362, 
        -52.77375, -52.81228, -52.85149, -52.89134, -52.93167, -52.97247, 
        -53.0135, -53.05429, -53.09459, -53.13403, -53.17219, -53.20784, 
        -53.24298, -53.27679, -53.30933, -53.34073, -53.37122, -53.40128, 
        -53.43138, -53.46224, -53.49425, -53.52752, -53.56209, -53.5981, 
        -53.63587, -53.67521, -53.71589, -53.7569, -53.79746, -53.8373, 
        -53.8766, -53.91527, -53.95354, -53.99123, -54.02759, -54.06482, 
        -54.10155, -54.13728, -54.17134, -54.20301, -54.23177, -54.25747, 
        -54.27995, -54.29987, -54.31777, -54.33404, -54.34949, -54.36459, 
        -54.37969, -54.39469, -54.40936, -54.42339, -54.43683, -54.44986, 
        -54.46273, -54.47557, -54.48843, -54.5015, -54.51502, -54.52838, 
        -54.54051, -54.55259, -54.56268, -54.56999, -54.57442, -54.57565, 
        -54.57358, -54.56868, -54.56184, -54.55307, -54.54283, -54.53139, 
        -54.51826, -54.50341, -54.48692, -54.46898, -54.44976, -54.4293, 
        -54.4077, -54.38494, -54.36077, -54.33536, -54.30831, -54.27969, 
        -54.24992, -54.2192, -54.1876, -54.15488, -54.12073, -54.08389, 
        -54.04622, -54.00697, -53.9664, -53.9251, -53.88305, -53.8395, 
        -53.79408, -53.74633, -53.69666, -53.64566, -53.59396, -53.54213, 
        -53.49068, -53.43974, -53.38969, -53.34075, -53.29284, -53.24603, 
        -53.20005, -53.15501, -53.11075, -53.06742, -53.02507, -52.98354, 
        -52.94222, -52.90041, -52.85743, -52.81298, -52.76688, -52.71932, 
        -52.67087, -52.6217, -52.57242, -52.52325, -52.47354, -52.42519, 
        -52.37706, -52.32869, -52.28008, -52.23127, -52.18228, -52.1334, 
        -52.08463, -52.03602, -51.98773, -51.94004, -51.89333, -51.84779, 
        -51.80344, -51.76027, -51.71781, -51.67588, -51.63425, -51.59249, 
        -51.55095, -51.50966, -51.46833, -51.42758, -51.38767, -51.34907, 
        -51.31227, -51.27778, -51.24601, -51.21742, -51.19198, -51.16955, 
        -51.14973, -51.13237, -51.1168, -51.10276, -51.08989, -51.07796, 
        -51.06697, -51.05737, -51.0499, -51.0453, -51.0442, -51.04675, 
        -51.05272,
  -48.12417, -48.2801, -48.42332, -48.55219, -48.66605, -48.76498, 
        -48.8491, -48.91879, -48.97484, -49.01845, -49.05162, -49.07706, 
        -49.0976, -49.11885, -49.14342, -49.17451, -49.21427, -49.26341, 
        -49.32185, -49.38807, -49.45974, -49.53383, -49.60743, -49.67823, 
        -49.74471, -49.80606, -49.86231, -49.91317, -49.96135, -50.00653, 
        -50.04933, -50.09034, -50.1299, -50.16799, -50.20472, -50.24015, 
        -50.27439, -50.30783, -50.34053, -50.37245, -50.4035, -50.43345, 
        -50.46201, -50.48785, -50.51285, -50.53622, -50.55844, -50.58004, 
        -50.60135, -50.62271, -50.64437, -50.66672, -50.68981, -50.71335, 
        -50.73719, -50.76137, -50.78581, -50.81045, -50.8355, -50.85977, 
        -50.88521, -50.9109, -50.93689, -50.96307, -50.98935, -51.01586, 
        -51.04229, -51.06866, -51.09493, -51.12074, -51.14575, -51.16964, 
        -51.19188, -51.21204, -51.22992, -51.24525, -51.25715, -51.26798, 
        -51.2771, -51.28534, -51.29369, -51.30335, -51.31517, -51.32965, 
        -51.34677, -51.36608, -51.3871, -51.40934, -51.43254, -51.45667, 
        -51.48192, -51.50855, -51.53681, -51.56706, -51.59921, -51.6319, 
        -51.66708, -51.70337, -51.74045, -51.77829, -51.81689, -51.85632, 
        -51.89627, -51.9362, -51.97555, -52.01391, -52.0512, -52.08742, 
        -52.12282, -52.15787, -52.19338, -52.23027, -52.26926, -52.31009, 
        -52.35116, -52.39365, -52.4359, -52.47735, -52.51739, -52.5554, 
        -52.59085, -52.62393, -52.65453, -52.6832, -52.71045, -52.73686, 
        -52.76322, -52.79087, -52.82034, -52.85225, -52.8866, -52.92306, 
        -52.96107, -53.0001, -53.03982, -53.07904, -53.11974, -53.16079, 
        -53.20222, -53.24358, -53.28451, -53.32514, -53.36465, -53.40294, 
        -53.43991, -53.47562, -53.51005, -53.54328, -53.57539, -53.60681, 
        -53.63818, -53.67019, -53.70334, -53.73785, -53.77361, -53.81075, 
        -53.84929, -53.88821, -53.92905, -53.97018, -54.01113, -54.0516, 
        -54.09168, -54.1314, -54.17075, -54.20963, -54.2482, -54.28647, 
        -54.3243, -54.36124, -54.39655, -54.42947, -54.45948, -54.48649, 
        -54.51052, -54.53196, -54.55135, -54.56934, -54.58656, -54.60349, 
        -54.6203, -54.63699, -54.65234, -54.66805, -54.68301, -54.69716, 
        -54.71103, -54.72449, -54.73712, -54.75031, -54.7641, -54.77742, 
        -54.79051, -54.80243, -54.81244, -54.81958, -54.82315, -54.82313, 
        -54.81963, -54.81318, -54.80455, -54.79441, -54.78352, -54.77161, 
        -54.75847, -54.74419, -54.72831, -54.71082, -54.6919, -54.67139, 
        -54.64833, -54.62482, -54.5998, -54.57312, -54.54464, -54.51441, 
        -54.48275, -54.45004, -54.41654, -54.38211, -54.34634, -54.30934, 
        -54.27061, -54.23039, -54.18901, -54.14665, -54.10332, -54.05845, 
        -54.01192, -53.96295, -53.91215, -53.85992, -53.8068, -53.75348, 
        -53.70055, -53.64816, -53.59673, -53.5467, -53.49817, -53.45108, 
        -53.40512, -53.36007, -53.31578, -53.27095, -53.22771, -53.1848, 
        -53.14172, -53.09786, -53.05272, -53.00589, -52.95754, -52.90792, 
        -52.85756, -52.80694, -52.75632, -52.70603, -52.65611, -52.60646, 
        -52.55686, -52.50705, -52.45668, -52.40608, -52.35538, -52.30488, 
        -52.25462, -52.20482, -52.15574, -52.10754, -52.06041, -52.01451, 
        -51.96973, -51.92587, -51.88261, -51.83956, -51.79639, -51.75263, 
        -51.7086, -51.66452, -51.62055, -51.57732, -51.53532, -51.49512, 
        -51.45732, -51.42128, -51.38931, -51.36043, -51.33464, -51.31151, 
        -51.29117, -51.27261, -51.25565, -51.23975, -51.22472, -51.21038, 
        -51.1969, -51.18503, -51.17573, -51.16974, -51.16761, -51.16941, 
        -51.17472,
  -48.10087, -48.26063, -48.4067, -48.53732, -48.65142, -48.74901, 
        -48.8293, -48.89441, -48.94417, -48.98013, -49.0047, -49.02118, 
        -49.03399, -49.04847, -49.06882, -49.09948, -49.143, -49.20046, 
        -49.27057, -49.35113, -49.43851, -49.52719, -49.61512, -49.69838, 
        -49.77505, -49.84451, -49.90688, -49.9632, -50.0148, -50.06298, 
        -50.10886, -50.15321, -50.19656, -50.23881, -50.27964, -50.31881, 
        -50.35624, -50.3909, -50.42506, -50.45772, -50.4893, -50.51986, 
        -50.54939, -50.57772, -50.6048, -50.63044, -50.65487, -50.67826, 
        -50.7011, -50.72343, -50.74596, -50.76884, -50.79239, -50.81538, 
        -50.8398, -50.86442, -50.88939, -50.91456, -50.9398, -50.96517, 
        -50.99053, -51.01603, -51.04168, -51.06742, -51.09364, -51.12024, 
        -51.14717, -51.17448, -51.20189, -51.22905, -51.25498, -51.28109, 
        -51.30573, -51.32854, -51.34918, -51.3674, -51.38313, -51.3967, 
        -51.40878, -51.41981, -51.43093, -51.44287, -51.45623, -51.47148, 
        -51.48838, -51.50668, -51.526, -51.54635, -51.56667, -51.58926, 
        -51.61337, -51.63927, -51.66733, -51.69791, -51.73061, -51.76569, 
        -51.80258, -51.84086, -51.8801, -51.92022, -51.96106, -52.00254, 
        -52.04456, -52.08656, -52.12827, -52.16929, -52.20922, -52.24699, 
        -52.28478, -52.3222, -52.3601, -52.39951, -52.44097, -52.48438, 
        -52.52915, -52.57425, -52.61897, -52.66256, -52.70433, -52.74361, 
        -52.77998, -52.8136, -52.8441, -52.87294, -52.90059, -52.92772, 
        -52.95526, -52.98248, -53.01283, -53.04557, -53.0806, -53.11745, 
        -53.1557, -53.1949, -53.23467, -53.27481, -53.31535, -53.35617, 
        -53.39748, -53.43886, -53.48045, -53.5216, -53.56245, -53.60232, 
        -53.64108, -53.67877, -53.71517, -53.7502, -53.78402, -53.81607, 
        -53.84903, -53.88256, -53.91721, -53.95321, -53.99047, -54.02885, 
        -54.0683, -54.1086, -54.14943, -54.19061, -54.23198, -54.27298, 
        -54.31384, -54.35439, -54.39457, -54.43434, -54.47371, -54.51269, 
        -54.5511, -54.58867, -54.62476, -54.65864, -54.68984, -54.71725, 
        -54.74302, -54.76646, -54.78801, -54.80822, -54.82763, -54.84668, 
        -54.86554, -54.88416, -54.90239, -54.92001, -54.93683, -54.95272, 
        -54.96782, -54.98183, -54.99528, -55.00902, -55.02285, -55.03631, 
        -55.04911, -55.06087, -55.0703, -55.07658, -55.07898, -55.07745, 
        -55.07228, -55.06322, -55.05323, -55.04209, -55.03022, -55.01782, 
        -55.00479, -54.99087, -54.97571, -54.95869, -54.93993, -54.91943, 
        -54.89686, -54.87275, -54.84702, -54.81948, -54.79005, -54.75877, 
        -54.7258, -54.69144, -54.65594, -54.61958, -54.58208, -54.54377, 
        -54.50389, -54.4629, -54.42075, -54.37728, -54.33252, -54.28622, 
        -54.23828, -54.18824, -54.13534, -54.0822, -54.02815, -53.97357, 
        -53.91943, -53.86574, -53.81309, -53.76193, -53.71252, -53.66483, 
        -53.61857, -53.57325, -53.52864, -53.48417, -53.43964, -53.39489, 
        -53.34953, -53.3032, -53.25552, -53.20636, -53.15583, -53.10425, 
        -53.05241, -53.00031, -52.9486, -52.89748, -52.84652, -52.79559, 
        -52.7445, -52.69301, -52.64111, -52.58908, -52.53669, -52.48452, 
        -52.43287, -52.38208, -52.33227, -52.28268, -52.2352, -52.18901, 
        -52.14371, -52.09909, -52.05482, -52.01045, -51.96555, -51.9199, 
        -51.87364, -51.82714, -51.78098, -51.73569, -51.69201, -51.65052, 
        -51.61173, -51.57599, -51.54346, -51.51415, -51.48801, -51.46445, 
        -51.44315, -51.42352, -51.40509, -51.38737, -51.37011, -51.35343, 
        -51.33765, -51.32383, -51.31293, -51.3057, -51.30247, -51.30328, 
        -51.30736,
  -48.09237, -48.25029, -48.39484, -48.52329, -48.63435, -48.72754, 
        -48.80302, -48.86128, -48.90269, -48.92929, -48.9437, -48.95028, 
        -48.95473, -48.96253, -48.9798, -49.01159, -49.05989, -49.12736, 
        -49.21131, -49.30829, -49.41286, -49.51933, -49.62275, -49.71912, 
        -49.80646, -49.88422, -49.95282, -50.01386, -50.06889, -50.12011, 
        -50.16904, -50.21588, -50.26305, -50.30951, -50.35463, -50.39768, 
        -50.4385, -50.47687, -50.51281, -50.54688, -50.5793, -50.61069, 
        -50.64132, -50.6712, -50.70029, -50.72829, -50.75521, -50.7798, 
        -50.8044, -50.82835, -50.85203, -50.87595, -50.90005, -50.92449, 
        -50.94928, -50.97437, -50.9995, -51.02486, -51.05024, -51.07558, 
        -51.101, -51.12651, -51.15199, -51.17772, -51.20287, -51.22961, 
        -51.25698, -51.2848, -51.31298, -51.34118, -51.36937, -51.39709, 
        -51.42364, -51.44866, -51.47173, -51.49276, -51.51146, -51.52814, 
        -51.54338, -51.55775, -51.57194, -51.5856, -51.60094, -51.61722, 
        -51.63425, -51.65186, -51.67007, -51.68889, -51.70871, -51.73001, 
        -51.75318, -51.77853, -51.80636, -51.83693, -51.8702, -51.90608, 
        -51.94415, -51.98378, -52.02456, -52.06649, -52.1084, -52.15211, 
        -52.19636, -52.2408, -52.28514, -52.32907, -52.37207, -52.41379, 
        -52.45437, -52.49446, -52.53508, -52.57715, -52.62116, -52.66703, 
        -52.71413, -52.76171, -52.80873, -52.85426, -52.89749, -52.93685, 
        -52.9742, -53.00834, -53.03969, -53.06927, -53.09761, -53.12553, 
        -53.15403, -53.18354, -53.21485, -53.24832, -53.28394, -53.32122, 
        -53.35968, -53.39881, -53.43831, -53.47808, -53.51827, -53.5588, 
        -53.59976, -53.64113, -53.68261, -53.72372, -53.7653, -53.80663, 
        -53.84705, -53.88639, -53.92442, -53.96106, -53.99648, -54.03117, 
        -54.0658, -54.10103, -54.13732, -54.17499, -54.21378, -54.25341, 
        -54.29387, -54.33477, -54.37597, -54.41752, -54.45918, -54.50084, 
        -54.54234, -54.58359, -54.62329, -54.66362, -54.70351, -54.74296, 
        -54.78172, -54.8196, -54.85628, -54.89098, -54.92326, -54.95308, 
        -54.98065, -55.00621, -55.03029, -55.05303, -55.07492, -55.09632, 
        -55.11736, -55.13805, -55.15837, -55.1779, -55.1965, -55.21425, 
        -55.23085, -55.24631, -55.26076, -55.27404, -55.2879, -55.30129, 
        -55.314, -55.32514, -55.33379, -55.33904, -55.34029, -55.33741, 
        -55.33082, -55.32149, -55.31036, -55.29838, -55.28597, -55.27333, 
        -55.2604, -55.24688, -55.23223, -55.21581, -55.1972, -55.17659, 
        -55.15376, -55.12922, -55.10299, -55.0747, -55.04444, -55.01228, 
        -54.9783, -54.94259, -54.90437, -54.86619, -54.82728, -54.78736, 
        -54.74683, -54.705, -54.66188, -54.61742, -54.5714, -54.52359, 
        -54.47393, -54.42252, -54.36945, -54.31556, -54.26059, -54.20513, 
        -54.14961, -54.09471, -54.04098, -53.98856, -53.93798, -53.88923, 
        -53.84204, -53.79588, -53.75032, -53.70457, -53.65822, -53.61152, 
        -53.56378, -53.51497, -53.46474, -53.41324, -53.3607, -53.30748, 
        -53.253, -53.19967, -53.14683, -53.09467, -53.04264, -52.99045, 
        -52.93807, -52.88535, -52.8321, -52.77856, -52.72483, -52.6713, 
        -52.61845, -52.56662, -52.51624, -52.46741, -52.41943, -52.37268, 
        -52.32676, -52.28131, -52.2359, -52.19012, -52.14353, -52.09606, 
        -52.04794, -51.99963, -51.9517, -51.90493, -51.86, -51.81736, 
        -51.7775, -51.74098, -51.7077, -51.67768, -51.65073, -51.62642, 
        -51.60414, -51.58327, -51.56328, -51.54367, -51.52432, -51.50553, 
        -51.48791, -51.47246, -51.46018, -51.45075, -51.44641, -51.44592, 
        -51.4486,
  -48.09911, -48.25195, -48.39016, -48.51178, -48.61594, -48.70153, 
        -48.76857, -48.81722, -48.84831, -48.86398, -48.86686, -48.86391, 
        -48.86029, -48.86316, -48.87925, -48.91405, -48.9711, -49.05073, 
        -49.15028, -49.26489, -49.38755, -49.51156, -49.6307, -49.74051, 
        -49.83875, -49.92376, -49.99859, -50.06433, -50.12304, -50.17735, 
        -50.22948, -50.28075, -50.33186, -50.38245, -50.43178, -50.47904, 
        -50.52338, -50.56476, -50.60309, -50.63886, -50.67265, -50.7042, 
        -50.73607, -50.76757, -50.79867, -50.82899, -50.85835, -50.88628, 
        -50.9131, -50.9389, -50.96421, -50.98927, -51.01425, -51.0394, 
        -51.06451, -51.0898, -51.1152, -51.1396, -51.16496, -51.19038, 
        -51.21603, -51.24155, -51.26724, -51.29321, -51.31957, -51.34656, 
        -51.37402, -51.40212, -51.43073, -51.45939, -51.48822, -51.51682, 
        -51.54473, -51.57149, -51.59676, -51.61916, -51.64077, -51.66067, 
        -51.67934, -51.69727, -51.71494, -51.73274, -51.75067, -51.76854, 
        -51.78631, -51.80395, -51.82162, -51.83969, -51.85865, -51.87913, 
        -51.90162, -51.92655, -51.95414, -51.98346, -52.01662, -52.05246, 
        -52.09085, -52.13119, -52.17314, -52.2162, -52.26096, -52.30684, 
        -52.35361, -52.40083, -52.44815, -52.49526, -52.54149, -52.58662, 
        -52.63042, -52.67348, -52.71697, -52.76178, -52.80737, -52.85556, 
        -52.90486, -52.95436, -53.00325, -53.05047, -53.09512, -53.13666, 
        -53.17489, -53.20995, -53.24236, -53.27283, -53.30224, -53.33145, 
        -53.36122, -53.39214, -53.4246, -53.45895, -53.49511, -53.53278, 
        -53.57137, -53.60953, -53.64882, -53.68821, -53.72784, -53.76792, 
        -53.80853, -53.84977, -53.89156, -53.93373, -53.9762, -54.01839, 
        -54.05993, -54.10049, -54.13979, -54.17765, -54.21435, -54.2505, 
        -54.28694, -54.32397, -54.36203, -54.40136, -54.44183, -54.48198, 
        -54.52344, -54.56525, -54.60707, -54.64926, -54.6916, -54.7341, 
        -54.77625, -54.81804, -54.85928, -54.89996, -54.94009, -54.97969, 
        -55.01865, -55.05672, -55.09356, -55.12883, -55.1622, -55.19346, 
        -55.22302, -55.25103, -55.27768, -55.30322, -55.32782, -55.3517, 
        -55.37398, -55.39661, -55.41888, -55.44042, -55.46104, -55.48077, 
        -55.49906, -55.51601, -55.53156, -55.54617, -55.56023, -55.57376, 
        -55.58626, -55.5968, -55.60455, -55.60874, -55.60878, -55.60484, 
        -55.59719, -55.58688, -55.57503, -55.56256, -55.54988, -55.53726, 
        -55.52458, -55.51152, -55.49741, -55.48048, -55.46211, -55.44118, 
        -55.41798, -55.39285, -55.36588, -55.3368, -55.30604, -55.27343, 
        -55.23882, -55.2023, -55.16396, -55.12418, -55.08376, -55.04277, 
        -55.00128, -54.95882, -54.91505, -54.86965, -54.82246, -54.77317, 
        -54.72185, -54.66899, -54.61491, -54.55993, -54.50415, -54.44773, 
        -54.39116, -54.33495, -54.28001, -54.22617, -54.17424, -54.12286, 
        -54.07401, -54.02599, -53.97852, -53.9309, -53.88266, -53.83354, 
        -53.78342, -53.73202, -53.67941, -53.62564, -53.57124, -53.51652, 
        -53.4618, -53.40733, -53.35336, -53.29993, -53.2468, -53.19361, 
        -53.14004, -53.08601, -53.03154, -52.97675, -52.92189, -52.86718, 
        -52.81316, -52.76055, -52.7097, -52.66047, -52.61217, -52.56469, 
        -52.51798, -52.47146, -52.42468, -52.37735, -52.32906, -52.27973, 
        -52.22996, -52.18042, -52.13139, -52.08255, -52.03649, -51.99261, 
        -51.95183, -51.91397, -51.87973, -51.84868, -51.82061, -51.79539, 
        -51.772, -51.7498, -51.72821, -51.70679, -51.68564, -51.6651, 
        -51.64601, -51.62928, -51.61579, -51.60619, -51.6007, -51.5989, 
        -51.60007,
  -48.12134, -48.26313, -48.38976, -48.50015, -48.59334, -48.66701, 
        -48.723, -48.75988, -48.77957, -48.78379, -48.7774, -48.76591, 
        -48.75628, -48.75655, -48.77425, -48.81508, -48.88234, -48.9758, 
        -49.09222, -49.22482, -49.36475, -49.50562, -49.63987, -49.76255, 
        -49.87112, -49.96527, -50.04634, -50.11673, -50.17942, -50.23724, 
        -50.29282, -50.34767, -50.40274, -50.45738, -50.51092, -50.56115, 
        -50.60935, -50.65387, -50.69504, -50.73301, -50.7687, -50.80268, 
        -50.83605, -50.86931, -50.9023, -50.93487, -50.96653, -50.99687, 
        -51.02606, -51.05396, -51.08107, -51.10644, -51.13265, -51.1586, 
        -51.18426, -51.20988, -51.23533, -51.26078, -51.28632, -51.31193, 
        -51.33778, -51.36383, -51.3899, -51.41629, -51.44294, -51.46998, 
        -51.49759, -51.52568, -51.5532, -51.58198, -51.61092, -51.63993, 
        -51.66863, -51.69661, -51.72346, -51.74894, -51.7732, -51.79627, 
        -51.81855, -51.8403, -51.86171, -51.88306, -51.90401, -51.92428, 
        -51.94363, -51.96209, -51.97918, -51.99738, -52.01633, -52.03672, 
        -52.05878, -52.08339, -52.11055, -52.14042, -52.17307, -52.20826, 
        -52.24623, -52.28629, -52.3283, -52.37221, -52.41806, -52.46603, 
        -52.51545, -52.56578, -52.61641, -52.6658, -52.71549, -52.76407, 
        -52.81144, -52.85795, -52.90449, -52.95224, -53.00133, -53.05172, 
        -53.10278, -53.1538, -53.20403, -53.25258, -53.29837, -53.34111, 
        -53.38036, -53.41663, -53.45038, -53.48235, -53.51321, -53.54283, 
        -53.57414, -53.60648, -53.64023, -53.67548, -53.71212, -53.75039, 
        -53.7893, -53.82858, -53.86781, -53.90687, -53.94621, -53.98597, 
        -54.02642, -54.06759, -54.1094, -54.15184, -54.1946, -54.23734, 
        -54.27952, -54.3207, -54.3606, -54.39816, -54.43607, -54.47367, 
        -54.51163, -54.55038, -54.59019, -54.63108, -54.67309, -54.71593, 
        -54.75893, -54.80183, -54.84468, -54.8878, -54.93113, -54.97445, 
        -55.0177, -55.06004, -55.10172, -55.14274, -55.18284, -55.22245, 
        -55.26145, -55.29961, -55.33566, -55.37145, -55.40586, -55.43879, 
        -55.47031, -55.50056, -55.52988, -55.55821, -55.58566, -55.61214, 
        -55.63763, -55.66242, -55.6865, -55.7099, -55.73233, -55.75391, 
        -55.77391, -55.7923, -55.80888, -55.82427, -55.83853, -55.85198, 
        -55.86396, -55.87402, -55.88107, -55.88437, -55.8836, -55.87777, 
        -55.86953, -55.85879, -55.84665, -55.83403, -55.82149, -55.80927, 
        -55.79708, -55.7844, -55.77073, -55.75501, -55.7367, -55.71538, 
        -55.69137, -55.66553, -55.63789, -55.60852, -55.57732, -55.54425, 
        -55.50941, -55.47245, -55.43348, -55.39283, -55.35115, -55.30909, 
        -55.26687, -55.22388, -55.17949, -55.13321, -55.08505, -55.0333, 
        -54.98071, -54.92669, -54.87129, -54.8152, -54.75818, -54.70065, 
        -54.64274, -54.58509, -54.52862, -54.4732, -54.41945, -54.36689, 
        -54.31556, -54.26535, -54.21536, -54.16532, -54.11464, -54.06294, 
        -54.0103, -53.95637, -53.90142, -53.84562, -53.78945, -53.73327, 
        -53.67734, -53.62185, -53.56688, -53.51226, -53.45802, -53.40374, 
        -53.34912, -53.29398, -53.23825, -53.18235, -53.12626, -53.0695, 
        -53.01465, -52.9613, -52.90985, -52.86008, -52.81152, -52.76339, 
        -52.71557, -52.6678, -52.61955, -52.57048, -52.52056, -52.46965, 
        -52.41841, -52.36785, -52.31804, -52.26949, -52.2226, -52.17782, 
        -52.13573, -52.09683, -52.0612, -52.02886, -51.99955, -51.97296, 
        -51.94818, -51.92442, -51.9011, -51.87801, -51.85534, -51.8335, 
        -51.81332, -51.79563, -51.78111, -51.77032, -51.76349, -51.76036, 
        -51.75994,
  -48.15198, -48.27782, -48.38876, -48.48373, -48.56223, -48.62302, 
        -48.66539, -48.68956, -48.69706, -48.69033, -48.67524, -48.6578, 
        -48.6455, -48.6469, -48.66895, -48.71919, -48.79934, -48.90854, 
        -49.04218, -49.19249, -49.35033, -49.50675, -49.6545, -49.78863, 
        -49.90654, -50.00832, -50.09524, -50.17037, -50.2373, -50.29902, 
        -50.35741, -50.41628, -50.47536, -50.53423, -50.59177, -50.647, 
        -50.69893, -50.74686, -50.79111, -50.83185, -50.86981, -50.90581, 
        -50.94094, -50.97596, -51.01088, -51.04449, -51.07834, -51.1111, 
        -51.1425, -51.17258, -51.20152, -51.22948, -51.25695, -51.28382, 
        -51.31036, -51.33651, -51.3623, -51.38804, -51.4138, -51.43981, 
        -51.46609, -51.49275, -51.51843, -51.54523, -51.57212, -51.59929, 
        -51.62679, -51.65471, -51.68294, -51.7115, -51.7403, -51.76928, 
        -51.79825, -51.82688, -51.85481, -51.88208, -51.90861, -51.93468, 
        -51.96045, -51.98613, -52.01075, -52.03598, -52.06047, -52.08368, 
        -52.10545, -52.12594, -52.14547, -52.16478, -52.18445, -52.20518, 
        -52.22756, -52.25179, -52.27843, -52.30745, -52.33908, -52.37332, 
        -52.40986, -52.44872, -52.48887, -52.53288, -52.57964, -52.62936, 
        -52.68138, -52.73476, -52.78878, -52.8428, -52.89581, -52.94823, 
        -52.99918, -53.04927, -53.09941, -53.15026, -53.20193, -53.25406, 
        -53.30655, -53.35886, -53.41014, -53.4597, -53.50534, -53.54903, 
        -53.58971, -53.62748, -53.66285, -53.69637, -53.72887, -53.76131, 
        -53.79412, -53.82792, -53.86285, -53.89904, -53.93673, -53.97557, 
        -54.01487, -54.05437, -54.09373, -54.13296, -54.17228, -54.21204, 
        -54.25248, -54.29281, -54.33482, -54.37735, -54.42022, -54.46296, 
        -54.50519, -54.54642, -54.58637, -54.6253, -54.66385, -54.70255, 
        -54.74189, -54.78226, -54.8238, -54.8666, -54.91036, -54.95462, 
        -54.99908, -55.04337, -55.08773, -55.13215, -55.17658, -55.2202, 
        -55.26431, -55.3075, -55.34961, -55.39071, -55.43094, -55.47056, 
        -55.5095, -55.54787, -55.5853, -55.62166, -55.65707, -55.69143, 
        -55.72485, -55.7575, -55.78935, -55.82047, -55.85064, -55.87972, 
        -55.90756, -55.93417, -55.95986, -55.98478, -56.009, -56.03246, 
        -56.05407, -56.07254, -56.09021, -56.10622, -56.12107, -56.13441, 
        -56.14636, -56.15599, -56.16255, -56.16526, -56.16379, -56.15852, 
        -56.1501, -56.13947, -56.12764, -56.11536, -56.10322, -56.09157, 
        -56.07994, -56.06771, -56.05415, -56.03826, -56.01944, -55.99754, 
        -55.97292, -55.94629, -55.91794, -55.88809, -55.85678, -55.8229, 
        -55.78794, -55.75094, -55.71165, -55.67061, -55.62855, -55.58585, 
        -55.54278, -55.49888, -55.45378, -55.40689, -55.3575, -55.30585, 
        -55.25188, -55.1967, -55.14037, -55.08279, -55.02433, -54.96517, 
        -54.90574, -54.84658, -54.7882, -54.73095, -54.67491, -54.61998, 
        -54.56609, -54.51282, -54.45992, -54.4069, -54.35346, -54.29927, 
        -54.24396, -54.1876, -54.13029, -54.07146, -54.01359, -53.95593, 
        -53.8987, -53.84203, -53.78597, -53.73046, -53.67517, -53.61988, 
        -53.56424, -53.50809, -53.45149, -53.39439, -53.3371, -53.28021, 
        -53.22453, -53.17059, -53.11859, -53.06829, -53.01902, -52.97013, 
        -52.92117, -52.87175, -52.82168, -52.77076, -52.71912, -52.66678, 
        -52.61459, -52.56315, -52.51277, -52.46373, -52.41628, -52.37072, 
        -52.32759, -52.28739, -52.25051, -52.21684, -52.18614, -52.15792, 
        -52.13128, -52.10567, -52.08057, -52.0559, -52.03096, -52.00824, 
        -51.98734, -51.96889, -51.95348, -51.94165, -51.93345, -51.92882, 
        -51.92664,
  -48.18597, -48.29266, -48.38448, -48.46061, -48.52094, -48.5649, 
        -48.5919, -48.60256, -48.5979, -48.58121, -48.56004, -48.54034, 
        -48.53026, -48.53782, -48.57102, -48.63452, -48.73023, -48.85608, 
        -49.00639, -49.17265, -49.34525, -49.51467, -49.67397, -49.81783, 
        -49.94297, -50.05146, -50.14426, -50.22443, -50.29589, -50.36216, 
        -50.42599, -50.48919, -50.55236, -50.61515, -50.67683, -50.73588, 
        -50.79149, -50.84296, -50.89037, -50.93419, -50.97378, -51.01244, 
        -51.05008, -51.08708, -51.12402, -51.1608, -51.19669, -51.23148, 
        -51.26493, -51.29687, -51.32742, -51.35696, -51.38564, -51.41375, 
        -51.44132, -51.46843, -51.49414, -51.52069, -51.54713, -51.57388, 
        -51.60097, -51.62819, -51.65548, -51.68256, -51.70968, -51.73685, 
        -51.76438, -51.79207, -51.81997, -51.84812, -51.87646, -51.90505, 
        -51.93376, -51.96143, -51.99001, -52.01849, -52.04698, -52.07584, 
        -52.10511, -52.13488, -52.16471, -52.19411, -52.22255, -52.24938, 
        -52.27443, -52.29766, -52.31947, -52.34071, -52.36184, -52.38355, 
        -52.40643, -52.42956, -52.45563, -52.48368, -52.5141, -52.54674, 
        -52.58146, -52.61855, -52.65839, -52.70176, -52.7489, -52.79963, 
        -52.85344, -52.90932, -52.96646, -53.02398, -53.08063, -53.13662, 
        -53.19137, -53.24561, -53.2987, -53.35256, -53.40677, -53.46105, 
        -53.51529, -53.56889, -53.62114, -53.67135, -53.71909, -53.76386, 
        -53.80564, -53.84478, -53.88171, -53.91694, -53.95131, -53.98552, 
        -54.02016, -54.0556, -54.092, -54.12955, -54.1681, -54.20636, 
        -54.24597, -54.28571, -54.32526, -54.36471, -54.40419, -54.44448, 
        -54.48505, -54.52661, -54.569, -54.6116, -54.65423, -54.69697, 
        -54.73909, -54.77985, -54.81959, -54.85854, -54.89765, -54.93703, 
        -54.97759, -55.01929, -55.06248, -55.10591, -55.15131, -55.19731, 
        -55.24352, -55.28955, -55.33549, -55.38128, -55.42702, -55.4726, 
        -55.51742, -55.56118, -55.60368, -55.645, -55.68542, -55.72525, 
        -55.76457, -55.80328, -55.84125, -55.87837, -55.91481, -55.95064, 
        -55.98594, -56.02074, -56.05501, -56.08775, -56.12067, -56.15233, 
        -56.18247, -56.21098, -56.23846, -56.26495, -56.29069, -56.31539, 
        -56.33838, -56.35913, -56.37822, -56.39519, -56.41036, -56.42414, 
        -56.43599, -56.44521, -56.45131, -56.45348, -56.45163, -56.44624, 
        -56.43801, -56.42792, -56.4168, -56.4054, -56.39408, -56.38308, 
        -56.37103, -56.359, -56.34513, -56.32869, -56.30916, -56.28655, 
        -56.26122, -56.23377, -56.20483, -56.17467, -56.14341, -56.11067, 
        -56.07598, -56.03913, -56.00009, -55.9591, -55.91682, -55.8736, 
        -55.82958, -55.78461, -55.73862, -55.69064, -55.64017, -55.58751, 
        -55.53269, -55.47629, -55.41873, -55.35976, -55.29976, -55.23902, 
        -55.17801, -55.11705, -55.05562, -54.99615, -54.93764, -54.88009, 
        -54.82344, -54.76722, -54.71131, -54.65532, -54.59914, -54.54236, 
        -54.48449, -54.42568, -54.3661, -54.30624, -54.24646, -54.18705, 
        -54.12831, -54.07027, -54.01331, -53.95692, -53.9007, -53.84459, 
        -53.78814, -53.73106, -53.67315, -53.61473, -53.55634, -53.49849, 
        -53.44189, -53.38708, -53.33421, -53.28296, -53.23266, -53.18262, 
        -53.13229, -53.08118, -53.02935, -52.97686, -52.92376, -52.86937, 
        -52.81639, -52.76427, -52.71337, -52.66381, -52.61577, -52.56947, 
        -52.52545, -52.48424, -52.44611, -52.41108, -52.37859, -52.34841, 
        -52.31956, -52.29187, -52.2649, -52.23875, -52.21379, -52.19038, 
        -52.16906, -52.15022, -52.1343, -52.12169, -52.11248, -52.10636, 
        -52.1026,
  -48.21521, -48.30035, -48.37068, -48.42575, -48.4649, -48.49015, 
        -48.50068, -48.49706, -48.48189, -48.45924, -48.43542, -48.41789, 
        -48.41478, -48.43415, -48.4821, -48.56273, -48.67679, -48.82096, 
        -48.98634, -49.16695, -49.35177, -49.53168, -49.69914, -49.85011, 
        -49.98271, -50.09712, -50.19527, -50.28071, -50.35734, -50.4287, 
        -50.49764, -50.56561, -50.63325, -50.70036, -50.76493, -50.82774, 
        -50.88671, -50.94162, -50.99245, -51.0396, -51.08356, -51.12513, 
        -51.16544, -51.20484, -51.24395, -51.28266, -51.32057, -51.35712, 
        -51.39224, -51.42598, -51.45712, -51.48815, -51.51831, -51.54785, 
        -51.5768, -51.60522, -51.63328, -51.66101, -51.68859, -51.71634, 
        -51.74429, -51.77237, -51.80019, -51.82777, -51.85505, -51.88237, 
        -51.90979, -51.9363, -51.96381, -51.99162, -52.01949, -52.04753, 
        -52.07567, -52.10394, -52.13264, -52.1619, -52.19215, -52.22355, 
        -52.25611, -52.28984, -52.32396, -52.35782, -52.39051, -52.42125, 
        -52.44907, -52.47575, -52.5007, -52.52443, -52.54749, -52.57077, 
        -52.59422, -52.61851, -52.64394, -52.67076, -52.69967, -52.7304, 
        -52.76317, -52.79824, -52.83625, -52.87853, -52.92533, -52.9766, 
        -53.0316, -53.08831, -53.14805, -53.20854, -53.26876, -53.32832, 
        -53.38707, -53.44539, -53.50332, -53.56091, -53.61803, -53.67455, 
        -53.73061, -53.7856, -53.83899, -53.89028, -53.93885, -53.9847, 
        -54.02773, -54.06834, -54.1068, -54.14273, -54.179, -54.21511, 
        -54.25175, -54.28898, -54.32688, -54.36566, -54.40504, -54.44484, 
        -54.48466, -54.52436, -54.56409, -54.60381, -54.64395, -54.68465, 
        -54.72597, -54.76789, -54.81044, -54.85335, -54.89586, -54.9381, 
        -54.97963, -55.01908, -55.05861, -55.09765, -55.13694, -55.17718, 
        -55.21824, -55.26101, -55.30544, -55.35142, -55.3984, -55.44609, 
        -55.49405, -55.54197, -55.58973, -55.63717, -55.68431, -55.73093, 
        -55.77657, -55.82085, -55.86369, -55.90524, -55.94588, -55.98611, 
        -56.02488, -56.06415, -56.10271, -56.14071, -56.17821, -56.21538, 
        -56.25239, -56.2892, -56.32585, -56.36211, -56.39756, -56.43174, 
        -56.46412, -56.49456, -56.52348, -56.55112, -56.57803, -56.60392, 
        -56.62814, -56.65039, -56.67055, -56.68884, -56.70494, -56.71908, 
        -56.73106, -56.74013, -56.74496, -56.74699, -56.74532, -56.74017, 
        -56.73257, -56.72349, -56.71347, -56.70321, -56.69307, -56.68271, 
        -56.67204, -56.65993, -56.64554, -56.62827, -56.60779, -56.5844, 
        -56.5583, -56.53022, -56.50069, -56.47011, -56.43881, -56.40624, 
        -56.37194, -56.33546, -56.29663, -56.25591, -56.21354, -56.16988, 
        -56.12506, -56.07895, -56.03064, -55.98161, -55.93001, -55.87616, 
        -55.82007, -55.76245, -55.70343, -55.64323, -55.58181, -55.51942, 
        -55.4566, -55.39378, -55.33152, -55.26979, -55.20867, -55.14859, 
        -55.08916, -55.03025, -54.97149, -54.91271, -54.85382, -54.79451, 
        -54.73431, -54.67317, -54.61133, -54.54939, -54.48761, -54.42631, 
        -54.36584, -54.30612, -54.248, -54.19079, -54.13395, -54.07701, 
        -54.01959, -53.96047, -53.90138, -53.84171, -53.78194, -53.72282, 
        -53.6652, -53.60944, -53.55554, -53.50306, -53.45127, -53.39964, 
        -53.34748, -53.29463, -53.24102, -53.18689, -53.13256, -53.07827, 
        -53.02456, -52.97189, -52.9203, -52.87011, -52.82146, -52.77457, 
        -52.72989, -52.68785, -52.64874, -52.61227, -52.57825, -52.54576, 
        -52.51461, -52.48471, -52.45592, -52.42842, -52.40251, -52.37862, 
        -52.35706, -52.33806, -52.32187, -52.30867, -52.29851, -52.29108, 
        -52.28561,
  -48.23288, -48.29507, -48.34272, -48.37577, -48.3945, -48.39993, 
        -48.39344, -48.37629, -48.35189, -48.32497, -48.3024, -48.29179, 
        -48.30045, -48.33521, -48.40285, -48.50421, -48.6384, -48.8007, 
        -48.98314, -49.17648, -49.37108, -49.55838, -49.73207, -49.88819, 
        -50.02538, -50.14449, -50.24776, -50.33871, -50.41992, -50.49681, 
        -50.57124, -50.64439, -50.71691, -50.78825, -50.85779, -50.92416, 
        -50.98663, -51.0449, -51.09925, -51.14986, -51.19737, -51.24243, 
        -51.28582, -51.32804, -51.36846, -51.40921, -51.44888, -51.48711, 
        -51.52389, -51.55917, -51.59298, -51.6255, -51.65722, -51.68826, 
        -51.71881, -51.74894, -51.77873, -51.80808, -51.83728, -51.86627, 
        -51.89537, -51.92334, -51.95198, -51.98002, -52.00778, -52.03519, 
        -52.06259, -52.09017, -52.11756, -52.14507, -52.17252, -52.19989, 
        -52.22737, -52.25512, -52.28363, -52.31335, -52.34488, -52.37861, 
        -52.4134, -52.45088, -52.48915, -52.52723, -52.56424, -52.59933, 
        -52.63218, -52.66268, -52.69099, -52.71786, -52.74346, -52.76834, 
        -52.79268, -52.81699, -52.8418, -52.86749, -52.89457, -52.92327, 
        -52.9528, -52.9859, -53.02238, -53.0632, -53.10927, -53.16011, 
        -53.21552, -53.27449, -53.33608, -53.39901, -53.46222, -53.52535, 
        -53.58809, -53.65047, -53.71237, -53.77358, -53.83402, -53.89341, 
        -53.9517, -54.00852, -54.06242, -54.11505, -54.16489, -54.21193, 
        -54.25621, -54.29821, -54.3382, -54.37682, -54.41493, -54.45312, 
        -54.49178, -54.53102, -54.57069, -54.61058, -54.6506, -54.69055, 
        -54.73029, -54.76987, -54.80956, -54.84954, -54.89009, -54.93044, 
        -54.97246, -55.01494, -55.05798, -55.10077, -55.14346, -55.18543, 
        -55.22656, -55.2666, -55.30598, -55.34505, -55.3847, -55.42504, 
        -55.46676, -55.51027, -55.55559, -55.60265, -55.65098, -55.7002, 
        -55.74989, -55.79963, -55.84923, -55.8975, -55.94619, -55.99394, 
        -56.04044, -56.08518, -56.12842, -56.17039, -56.21156, -56.25239, 
        -56.2929, -56.33276, -56.37208, -56.41089, -56.44951, -56.48797, 
        -56.52649, -56.56507, -56.60373, -56.64235, -56.68029, -56.71686, 
        -56.7513, -56.78352, -56.814, -56.84315, -56.87013, -56.89697, 
        -56.92222, -56.94567, -56.96711, -56.98643, -57.0035, -57.01818, 
        -57.0303, -57.03948, -57.04531, -57.04754, -57.04626, -57.0421, 
        -57.03572, -57.02797, -57.01937, -57.01029, -57.0012, -56.99192, 
        -56.98154, -56.96906, -56.9539, -56.93576, -56.91447, -56.89028, 
        -56.86343, -56.83462, -56.80359, -56.77273, -56.74114, -56.70847, 
        -56.67417, -56.63796, -56.59953, -56.55903, -56.51669, -56.47263, 
        -56.42708, -56.3796, -56.33087, -56.28006, -56.22715, -56.17177, 
        -56.11432, -56.0552, -55.99486, -55.9331, -55.87032, -55.8065, 
        -55.74241, -55.67766, -55.61338, -55.54976, -55.48669, -55.42426, 
        -55.36229, -55.30066, -55.23936, -55.17821, -55.11693, -55.05431, 
        -54.99187, -54.92869, -54.86485, -54.8008, -54.73684, -54.67333, 
        -54.61082, -54.5496, -54.49, -54.43151, -54.37378, -54.3161, 
        -54.25774, -54.19832, -54.13774, -54.0764, -54.0152, -53.95485, 
        -53.89608, -53.83916, -53.78384, -53.72969, -53.67606, -53.62246, 
        -53.5683, -53.51359, -53.45839, -53.40281, -53.34742, -53.29222, 
        -53.23765, -53.1839, -53.13165, -53.08064, -53.03122, -52.98376, 
        -52.93864, -52.89606, -52.85612, -52.81842, -52.78243, -52.74701, 
        -52.71374, -52.6818, -52.65126, -52.62243, -52.59565, -52.57129, 
        -52.54953, -52.53047, -52.51415, -52.50059, -52.48966, -52.48098, 
        -52.47393,
  -48.23722, -48.27668, -48.30119, -48.31138, -48.30854, -48.29399, 
        -48.27029, -48.2407, -48.20805, -48.18014, -48.16286, -48.1636, 
        -48.18911, -48.24556, -48.33583, -48.45999, -48.61525, -48.79564, 
        -48.99288, -49.19714, -49.39942, -49.59229, -49.7702, -49.929, 
        -50.0699, -50.19315, -50.30117, -50.39751, -50.48552, -50.56836, 
        -50.64861, -50.72712, -50.80433, -50.88013, -50.95345, -51.02361, 
        -51.08959, -51.15154, -51.20857, -51.26301, -51.31411, -51.36282, 
        -51.40966, -51.45499, -51.49909, -51.54192, -51.58337, -51.62323, 
        -51.6615, -51.69825, -51.73341, -51.76759, -51.80093, -51.83387, 
        -51.86552, -51.89767, -51.92943, -51.96061, -51.99137, -52.02195, 
        -52.05242, -52.08253, -52.11209, -52.1412, -52.16964, -52.19775, 
        -52.22554, -52.25331, -52.28084, -52.30816, -52.33525, -52.36112, 
        -52.38807, -52.41539, -52.44371, -52.47387, -52.50666, -52.54247, 
        -52.58096, -52.62165, -52.66363, -52.70577, -52.74694, -52.78615, 
        -52.82294, -52.85728, -52.88927, -52.91934, -52.94758, -52.97324, 
        -52.9988, -53.02348, -53.04779, -53.07218, -53.09739, -53.12402, 
        -53.15245, -53.18357, -53.21825, -53.25754, -53.3024, -53.35248, 
        -53.40762, -53.46709, -53.52981, -53.59476, -53.66073, -53.72717, 
        -53.79248, -53.85856, -53.9245, -53.98967, -54.05383, -54.11656, 
        -54.17754, -54.2368, -54.29371, -54.34801, -54.39936, -54.44757, 
        -54.49321, -54.53655, -54.57824, -54.6187, -54.65877, -54.69919, 
        -54.74012, -54.78137, -54.82265, -54.86245, -54.90287, -54.94273, 
        -54.9822, -55.02144, -55.06088, -55.10092, -55.14177, -55.18357, 
        -55.2261, -55.26907, -55.31232, -55.35541, -55.39798, -55.43974, 
        -55.48057, -55.52055, -55.55978, -55.59878, -55.63822, -55.67873, 
        -55.72086, -55.76397, -55.81014, -55.85838, -55.90795, -55.95863, 
        -56.00997, -56.06145, -56.11293, -56.16404, -56.21431, -56.26356, 
        -56.31114, -56.35689, -56.4009, -56.44363, -56.48545, -56.5271, 
        -56.56834, -56.60891, -56.64899, -56.68866, -56.72822, -56.76779, 
        -56.80755, -56.84668, -56.88712, -56.92776, -56.96792, -57.00665, 
        -57.04323, -57.07743, -57.10968, -57.14018, -57.16941, -57.1973, 
        -57.22349, -57.24788, -57.27037, -57.29042, -57.30804, -57.32306, 
        -57.33536, -57.34457, -57.35056, -57.35326, -57.35283, -57.34985, 
        -57.34489, -57.33875, -57.33171, -57.32433, -57.31564, -57.30714, 
        -57.29683, -57.28419, -57.2685, -57.24967, -57.2275, -57.20242, 
        -57.17502, -57.1459, -57.11523, -57.08392, -57.05198, -57.01914, 
        -56.98478, -56.94859, -56.9102, -56.86949, -56.82676, -56.78198, 
        -56.73532, -56.68655, -56.63578, -56.58294, -56.52808, -56.47119, 
        -56.41225, -56.35172, -56.28994, -56.22707, -56.16319, -56.09719, 
        -56.03168, -55.96581, -55.90039, -55.8353, -55.77043, -55.70601, 
        -55.64194, -55.5781, -55.51451, -55.45101, -55.38746, -55.32369, 
        -55.25927, -55.19415, -55.12833, -55.06221, -54.99606, -54.93045, 
        -54.86588, -54.80272, -54.74122, -54.68128, -54.62223, -54.56332, 
        -54.5035, -54.44252, -54.38039, -54.3175, -54.25477, -54.19297, 
        -54.13279, -54.07435, -54.01733, -53.9613, -53.90557, -53.8497, 
        -53.79338, -53.7359, -53.67904, -53.62204, -53.5653, -53.50888, 
        -53.45329, -53.39875, -53.34547, -53.29364, -53.24354, -53.19565, 
        -53.1501, -53.10696, -53.06612, -53.02719, -52.98973, -52.9535, 
        -52.91837, -52.88461, -52.85256, -52.82253, -52.79485, -52.76989, 
        -52.74781, -52.72851, -52.71192, -52.69794, -52.68632, -52.67661, 
        -52.6683,
  -48.2263, -48.24348, -48.24414, -48.2318, -48.20724, -48.17315, 
        -48.13304, -48.09211, -48.05562, -48.02964, -48.02135, -48.03775, 
        -48.08398, -48.16433, -48.27987, -48.42832, -48.60518, -48.80203, 
        -49.01239, -49.22587, -49.4342, -49.63068, -49.81107, -49.97335, 
        -50.11725, -50.24456, -50.35777, -50.45983, -50.55405, -50.64309, 
        -50.72903, -50.8129, -50.89402, -50.97385, -51.0509, -51.12444, 
        -51.19413, -51.25991, -51.32181, -51.38028, -51.4357, -51.4883, 
        -51.5388, -51.58738, -51.63427, -51.6792, -51.72247, -51.76387, 
        -51.80258, -51.84085, -51.87782, -51.91369, -51.94881, -51.98363, 
        -52.01838, -52.05291, -52.08686, -52.12031, -52.15302, -52.18533, 
        -52.21714, -52.24859, -52.27964, -52.30999, -52.33982, -52.36795, 
        -52.39672, -52.42497, -52.45291, -52.48043, -52.50746, -52.53419, 
        -52.56084, -52.58802, -52.61657, -52.64734, -52.68125, -52.71865, 
        -52.75945, -52.80302, -52.8482, -52.89383, -52.93856, -52.9805, 
        -53.02113, -53.05912, -53.09461, -53.12765, -53.15849, -53.18733, 
        -53.21416, -53.23935, -53.26324, -53.28664, -53.31041, -53.33514, 
        -53.36177, -53.39109, -53.42418, -53.46207, -53.50523, -53.55306, 
        -53.6073, -53.66652, -53.72995, -53.7962, -53.86432, -53.93331, 
        -54.00281, -54.07265, -54.14233, -54.21152, -54.27952, -54.34593, 
        -54.41043, -54.47248, -54.53183, -54.58804, -54.64105, -54.69101, 
        -54.73813, -54.78205, -54.82531, -54.86772, -54.91011, -54.95281, 
        -54.99594, -55.03901, -55.08162, -55.12337, -55.16397, -55.2036, 
        -55.24254, -55.28137, -55.32066, -55.36066, -55.40165, -55.44362, 
        -55.48643, -55.52982, -55.5733, -55.6165, -55.65904, -55.6997, 
        -55.74043, -55.78025, -55.81941, -55.85838, -55.89782, -55.93842, 
        -55.98084, -56.02542, -56.0723, -56.12127, -56.17186, -56.22374, 
        -56.27638, -56.32952, -56.38278, -56.43571, -56.48784, -56.53858, 
        -56.58748, -56.63439, -56.67954, -56.72338, -56.76549, -56.80812, 
        -56.85024, -56.89175, -56.93261, -56.97313, -57.01354, -57.05407, 
        -57.09498, -57.13634, -57.17833, -57.22062, -57.26257, -57.30328, 
        -57.34185, -57.37801, -57.41189, -57.44391, -57.47434, -57.50315, 
        -57.53023, -57.55539, -57.57845, -57.59913, -57.61712, -57.63235, 
        -57.64372, -57.65319, -57.65977, -57.66331, -57.66407, -57.6624, 
        -57.65897, -57.65445, -57.64915, -57.64336, -57.63678, -57.6289, 
        -57.619, -57.60618, -57.59011, -57.57058, -57.54785, -57.52239, 
        -57.49458, -57.46506, -57.43422, -57.40258, -57.37027, -57.33692, 
        -57.30217, -57.2655, -57.22665, -57.18554, -57.14207, -57.09533, 
        -57.04712, -56.99646, -56.94353, -56.8884, -56.8314, -56.77249, 
        -56.71193, -56.6501, -56.58709, -56.52314, -56.45812, -56.39222, 
        -56.32581, -56.25915, -56.19276, -56.12661, -56.06072, -55.99503, 
        -55.9293, -55.86363, -55.79798, -55.73243, -55.66697, -55.60124, 
        -55.53502, -55.46801, -55.40032, -55.33224, -55.26401, -55.19617, 
        -55.12922, -55.0638, -55.00026, -54.93837, -54.87655, -54.8158, 
        -54.7543, -54.69163, -54.62771, -54.56315, -54.49877, -54.43548, 
        -54.3738, -54.31361, -54.25459, -54.19622, -54.13814, -54.08007, 
        -54.02178, -53.96333, -53.90474, -53.84622, -53.78809, -53.73053, 
        -53.67384, -53.61821, -53.56389, -53.51122, -53.46054, -53.41218, 
        -53.36625, -53.32262, -53.28096, -53.24082, -53.20184, -53.16386, 
        -53.12707, -53.09179, -53.0584, -53.02728, -52.99873, -52.97304, 
        -52.95032, -52.93053, -52.91351, -52.89904, -52.88678, -52.87628, 
        -52.867,
  -48.19993, -48.19596, -48.17577, -48.14163, -48.09614, -48.04331, 
        -47.98818, -47.93727, -47.89754, -47.87609, -47.8796, -47.91443, 
        -47.98347, -48.09016, -48.23215, -48.40537, -48.60313, -48.81746, 
        -49.03942, -49.26058, -49.47348, -49.6727, -49.85497, -50.01929, 
        -50.16613, -50.2975, -50.41605, -50.52342, -50.62431, -50.71991, 
        -50.81174, -50.90068, -50.98732, -51.07117, -51.15188, -51.22921, 
        -51.30246, -51.37185, -51.43771, -51.5005, -51.56016, -51.617, 
        -51.67143, -51.7225, -51.77229, -51.81952, -51.86448, -51.9073, 
        -51.94859, -51.98858, -52.02744, -52.0652, -52.10244, -52.13934, 
        -52.17619, -52.21309, -52.24956, -52.28521, -52.3201, -52.35338, 
        -52.38698, -52.42015, -52.45303, -52.48528, -52.51698, -52.54782, 
        -52.57796, -52.60746, -52.63614, -52.66421, -52.6916, -52.71859, 
        -52.74557, -52.77318, -52.80231, -52.83388, -52.86792, -52.90686, 
        -52.94956, -52.99531, -53.04291, -53.0912, -53.13891, -53.18504, 
        -53.22893, -53.27011, -53.30868, -53.34468, -53.37812, -53.40902, 
        -53.43723, -53.46313, -53.48717, -53.51009, -53.53281, -53.55516, 
        -53.58035, -53.60838, -53.64023, -53.67669, -53.71816, -53.76527, 
        -53.81817, -53.87661, -53.93985, -54.0066, -54.07598, -54.14709, 
        -54.21934, -54.29239, -54.36561, -54.43861, -54.51066, -54.58105, 
        -54.64819, -54.71339, -54.77542, -54.83398, -54.88902, -54.94075, 
        -54.98952, -55.03618, -55.08146, -55.12615, -55.17093, -55.21593, 
        -55.26111, -55.30591, -55.34969, -55.39202, -55.43264, -55.47197, 
        -55.51056, -55.54913, -55.58829, -55.62725, -55.66826, -55.7103, 
        -55.75323, -55.79675, -55.84033, -55.88356, -55.92606, -55.96761, 
        -56.00819, -56.04792, -56.087, -56.12592, -56.16535, -56.206, 
        -56.24866, -56.29366, -56.34105, -56.39059, -56.44192, -56.49469, 
        -56.54845, -56.60192, -56.65677, -56.71149, -56.76545, -56.8179, 
        -56.86835, -56.9167, -56.96326, -57.00854, -57.05309, -57.09708, 
        -57.14041, -57.18297, -57.22477, -57.2662, -57.30756, -57.34908, 
        -57.39096, -57.43335, -57.47644, -57.52, -57.56335, -57.60559, 
        -57.64586, -57.68382, -57.71846, -57.75196, -57.78352, -57.81314, 
        -57.84089, -57.86665, -57.89022, -57.91128, -57.9295, -57.94486, 
        -57.95744, -57.96734, -57.97461, -57.97915, -57.98115, -57.98094, 
        -57.97906, -57.9761, -57.97229, -57.96777, -57.9622, -57.95493, 
        -57.94524, -57.93235, -57.91607, -57.89634, -57.87344, -57.84784, 
        -57.81895, -57.78941, -57.75861, -57.7268, -57.69402, -57.65996, 
        -57.62441, -57.58699, -57.5474, -57.50545, -57.46088, -57.4137, 
        -57.36373, -57.3109, -57.25547, -57.19771, -57.13821, -57.07727, 
        -57.01512, -56.95198, -56.88781, -56.82286, -56.75706, -56.69046, 
        -56.62337, -56.55607, -56.48903, -56.42236, -56.35589, -56.28938, 
        -56.22255, -56.15546, -56.08723, -56.01995, -55.95264, -55.88506, 
        -55.81702, -55.74829, -55.67889, -55.60896, -55.53866, -55.46856, 
        -55.39927, -55.33144, -55.26549, -55.20121, -55.13807, -55.0751, 
        -55.01149, -54.9468, -54.88101, -54.81474, -54.74878, -54.68396, 
        -54.62059, -54.55844, -54.49723, -54.43652, -54.37607, -54.31573, 
        -54.25533, -54.19495, -54.13463, -54.07458, -54.01504, -53.95624, 
        -53.89843, -53.8418, -53.7866, -53.7332, -53.68197, -53.63319, 
        -53.58678, -53.54145, -53.49876, -53.45725, -53.41666, -53.37704, 
        -53.33869, -53.30204, -53.26747, -53.23532, -53.20591, -53.17942, 
        -53.15593, -53.13541, -53.11773, -53.10263, -53.08976, -53.07862, 
        -53.06867,
  -48.16255, -48.13873, -48.09771, -48.04301, -47.97805, -47.90815, 
        -47.8386, -47.77946, -47.73808, -47.72301, -47.74025, -47.7954, 
        -47.89059, -48.02447, -48.19301, -48.39003, -48.60719, -48.83659, 
        -49.06898, -49.29651, -49.51317, -49.71374, -49.89799, -50.0648, 
        -50.21523, -50.35117, -50.47553, -50.59053, -50.69836, -50.80046, 
        -50.8983, -50.99261, -51.08364, -51.17155, -51.25597, -51.33681, 
        -51.41356, -51.48583, -51.55596, -51.62244, -51.68636, -51.74759, 
        -51.80639, -51.86192, -51.91465, -51.96425, -52.01101, -52.05546, 
        -52.09836, -52.14032, -52.18087, -52.22104, -52.26056, -52.29874, 
        -52.33778, -52.37667, -52.41557, -52.4537, -52.49107, -52.52757, 
        -52.56337, -52.5988, -52.63386, -52.66851, -52.70266, -52.73591, 
        -52.76824, -52.7994, -52.82939, -52.85852, -52.88567, -52.91354, 
        -52.94152, -52.97015, -53.00046, -53.03317, -53.06958, -53.10991, 
        -53.15399, -53.20119, -53.25043, -53.30069, -53.35039, -53.39883, 
        -53.44526, -53.48914, -53.53048, -53.5691, -53.6039, -53.63668, 
        -53.66649, -53.69364, -53.71844, -53.74148, -53.76391, -53.78671, 
        -53.81124, -53.83851, -53.86934, -53.9045, -53.94436, -53.98978, 
        -54.04096, -54.09788, -54.15998, -54.22641, -54.29633, -54.36785, 
        -54.44209, -54.5177, -54.59422, -54.67094, -54.74683, -54.82095, 
        -54.8927, -54.96128, -55.02625, -55.08754, -55.14469, -55.19831, 
        -55.24897, -55.29775, -55.34536, -55.39247, -55.43975, -55.48713, 
        -55.53436, -55.57965, -55.62428, -55.66696, -55.70762, -55.74686, 
        -55.78529, -55.82379, -55.86308, -55.90315, -55.94431, -55.98638, 
        -56.02924, -56.07269, -56.11623, -56.15934, -56.2016, -56.24286, 
        -56.28324, -56.32299, -56.36183, -56.40069, -56.44047, -56.47977, 
        -56.52257, -56.56786, -56.6156, -56.66559, -56.71743, -56.77082, 
        -56.8254, -56.88095, -56.93717, -56.99347, -57.04916, -57.10322, 
        -57.15533, -57.20521, -57.25343, -57.30036, -57.3466, -57.39214, 
        -57.4368, -57.48059, -57.52355, -57.5663, -57.60884, -57.65042, 
        -57.69327, -57.73669, -57.78066, -57.82498, -57.86907, -57.91224, 
        -57.95382, -57.99338, -58.03062, -58.06545, -58.09801, -58.1283, 
        -58.15684, -58.18315, -58.2071, -58.22847, -58.24694, -58.26255, 
        -58.27538, -58.28564, -58.29358, -58.29916, -58.30239, -58.30357, 
        -58.30299, -58.30034, -58.29783, -58.2944, -58.2895, -58.28261, 
        -58.273, -58.26023, -58.24411, -58.22452, -58.20172, -58.17628, 
        -58.14869, -58.11953, -58.08904, -58.05713, -58.02389, -57.9891, 
        -57.95266, -57.91426, -57.87358, -57.8305, -57.78463, -57.73582, 
        -57.68383, -57.62847, -57.57041, -57.51008, -57.44783, -57.38474, 
        -57.32083, -57.25644, -57.1902, -57.12456, -57.05835, -56.99111, 
        -56.92352, -56.85582, -56.78836, -56.72128, -56.65434, -56.58725, 
        -56.51978, -56.45179, -56.38332, -56.31448, -56.24534, -56.17607, 
        -56.10627, -56.03575, -55.96469, -55.89299, -55.82083, -55.74866, 
        -55.67722, -55.6069, -55.5383, -55.47129, -55.40544, -55.33978, 
        -55.27361, -55.20667, -55.1391, -55.07125, -55.0037, -54.93733, 
        -54.87225, -54.80799, -54.74468, -54.68057, -54.61774, -54.5551, 
        -54.49259, -54.43027, -54.36822, -54.30657, -54.24558, -54.18567, 
        -54.12696, -54.06953, -54.01364, -53.9596, -53.90798, -53.85882, 
        -53.81167, -53.76615, -53.72202, -53.67885, -53.6365, -53.5952, 
        -53.55532, -53.5174, -53.48164, -53.44859, -53.41841, -53.39118, 
        -53.3669, -53.34551, -53.32698, -53.3112, -53.29763, -53.286, 
        -53.27565,
  -48.11464, -48.07104, -48.01121, -47.93768, -47.85533, -47.77057, 
        -47.69112, -47.62644, -47.58586, -47.57822, -47.6103, -47.68545, 
        -47.80432, -47.96374, -48.15707, -48.37626, -48.61104, -48.85426, 
        -49.09653, -49.33061, -49.55122, -49.75547, -49.94225, -50.11211, 
        -50.2667, -50.40812, -50.53875, -50.66054, -50.77533, -50.88419, 
        -50.9882, -51.08688, -51.18267, -51.27457, -51.36251, -51.44674, 
        -51.52736, -51.60462, -51.67866, -51.7495, -51.81764, -51.88303, 
        -51.94552, -52.0048, -52.06044, -52.11262, -52.16166, -52.20703, 
        -52.25183, -52.29568, -52.33867, -52.38111, -52.42284, -52.46408, 
        -52.50505, -52.54594, -52.58702, -52.62759, -52.66741, -52.7064, 
        -52.74478, -52.78294, -52.82074, -52.85823, -52.89424, -52.93023, 
        -52.96509, -52.99852, -53.03059, -53.06125, -53.09104, -53.12041, 
        -53.15003, -53.18045, -53.21243, -53.24684, -53.28473, -53.32635, 
        -53.3716, -53.41982, -53.47002, -53.52041, -53.57166, -53.62184, 
        -53.67012, -53.71598, -53.75951, -53.8003, -53.83823, -53.87299, 
        -53.90448, -53.93319, -53.95924, -53.98338, -54.00638, -54.02935, 
        -54.05395, -54.081, -54.11142, -54.14567, -54.18322, -54.22709, 
        -54.27647, -54.33163, -54.39212, -54.45718, -54.52653, -54.59915, 
        -54.67458, -54.75215, -54.83111, -54.91088, -54.99008, -55.06774, 
        -55.14283, -55.21455, -55.28274, -55.3467, -55.40649, -55.46144, 
        -55.51431, -55.56549, -55.61554, -55.66521, -55.71476, -55.76408, 
        -55.81304, -55.8606, -55.9062, -55.9494, -55.99034, -56.0299, 
        -56.06873, -56.10777, -56.14749, -56.18808, -56.22971, -56.27207, 
        -56.31509, -56.35848, -56.40182, -56.44368, -56.48562, -56.52658, 
        -56.56666, -56.60605, -56.64494, -56.68371, -56.72306, -56.76377, 
        -56.80663, -56.85185, -56.89957, -56.94956, -57.00158, -57.0553, 
        -57.11034, -57.16657, -57.22366, -57.28106, -57.33795, -57.39344, 
        -57.44697, -57.49847, -57.54726, -57.59586, -57.64371, -57.69082, 
        -57.73707, -57.78236, -57.82684, -57.87102, -57.91504, -57.95908, 
        -58.00318, -58.04746, -58.0922, -58.13704, -58.18163, -58.22529, 
        -58.26748, -58.3079, -58.34606, -58.38183, -58.41519, -58.44626, 
        -58.47533, -58.50216, -58.52661, -58.54736, -58.56618, -58.58218, 
        -58.59547, -58.6064, -58.61512, -58.62164, -58.6261, -58.62854, 
        -58.62925, -58.62863, -58.62689, -58.6241, -58.61965, -58.61303, 
        -58.60358, -58.59087, -58.57501, -58.55574, -58.53341, -58.50841, 
        -58.48129, -58.45271, -58.42257, -58.39085, -58.35736, -58.32195, 
        -58.28472, -58.24531, -58.20257, -58.15815, -58.11072, -58.06025, 
        -58.00624, -57.94878, -57.88823, -57.82528, -57.76109, -57.69599, 
        -57.63041, -57.56444, -57.49811, -57.43169, -57.36479, -57.29735, 
        -57.22941, -57.16123, -57.09338, -57.02578, -56.95828, -56.8905, 
        -56.82206, -56.75309, -56.68344, -56.61332, -56.54271, -56.47163, 
        -56.40019, -56.32813, -56.25547, -56.18217, -56.10829, -56.03439, 
        -55.95985, -55.88729, -55.81609, -55.74625, -55.67753, -55.60913, 
        -55.54048, -55.4713, -55.40168, -55.33218, -55.26322, -55.19531, 
        -55.12848, -55.06246, -54.99704, -54.93184, -54.86673, -54.80169, 
        -54.73679, -54.67225, -54.60817, -54.54483, -54.48246, -54.42134, 
        -54.36171, -54.30363, -54.2473, -54.19294, -54.14076, -54.09077, 
        -54.04257, -53.99577, -53.94999, -53.90504, -53.86104, -53.81822, 
        -53.777, -53.7378, -53.70105, -53.66714, -53.63622, -53.60831, 
        -53.58332, -53.56117, -53.54182, -53.52417, -53.50996, -53.49775, 
        -53.48693,
  -48.05844, -47.99828, -47.92125, -47.83097, -47.73374, -47.63678, 
        -47.54923, -47.48116, -47.44302, -47.44391, -47.48946, -47.58389, 
        -47.72508, -47.90751, -48.12272, -48.36149, -48.61318, -48.86863, 
        -49.11996, -49.36056, -49.58606, -49.79432, -49.98509, -50.15941, 
        -50.31958, -50.46635, -50.60412, -50.73325, -50.85513, -50.97057, 
        -51.08054, -51.18558, -51.28615, -51.3822, -51.47404, -51.5619, 
        -51.64618, -51.72726, -51.80516, -51.88018, -51.95238, -52.02056, 
        -52.08666, -52.1492, -52.20796, -52.26302, -52.31469, -52.36375, 
        -52.41106, -52.45739, -52.50285, -52.54743, -52.5914, -52.63449, 
        -52.67714, -52.71993, -52.76273, -52.80558, -52.84713, -52.88893, 
        -52.93023, -52.97144, -53.01238, -53.05299, -53.09312, -53.1322, 
        -53.17005, -53.20634, -53.24078, -53.27377, -53.30573, -53.33747, 
        -53.36926, -53.40194, -53.43621, -53.47175, -53.51143, -53.55435, 
        -53.60042, -53.64933, -53.70012, -53.75211, -53.80407, -53.8552, 
        -53.90466, -53.95206, -53.99732, -54.0399, -54.07959, -54.1163, 
        -54.15001, -54.18076, -54.20885, -54.2338, -54.25846, -54.28279, 
        -54.30838, -54.33596, -54.36638, -54.40028, -54.43804, -54.48056, 
        -54.52795, -54.5806, -54.63858, -54.70142, -54.76905, -54.84072, 
        -54.91615, -54.99491, -55.07594, -55.15819, -55.23912, -55.3196, 
        -55.39776, -55.47271, -55.54406, -55.61092, -55.67335, -55.7319, 
        -55.7874, -55.84121, -55.89377, -55.94566, -55.99726, -56.04834, 
        -56.0987, -56.14731, -56.1936, -56.23753, -56.27925, -56.31965, 
        -56.35935, -56.39827, -56.43902, -56.48053, -56.52301, -56.56577, 
        -56.60882, -56.65208, -56.69515, -56.73767, -56.77919, -56.8197, 
        -56.85937, -56.89846, -56.93716, -56.97588, -57.01525, -57.05606, 
        -57.09927, -57.14405, -57.19169, -57.24172, -57.2939, -57.34659, 
        -57.40178, -57.45823, -57.51552, -57.57333, -57.63083, -57.68715, 
        -57.74183, -57.79473, -57.84615, -57.8965, -57.94605, -57.99479, 
        -58.04275, -58.08972, -58.13601, -58.18205, -58.22784, -58.27343, 
        -58.31891, -58.36427, -58.40968, -58.45481, -58.49939, -58.54313, 
        -58.58455, -58.62541, -58.66413, -58.70042, -58.73424, -58.76605, 
        -58.79572, -58.82297, -58.84771, -58.86987, -58.88907, -58.90545, 
        -58.91921, -58.93065, -58.94018, -58.94762, -58.9532, -58.95701, 
        -58.95836, -58.95852, -58.95739, -58.95507, -58.95066, -58.94408, 
        -58.93476, -58.92231, -58.90683, -58.88702, -58.8651, -58.84071, 
        -58.81433, -58.78651, -58.75693, -58.72545, -58.69195, -58.65619, 
        -58.61824, -58.57783, -58.53494, -58.48916, -58.44033, -58.38827, 
        -58.33248, -58.27306, -58.21057, -58.14577, -58.07977, -58.0129, 
        -57.94563, -57.87836, -57.81118, -57.74402, -57.67671, -57.609, 
        -57.54088, -57.47228, -57.40398, -57.33564, -57.26714, -57.19737, 
        -57.12797, -57.05793, -56.98707, -56.9155, -56.84336, -56.77068, 
        -56.69762, -56.62399, -56.54984, -56.47528, -56.4, -56.32459, 
        -56.24934, -56.17464, -56.10099, -56.02839, -55.95679, -55.8856, 
        -55.81439, -55.74307, -55.67153, -55.6004, -55.52991, -55.46036, 
        -55.3918, -55.32399, -55.25668, -55.18937, -55.12204, -55.05461, 
        -54.98729, -54.92046, -54.85435, -54.78925, -54.72548, -54.66331, 
        -54.60292, -54.54435, -54.48765, -54.43195, -54.37916, -54.32843, 
        -54.27884, -54.2304, -54.1827, -54.13592, -54.09036, -54.04623, 
        -54.00376, -53.96333, -53.92542, -53.89046, -53.85881, -53.83024, 
        -53.80473, -53.78193, -53.76183, -53.74438, -53.72945, -53.71664, 
        -53.70515,
  -47.99515, -47.91883, -47.82654, -47.72243, -47.61351, -47.50687, 
        -47.41473, -47.34671, -47.31314, -47.32327, -47.38317, -47.49443, 
        -47.65425, -47.85572, -48.08932, -48.34434, -48.60994, -48.87667, 
        -49.1367, -49.38457, -49.61511, -49.82885, -50.02512, -50.20559, 
        -50.37239, -50.52769, -50.67311, -50.80997, -50.93925, -51.06163, 
        -51.17775, -51.28815, -51.39335, -51.49385, -51.5899, -51.68073, 
        -51.76879, -51.85347, -51.93534, -52.01437, -52.09044, -52.1633, 
        -52.2328, -52.29853, -52.36019, -52.41817, -52.47293, -52.52528, 
        -52.57562, -52.62494, -52.67298, -52.71901, -52.7648, -52.80974, 
        -52.8541, -52.89824, -52.9427, -52.98738, -53.03234, -53.07721, 
        -53.12169, -53.16615, -53.21041, -53.25449, -53.29785, -53.34018, 
        -53.38122, -53.42059, -53.45704, -53.49295, -53.52781, -53.56224, 
        -53.59686, -53.63213, -53.66899, -53.70786, -53.74936, -53.7937, 
        -53.84089, -53.89043, -53.9417, -53.99395, -54.04631, -54.09805, 
        -54.14841, -54.19696, -54.24245, -54.28667, -54.32832, -54.36711, 
        -54.40302, -54.43621, -54.4667, -54.49543, -54.52251, -54.54902, 
        -54.5763, -54.60517, -54.63655, -54.67067, -54.70799, -54.74917, 
        -54.79459, -54.84488, -54.89996, -54.95888, -55.02378, -55.09344, 
        -55.16783, -55.24665, -55.32852, -55.41218, -55.49617, -55.57927, 
        -55.66022, -55.7381, -55.81229, -55.88207, -55.94754, -56.00895, 
        -56.06724, -56.12349, -56.1783, -56.23236, -56.28569, -56.33711, 
        -56.38851, -56.43791, -56.48531, -56.5302, -56.57302, -56.61454, 
        -56.65551, -56.6969, -56.73904, -56.78183, -56.82508, -56.86826, 
        -56.91159, -56.95493, -56.9977, -57.03992, -57.08117, -57.12156, 
        -57.16107, -57.20016, -57.23902, -57.27707, -57.31678, -57.3578, 
        -57.40062, -57.44566, -57.49316, -57.54277, -57.59442, -57.64782, 
        -57.70275, -57.75888, -57.81555, -57.87294, -57.9303, -57.98688, 
        -58.04221, -58.09614, -58.1489, -58.20085, -58.25227, -58.3028, 
        -58.35265, -58.40168, -58.44908, -58.4971, -58.54473, -58.59203, 
        -58.63886, -58.68526, -58.73119, -58.77654, -58.82111, -58.86458, 
        -58.90676, -58.94745, -58.98604, -59.02249, -59.05665, -59.0887, 
        -59.11868, -59.14634, -59.17154, -59.19381, -59.21326, -59.23013, 
        -59.24459, -59.25702, -59.26733, -59.27622, -59.28273, -59.28632, 
        -59.28859, -59.28917, -59.28825, -59.28557, -59.2809, -59.27403, 
        -59.26455, -59.25218, -59.23682, -59.21838, -59.1972, -59.17358, 
        -59.14805, -59.12089, -59.09182, -59.06075, -59.0273, -58.99133, 
        -58.95282, -58.91163, -58.86785, -58.821, -58.77113, -58.71799, 
        -58.66122, -58.6009, -58.53738, -58.47171, -58.40443, -58.33524, 
        -58.26681, -58.19834, -58.1301, -58.06212, -57.99414, -57.92603, 
        -57.8575, -57.78868, -57.71941, -57.65007, -57.58049, -57.5105, 
        -57.43973, -57.36819, -57.29585, -57.22297, -57.1493, -57.07502, 
        -57.00054, -56.92537, -56.85022, -56.7744, -56.69802, -56.62128, 
        -56.54455, -56.46816, -56.39241, -56.3175, -56.2434, -56.16971, 
        -56.09623, -56.02267, -55.94915, -55.87603, -55.80364, -55.73125, 
        -55.66082, -55.59104, -55.52175, -55.45245, -55.38295, -55.31317, 
        -55.24357, -55.17452, -55.10637, -55.0396, -54.97448, -54.91124, 
        -54.85, -54.79076, -54.73351, -54.67822, -54.62473, -54.57278, 
        -54.52187, -54.47173, -54.42237, -54.37407, -54.32719, -54.28204, 
        -54.23845, -54.19672, -54.15768, -54.1217, -54.08916, -54.05976, 
        -54.03349, -54.01001, -53.98919, -53.97098, -53.9553, -53.94197, 
        -53.9299,
  -47.92444, -47.83326, -47.72739, -47.61215, -47.49533, -47.38498, 
        -47.29202, -47.22683, -47.19989, -47.2197, -47.29176, -47.41708, 
        -47.59191, -47.80798, -48.05443, -48.32214, -48.59908, -48.87561, 
        -49.14455, -49.40003, -49.63901, -49.86007, -50.06378, -50.25209, 
        -50.42712, -50.59072, -50.74447, -50.88939, -51.02624, -51.15559, 
        -51.27708, -51.39311, -51.50334, -51.60859, -51.70901, -51.80516, 
        -51.89749, -51.98617, -52.07188, -52.15451, -52.23417, -52.31056, 
        -52.38326, -52.45195, -52.51669, -52.57765, -52.63465, -52.6903, 
        -52.74431, -52.79681, -52.84795, -52.89742, -52.94534, -52.99194, 
        -53.03777, -53.08315, -53.12892, -53.17538, -53.22258, -53.27022, 
        -53.31813, -53.36618, -53.41299, -53.46045, -53.50719, -53.55288, 
        -53.59704, -53.63982, -53.68071, -53.72004, -53.75824, -53.79576, 
        -53.83338, -53.87162, -53.91119, -53.95259, -53.99617, -54.04205, 
        -54.09028, -54.1405, -54.19128, -54.24385, -54.29644, -54.34844, 
        -54.39933, -54.44885, -54.49657, -54.54219, -54.58563, -54.62661, 
        -54.66511, -54.70131, -54.73503, -54.76682, -54.79705, -54.82675, 
        -54.85662, -54.88746, -54.91924, -54.95411, -54.99156, -55.03183, 
        -55.07541, -55.12307, -55.17496, -55.23157, -55.2931, -55.35986, 
        -55.43228, -55.50999, -55.59192, -55.67633, -55.76168, -55.84669, 
        -55.92995, -56.01059, -56.08751, -56.16002, -56.22725, -56.29144, 
        -56.3525, -56.41117, -56.4681, -56.52387, -56.57858, -56.63229, 
        -56.68456, -56.73485, -56.78302, -56.8291, -56.87336, -56.91641, 
        -56.95888, -57.00183, -57.04546, -57.08963, -57.13382, -57.17765, 
        -57.22122, -57.26365, -57.30655, -57.34874, -57.38984, -57.42989, 
        -57.46963, -57.50885, -57.54823, -57.58797, -57.62848, -57.67011, 
        -57.71322, -57.7582, -57.80532, -57.85453, -57.90574, -57.95857, 
        -58.01277, -58.0681, -58.12375, -58.18005, -58.23651, -58.29154, 
        -58.3469, -58.40144, -58.4553, -58.50874, -58.56181, -58.61435, 
        -58.66627, -58.71752, -58.76825, -58.81837, -58.86786, -58.91665, 
        -58.96467, -59.01199, -59.05846, -59.10392, -59.14827, -59.1911, 
        -59.23262, -59.27259, -59.31071, -59.34683, -59.3809, -59.41304, 
        -59.44319, -59.46991, -59.49503, -59.51731, -59.53694, -59.55409, 
        -59.56945, -59.583, -59.59476, -59.60453, -59.6123, -59.61752, 
        -59.62036, -59.62094, -59.61966, -59.61631, -59.61086, -59.60324, 
        -59.59333, -59.58087, -59.56555, -59.54742, -59.5268, -59.50398, 
        -59.47932, -59.45283, -59.42423, -59.39348, -59.36023, -59.32346, 
        -59.28461, -59.24288, -59.19832, -59.15084, -59.1005, -59.04702, 
        -58.99006, -58.92985, -58.86638, -58.80054, -58.73285, -58.66398, 
        -58.59474, -58.52547, -58.45658, -58.388, -58.31934, -58.25067, 
        -58.18162, -58.11229, -58.04211, -57.9716, -57.90066, -57.82912, 
        -57.75684, -57.68368, -57.60962, -57.53489, -57.4596, -57.38395, 
        -57.308, -57.23172, -57.15515, -57.07743, -57.00019, -56.92243, 
        -56.84452, -56.7667, -56.68928, -56.61257, -56.53647, -56.4607, 
        -56.38504, -56.30935, -56.23377, -56.15854, -56.08393, -56.01029, 
        -55.93763, -55.86575, -55.79436, -55.72305, -55.65166, -55.57983, 
        -55.50817, -55.43716, -55.36702, -55.2986, -55.23202, -55.16766, 
        -55.10548, -55.04531, -54.98727, -54.93116, -54.87673, -54.82351, 
        -54.77116, -54.71953, -54.66865, -54.61913, -54.57117, -54.52503, 
        -54.48089, -54.43858, -54.3982, -54.36087, -54.326, -54.29573, 
        -54.26877, -54.24457, -54.22319, -54.20414, -54.18764, -54.17331, 
        -54.16077,
  -47.84868, -47.74388, -47.62659, -47.5038, -47.38202, -47.27095, 
        -47.18093, -47.1221, -47.10384, -47.13266, -47.2154, -47.35148, 
        -47.53662, -47.76315, -48.02023, -48.29688, -48.58298, -48.86827, 
        -49.14575, -49.40987, -49.6573, -49.88739, -50.10041, -50.29805, 
        -50.48145, -50.6543, -50.81685, -50.96998, -51.11457, -51.25092, 
        -51.37978, -51.50175, -51.61745, -51.72773, -51.83317, -51.93393, 
        -52.03087, -52.1241, -52.21386, -52.30026, -52.38237, -52.4618, 
        -52.53744, -52.60917, -52.67697, -52.74119, -52.80262, -52.86182, 
        -52.9194, -52.97533, -53.02943, -53.08163, -53.13169, -53.18022, 
        -53.22747, -53.27436, -53.32043, -53.36839, -53.41742, -53.46776, 
        -53.5191, -53.57083, -53.62222, -53.67321, -53.72336, -53.77236, 
        -53.82006, -53.86608, -53.91039, -53.95349, -53.99521, -54.03619, 
        -54.07705, -54.11746, -54.15974, -54.20357, -54.24928, -54.29684, 
        -54.34626, -54.39734, -54.44969, -54.50269, -54.5556, -54.60787, 
        -54.65928, -54.7096, -54.75851, -54.80569, -54.85107, -54.89443, 
        -54.93582, -54.97417, -55.01148, -55.04701, -55.08103, -55.11435, 
        -55.14743, -55.18099, -55.21566, -55.25172, -55.28951, -55.32925, 
        -55.37138, -55.41677, -55.46574, -55.5188, -55.57684, -55.64042, 
        -55.71017, -55.78584, -55.86561, -55.94982, -56.03592, -56.12235, 
        -56.20757, -56.29036, -56.36972, -56.44469, -56.51551, -56.5822, 
        -56.64563, -56.70645, -56.76522, -56.82256, -56.87857, -56.93336, 
        -56.98658, -57.03784, -57.08709, -57.13428, -57.17976, -57.22331, 
        -57.26734, -57.31187, -57.35698, -57.40224, -57.44727, -57.49161, 
        -57.53542, -57.57882, -57.622, -57.66447, -57.70543, -57.74592, 
        -57.78598, -57.82602, -57.8666, -57.90739, -57.94894, -57.99158, 
        -58.03542, -58.08057, -58.12743, -58.17528, -58.22601, -58.27825, 
        -58.33174, -58.38557, -58.43996, -58.49482, -58.54952, -58.60441, 
        -58.65918, -58.71385, -58.76844, -58.82309, -58.87773, -58.93215, 
        -58.98625, -59.03974, -59.09271, -59.14493, -59.19609, -59.24615, 
        -59.29505, -59.34304, -59.38995, -59.43439, -59.4782, -59.52032, 
        -59.56059, -59.59937, -59.63647, -59.67188, -59.70552, -59.73741, 
        -59.76738, -59.79491, -59.8197, -59.84175, -59.8614, -59.8791, 
        -59.89515, -59.90989, -59.92296, -59.93397, -59.94254, -59.94833, 
        -59.95141, -59.95176, -59.94965, -59.94516, -59.93855, -59.9299, 
        -59.91801, -59.90482, -59.88929, -59.8713, -59.85127, -59.82915, 
        -59.80518, -59.77919, -59.75096, -59.72043, -59.68736, -59.65162, 
        -59.61289, -59.57113, -59.5263, -59.47873, -59.42854, -59.37558, 
        -59.31955, -59.2604, -59.19802, -59.13291, -59.06579, -58.99691, 
        -58.92749, -58.85793, -58.78871, -58.71963, -58.65053, -58.5813, 
        -58.51156, -58.4414, -58.36955, -58.29794, -58.22562, -58.15242, 
        -58.07829, -58.00332, -57.92741, -57.85088, -57.77389, -57.69669, 
        -57.61932, -57.54172, -57.46426, -57.38649, -57.30842, -57.22994, 
        -57.15114, -57.07233, -56.99377, -56.91567, -56.83797, -56.76049, 
        -56.68284, -56.60508, -56.52729, -56.44992, -56.3727, -56.29658, 
        -56.22131, -56.14713, -56.07359, -56.00037, -55.92706, -55.85364, 
        -55.78012, -55.70724, -55.63549, -55.56539, -55.49734, -55.43071, 
        -55.3673, -55.30609, -55.24728, -55.19003, -55.13425, -55.07963, 
        -55.02573, -54.97301, -54.92107, -54.87046, -54.8218, -54.775, 
        -54.7301, -54.68661, -54.64534, -54.6069, -54.57188, -54.54051, 
        -54.51257, -54.48773, -54.46548, -54.44581, -54.42858, -54.4131, 
        -54.39928,
  -47.76804, -47.65059, -47.52424, -47.39677, -47.2731, -47.16492, 
        -47.08161, -47.03194, -47.02396, -47.0641, -47.15602, -47.29979, 
        -47.49143, -47.72368, -47.98635, -48.26908, -48.56178, -48.85487, 
        -49.14091, -49.41337, -49.67056, -49.9109, -50.13463, -50.34291, 
        -50.53764, -50.72034, -50.89188, -51.0535, -51.20563, -51.34888, 
        -51.48431, -51.61253, -51.73425, -51.85011, -51.9598, -52.06588, 
        -52.16771, -52.26569, -52.35998, -52.45042, -52.53688, -52.61934, 
        -52.69761, -52.77232, -52.84328, -52.91104, -52.97618, -53.03919, 
        -53.10033, -53.15979, -53.21583, -53.27084, -53.32333, -53.37379, 
        -53.42284, -53.47119, -53.52005, -53.56976, -53.62077, -53.67344, 
        -53.72756, -53.78278, -53.83789, -53.89258, -53.94606, -53.99844, 
        -54.04926, -54.09774, -54.14573, -54.19236, -54.23768, -54.28211, 
        -54.32618, -54.37074, -54.41587, -54.46217, -54.5099, -54.55919, 
        -54.61011, -54.66215, -54.71513, -54.7685, -54.82186, -54.87479, 
        -54.92699, -54.97716, -55.02724, -55.07624, -55.12386, -55.16975, 
        -55.21412, -55.25692, -55.298, -55.33763, -55.37579, -55.41297, 
        -55.44965, -55.48632, -55.52342, -55.56094, -55.5993, -55.63882, 
        -55.68006, -55.72277, -55.76917, -55.81936, -55.87416, -55.93467, 
        -56.00138, -56.0742, -56.15295, -56.23608, -56.3222, -56.40954, 
        -56.49605, -56.58055, -56.66184, -56.73896, -56.81201, -56.88078, 
        -56.94613, -57.0087, -57.06916, -57.12712, -57.18446, -57.24035, 
        -57.29458, -57.34691, -57.3973, -57.44527, -57.49181, -57.53753, 
        -57.58286, -57.6288, -57.67479, -57.72097, -57.76663, -57.81128, 
        -57.85537, -57.89893, -57.94212, -57.98473, -58.02675, -58.06799, 
        -58.10891, -58.14894, -58.19072, -58.23326, -58.27661, -58.32091, 
        -58.36534, -58.411, -58.45818, -58.50672, -58.55703, -58.60875, 
        -58.66102, -58.71372, -58.76653, -58.81957, -58.87247, -58.9258, 
        -58.97948, -59.03377, -59.0886, -59.14405, -59.19991, -59.25594, 
        -59.31092, -59.36658, -59.42152, -59.47557, -59.52819, -59.57919, 
        -59.62875, -59.67707, -59.72403, -59.7692, -59.81227, -59.85307, 
        -59.89198, -59.92924, -59.96498, -59.99937, -60.03224, -60.06352, 
        -60.09289, -60.11987, -60.14417, -60.16579, -60.18544, -60.20349, 
        -60.22037, -60.23611, -60.24917, -60.26104, -60.27016, -60.27641, 
        -60.27937, -60.27915, -60.27599, -60.27, -60.26182, -60.25167, 
        -60.2395, -60.22516, -60.20883, -60.19103, -60.17127, -60.14957, 
        -60.12607, -60.10038, -60.0723, -60.0418, -60.0088, -59.97311, 
        -59.93449, -59.89292, -59.8486, -59.80159, -59.75232, -59.7007, 
        -59.64647, -59.58928, -59.52783, -59.46424, -59.39824, -59.33055, 
        -59.26164, -59.19232, -59.12315, -59.05388, -58.98448, -58.91499, 
        -58.84495, -58.77435, -58.70284, -58.63027, -58.55675, -58.48201, 
        -58.40613, -58.32919, -58.2514, -58.17323, -58.09453, -58.0157, 
        -57.93682, -57.85797, -57.77926, -57.70035, -57.62138, -57.54227, 
        -57.46292, -57.38353, -57.30424, -57.22519, -57.14615, -57.06689, 
        -56.98743, -56.9067, -56.82681, -56.74696, -56.66737, -56.58867, 
        -56.5108, -56.43412, -56.35841, -56.28325, -56.20826, -56.13321, 
        -56.05826, -55.98385, -55.91056, -55.83893, -55.76937, -55.70219, 
        -55.6374, -55.57528, -55.51515, -55.45671, -55.3995, -55.34357, 
        -55.28862, -55.23464, -55.18182, -55.13056, -55.08105, -55.03368, 
        -54.98798, -54.94389, -54.90171, -54.86222, -54.8259, -54.79332, 
        -54.76431, -54.7385, -54.71547, -54.69497, -54.67656, -54.66004, 
        -54.64498,
  -47.68504, -47.55705, -47.42368, -47.29376, -47.17342, -47.07183, 
        -46.99782, -46.95932, -46.96262, -47.01267, -47.1119, -47.26052, 
        -47.45507, -47.688, -47.95275, -48.23882, -48.53633, -48.83616, 
        -49.13068, -49.41393, -49.68233, -49.93386, -50.1694, -50.38924, 
        -50.595, -50.78762, -50.9685, -51.13832, -51.29705, -51.44753, 
        -51.58969, -51.7243, -51.8522, -51.97411, -52.09063, -52.20237, 
        -52.30954, -52.41267, -52.51176, -52.60643, -52.69674, -52.78224, 
        -52.86339, -52.94104, -53.01418, -53.08545, -53.15457, -53.22142, 
        -53.28638, -53.34919, -53.40954, -53.46744, -53.52253, -53.57529, 
        -53.62638, -53.67672, -53.72747, -53.7792, -53.83257, -53.88749, 
        -53.94413, -54.00119, -54.0597, -54.1179, -54.17479, -54.23039, 
        -54.28453, -54.33741, -54.38872, -54.43879, -54.4875, -54.53532, 
        -54.58268, -54.63018, -54.67818, -54.72704, -54.77685, -54.82806, 
        -54.87931, -54.93235, -54.98613, -55.0401, -55.09407, -55.14768, 
        -55.20074, -55.25329, -55.30478, -55.35564, -55.40557, -55.45437, 
        -55.502, -55.54833, -55.59315, -55.63679, -55.67927, -55.72054, 
        -55.75994, -55.79982, -55.83932, -55.87865, -55.91815, -55.95793, 
        -55.99881, -56.04142, -56.08649, -56.13454, -56.18676, -56.24398, 
        -56.30747, -56.37753, -56.45374, -56.53515, -56.62043, -56.70773, 
        -56.79508, -56.88085, -56.96241, -57.04122, -57.11588, -57.18647, 
        -57.25355, -57.31763, -57.37964, -57.43996, -57.49873, -57.55595, 
        -57.61127, -57.66459, -57.71566, -57.76457, -57.81203, -57.85829, 
        -57.90439, -57.95093, -57.99764, -58.04425, -58.09013, -58.13425, 
        -58.17864, -58.2226, -58.26624, -58.30936, -58.35207, -58.39423, 
        -58.43654, -58.47944, -58.52293, -58.56743, -58.61276, -58.65845, 
        -58.70444, -58.75094, -58.79858, -58.84721, -58.89712, -58.94815, 
        -58.9994, -59.05096, -59.10228, -59.15242, -59.20369, -59.25543, 
        -59.30794, -59.36147, -59.41609, -59.47175, -59.52827, -59.58532, 
        -59.6426, -59.69975, -59.75628, -59.8115, -59.86504, -59.91671, 
        -59.96665, -60.01504, -60.06169, -60.10629, -60.14826, -60.1877, 
        -60.225, -60.26059, -60.29491, -60.32806, -60.35893, -60.3893, 
        -60.41778, -60.44383, -60.4673, -60.48851, -60.50804, -60.52611, 
        -60.54335, -60.55968, -60.57407, -60.58628, -60.59563, -60.60178, 
        -60.60441, -60.60344, -60.59911, -60.59144, -60.58142, -60.56936, 
        -60.5556, -60.54009, -60.52286, -60.50461, -60.4849, -60.46359, 
        -60.4403, -60.41453, -60.38623, -60.35447, -60.3213, -60.28562, 
        -60.24715, -60.20604, -60.16238, -60.1166, -60.0689, -60.01921, 
        -59.96726, -59.91249, -59.85451, -59.79335, -59.7293, -59.66318, 
        -59.59565, -59.52734, -59.45872, -59.38984, -59.32078, -59.25142, 
        -59.18149, -59.11083, -59.03916, -58.96604, -58.89161, -58.81579, 
        -58.73841, -58.65984, -58.58044, -58.50052, -58.42019, -58.33979, 
        -58.25835, -58.17806, -58.09787, -58.01778, -57.93778, -57.85778, 
        -57.77787, -57.69812, -57.61848, -57.53856, -57.45837, -57.37766, 
        -57.29636, -57.21472, -57.13284, -57.05083, -56.9691, -56.88788, 
        -56.80769, -56.72876, -56.65079, -56.57372, -56.49699, -56.42049, 
        -56.34422, -56.26846, -56.19374, -56.12054, -56.04934, -55.98056, 
        -55.91428, -55.85096, -55.78948, -55.73034, -55.67231, -55.61528, 
        -55.55929, -55.50425, -55.45044, -55.39828, -55.348, -55.29877, 
        -55.25232, -55.20777, -55.16493, -55.12449, -55.08718, -55.05343, 
        -55.02321, -54.99634, -54.9722, -54.95048, -54.93086, -54.91294, 
        -54.89616,
  -47.60523, -47.46841, -47.33127, -47.20113, -47.08566, -46.99323, 
        -46.93077, -46.90443, -46.91824, -46.97717, -47.08219, -47.23287, 
        -47.4267, -47.65909, -47.92295, -48.20997, -48.51083, -48.81675, 
        -49.1195, -49.41299, -49.69284, -49.95667, -50.2045, -50.43562, 
        -50.65254, -50.85549, -51.04541, -51.22347, -51.39047, -51.54797, 
        -51.69716, -51.83849, -51.97299, -52.10132, -52.22412, -52.34196, 
        -52.45499, -52.56362, -52.66664, -52.76583, -52.8602, -52.9493, 
        -53.03394, -53.11442, -53.19189, -53.26706, -53.33995, -53.41088, 
        -53.47978, -53.54626, -53.60992, -53.67072, -53.72866, -53.7842, 
        -53.83786, -53.88963, -53.9427, -53.99677, -54.05227, -54.10961, 
        -54.16872, -54.22933, -54.29067, -54.35179, -54.41188, -54.47068, 
        -54.52808, -54.584, -54.63868, -54.69186, -54.74385, -54.79502, 
        -54.8446, -54.89498, -54.94566, -54.99702, -55.04914, -55.10212, 
        -55.15572, -55.20988, -55.26439, -55.31912, -55.37395, -55.42846, 
        -55.48262, -55.53656, -55.58997, -55.64304, -55.6955, -55.74719, 
        -55.79702, -55.84675, -55.89526, -55.9428, -55.98887, -56.0342, 
        -56.07835, -56.12149, -56.16355, -56.20483, -56.24578, -56.28664, 
        -56.32819, -56.37067, -56.41502, -56.46199, -56.512, -56.56718, 
        -56.62782, -56.6936, -56.76694, -56.84611, -56.92996, -57.01655, 
        -57.10378, -57.18998, -57.27354, -57.3536, -57.42952, -57.50142, 
        -57.56992, -57.63551, -57.69897, -57.76057, -57.82063, -57.87902, 
        -57.93559, -57.99015, -58.04204, -58.09036, -58.138, -58.18465, 
        -58.23111, -58.27774, -58.32446, -58.37112, -58.41712, -58.46261, 
        -58.50756, -58.55215, -58.59653, -58.6405, -58.68412, -58.72761, 
        -58.77155, -58.81634, -58.86206, -58.90863, -58.95576, -59.0032, 
        -59.05067, -59.09753, -59.1457, -59.1945, -59.24404, -59.29417, 
        -59.34456, -59.39497, -59.44524, -59.49526, -59.54545, -59.59602, 
        -59.64739, -59.69992, -59.75379, -59.80903, -59.86548, -59.92263, 
        -59.98029, -60.03799, -60.09513, -60.15082, -60.20473, -60.25661, 
        -60.30651, -60.3537, -60.39982, -60.4435, -60.4843, -60.52228, 
        -60.55817, -60.59225, -60.62522, -60.65696, -60.68743, -60.7164, 
        -60.74347, -60.76836, -60.79099, -60.81162, -60.83068, -60.84876, 
        -60.86554, -60.88184, -60.89602, -60.90783, -60.9167, -60.92226, 
        -60.92413, -60.92213, -60.91636, -60.90715, -60.89423, -60.88019, 
        -60.86452, -60.84756, -60.82952, -60.8107, -60.79084, -60.7695, 
        -60.74611, -60.72005, -60.69135, -60.66011, -60.62648, -60.59061, 
        -60.55235, -60.51183, -60.46905, -60.42457, -60.37863, -60.33113, 
        -60.2817, -60.22949, -60.17413, -60.11566, -60.05418, -59.99052, 
        -59.92512, -59.85847, -59.79108, -59.72335, -59.65512, -59.58552, 
        -59.51626, -59.44623, -59.37487, -59.30199, -59.22713, -59.15072, 
        -59.07242, -58.99266, -58.91186, -58.83043, -58.74851, -58.66669, 
        -58.5848, -58.50301, -58.4213, -58.33969, -58.25832, -58.1773, 
        -58.09683, -58.01673, -57.93664, -57.85615, -57.77484, -57.69269, 
        -57.60981, -57.52645, -57.44284, -57.35911, -57.27554, -57.19246, 
        -57.1103, -57.0292, -56.94936, -56.87032, -56.79192, -56.71394, 
        -56.63638, -56.55834, -56.48218, -56.40734, -56.33442, -56.264, 
        -56.19644, -56.13181, -56.06968, -56.00953, -55.95079, -55.89305, 
        -55.83619, -55.78024, -55.72543, -55.67214, -55.62077, -55.57158, 
        -55.52459, -55.47976, -55.4366, -55.39581, -55.35785, -55.32316, 
        -55.29179, -55.26335, -55.23767, -55.21436, -55.19312, -55.1736, 
        -55.15485,
  -47.53318, -47.38988, -47.25053, -47.12199, -47.01379, -46.93169, 
        -46.88103, -46.8671, -46.89241, -46.95926, -47.06821, -47.21913, 
        -47.41068, -47.63953, -47.89983, -48.18562, -48.4879, -48.79726, 
        -49.10769, -49.41103, -49.70233, -49.97918, -50.23982, -50.48425, 
        -50.71276, -50.92603, -51.12507, -51.31119, -51.48567, -51.65016, 
        -51.80595, -51.95422, -52.09566, -52.22974, -52.35917, -52.48339, 
        -52.60273, -52.71718, -52.82657, -52.93064, -53.02935, -53.12236, 
        -53.21079, -53.29503, -53.37617, -53.45494, -53.53175, -53.6068, 
        -53.6797, -53.74906, -53.81638, -53.88035, -53.94129, -53.99979, 
        -54.05654, -54.11228, -54.16806, -54.22461, -54.28258, -54.34219, 
        -54.40363, -54.4666, -54.53059, -54.59437, -54.65727, -54.71784, 
        -54.77806, -54.83683, -54.89436, -54.95066, -55.00591, -55.06002, 
        -55.11364, -55.16702, -55.22047, -55.27427, -55.32842, -55.38291, 
        -55.43785, -55.49303, -55.54848, -55.60404, -55.65985, -55.71462, 
        -55.77007, -55.82557, -55.88075, -55.93604, -55.99105, -56.0456, 
        -56.09933, -56.15247, -56.20454, -56.25562, -56.30563, -56.35455, 
        -56.40211, -56.44849, -56.49356, -56.53743, -56.58044, -56.62283, 
        -56.66443, -56.70774, -56.7523, -56.79881, -56.84778, -56.90112, 
        -56.95934, -57.02347, -57.09404, -57.17064, -57.25243, -57.33765, 
        -57.42419, -57.51022, -57.594, -57.67471, -57.75169, -57.82485, 
        -57.89456, -57.96041, -58.02491, -58.08762, -58.14883, -58.20855, 
        -58.2662, -58.32144, -58.37387, -58.42366, -58.47153, -58.51836, 
        -58.56495, -58.61139, -58.65791, -58.70433, -58.75039, -58.79624, 
        -58.84196, -58.88747, -58.93275, -58.97774, -59.02262, -59.06661, 
        -59.11235, -59.15912, -59.20692, -59.25554, -59.3046, -59.35375, 
        -59.40277, -59.4517, -59.50058, -59.5496, -59.59885, -59.6483, 
        -59.69792, -59.7479, -59.79705, -59.84682, -59.89656, -59.94638, 
        -59.99688, -60.04839, -60.1012, -60.15533, -60.20969, -60.26596, 
        -60.32275, -60.37972, -60.43623, -60.49146, -60.54502, -60.59653, 
        -60.64605, -60.69365, -60.73883, -60.78152, -60.82119, -60.85809, 
        -60.89268, -60.92543, -60.95696, -60.98718, -61.01598, -61.04318, 
        -61.06849, -61.09188, -61.1134, -61.13326, -61.15177, -61.16895, 
        -61.18421, -61.19932, -61.21221, -61.22293, -61.23043, -61.23473, 
        -61.23553, -61.23243, -61.22538, -61.21478, -61.20132, -61.18573, 
        -61.16861, -61.1505, -61.1315, -61.11203, -61.09163, -61.06982, 
        -61.04572, -61.019, -60.98965, -60.95786, -60.92382, -60.88762, 
        -60.84932, -60.8091, -60.76719, -60.72396, -60.67971, -60.63315, 
        -60.58585, -60.53607, -60.48325, -60.42739, -60.36868, -60.30768, 
        -60.24486, -60.18063, -60.11532, -60.04915, -59.98247, -59.91528, 
        -59.84745, -59.77871, -59.70852, -59.63649, -59.56225, -59.48573, 
        -59.40714, -59.32674, -59.24509, -59.16254, -59.07944, -58.99611, 
        -58.91294, -58.82983, -58.74673, -58.66365, -58.58083, -58.49859, 
        -58.41722, -58.33652, -58.25591, -58.17474, -58.09147, -58.00814, 
        -57.92399, -57.83919, -57.75411, -57.66895, -57.58381, -57.49924, 
        -57.41557, -57.33298, -57.25153, -57.17093, -57.09106, -57.01179, 
        -56.93298, -56.85469, -56.77725, -56.7009, -56.62641, -56.55453, 
        -56.48566, -56.41997, -56.35681, -56.29575, -56.23626, -56.1778, 
        -56.1201, -56.06334, -56.00769, -55.95351, -55.90128, -55.85118, 
        -55.80376, -55.75886, -55.71579, -55.67507, -55.63678, -55.60137, 
        -55.56878, -55.53888, -55.51137, -55.48599, -55.46268, -55.44099, 
        -55.42023,
  -47.47217, -47.32463, -47.18516, -47.06231, -46.96275, -46.89157, 
        -46.85313, -46.85056, -46.88514, -46.95803, -47.06944, -47.21904, 
        -47.40546, -47.62891, -47.88411, -48.16661, -48.46887, -48.78262, 
        -49.09945, -49.41235, -49.71532, -50.00455, -50.27813, -50.53505, 
        -50.77505, -50.99844, -51.20643, -51.39949, -51.58136, -51.75283, 
        -51.91552, -52.07075, -52.21925, -52.36136, -52.49762, -52.6287, 
        -52.75449, -52.87504, -52.99023, -53.09964, -53.20308, -53.3008, 
        -53.39338, -53.48077, -53.566, -53.64888, -53.7298, -53.80888, 
        -53.88591, -53.95991, -54.03093, -54.09871, -54.16311, -54.2248, 
        -54.28462, -54.34349, -54.40231, -54.46164, -54.52226, -54.58347, 
        -54.64726, -54.71263, -54.77879, -54.84488, -54.91037, -54.97432, 
        -55.03672, -55.09799, -55.15829, -55.21724, -55.27527, -55.33261, 
        -55.38894, -55.44519, -55.50108, -55.55708, -55.61302, -55.66814, 
        -55.72437, -55.78043, -55.83679, -55.89358, -55.95067, -56.0079, 
        -56.06504, -56.12207, -56.17925, -56.23648, -56.29377, -56.35063, 
        -56.40709, -56.46331, -56.51851, -56.57304, -56.6266, -56.67806, 
        -56.72928, -56.77915, -56.82746, -56.87415, -56.91971, -56.96432, 
        -57.0087, -57.05336, -57.09853, -57.14516, -57.19398, -57.24619, 
        -57.30283, -57.36478, -57.43287, -57.50709, -57.58667, -57.67021, 
        -57.75426, -57.83944, -57.92309, -58.00413, -58.08179, -58.15574, 
        -58.2262, -58.29393, -58.35917, -58.42265, -58.48453, -58.54509, 
        -58.6037, -58.65975, -58.713, -58.76316, -58.81146, -58.85863, 
        -58.90527, -58.95169, -58.99791, -59.04308, -59.08925, -59.13556, 
        -59.18211, -59.22857, -59.27513, -59.32148, -59.36784, -59.41455, 
        -59.46207, -59.51093, -59.56059, -59.61111, -59.66191, -59.71251, 
        -59.76272, -59.81257, -59.86211, -59.91141, -59.96056, -60.00962, 
        -60.05912, -60.10678, -60.15618, -60.20599, -60.25565, -60.30518, 
        -60.35497, -60.4054, -60.45673, -60.5091, -60.56239, -60.61659, 
        -60.67165, -60.72636, -60.78119, -60.83476, -60.88701, -60.93753, 
        -60.98618, -61.03271, -61.07695, -61.11853, -61.15718, -61.19305, 
        -61.22663, -61.25826, -61.2875, -61.31611, -61.34306, -61.36831, 
        -61.39157, -61.41308, -61.43316, -61.45187, -61.46935, -61.4856, 
        -61.50048, -61.51356, -61.52469, -61.53341, -61.53911, -61.54173, 
        -61.54089, -61.53626, -61.52794, -61.51624, -61.50171, -61.48504, 
        -61.46687, -61.44773, -61.42796, -61.40764, -61.38638, -61.36353, 
        -61.33746, -61.30986, -61.27964, -61.24715, -61.21249, -61.17594, 
        -61.1375, -61.09752, -61.05614, -61.01384, -60.97085, -60.92692, 
        -60.88138, -60.83361, -60.78278, -60.72913, -60.67295, -60.61478, 
        -60.55486, -60.49334, -60.4304, -60.36646, -60.30189, -60.23684, 
        -60.17085, -60.10392, -60.03547, -59.96489, -59.8919, -59.81618, 
        -59.73807, -59.65784, -59.57492, -59.49178, -59.40782, -59.32362, 
        -59.23943, -59.15525, -59.07095, -58.98651, -58.90231, -58.81886, 
        -58.73645, -58.6549, -58.57353, -58.4916, -58.40854, -58.32434, 
        -58.2391, -58.15323, -58.06697, -57.98058, -57.89422, -57.80855, 
        -57.72379, -57.64006, -57.55741, -57.47574, -57.39479, -57.3144, 
        -57.23452, -57.15509, -57.07634, -56.99875, -56.92291, -56.8497, 
        -56.77954, -56.7124, -56.6481, -56.58617, -56.52586, -56.46666, 
        -56.40817, -56.34975, -56.29333, -56.23846, -56.18564, -56.13533, 
        -56.08777, -56.04285, -56.00024, -55.95977, -55.92134, -55.88525, 
        -55.85165, -55.82016, -55.7908, -55.76342, -55.73794, -55.71411, 
        -55.69126,
  -47.42846, -47.27889, -47.14169, -47.02431, -46.93339, -46.87293, 
        -46.84587, -46.85244, -46.89506, -46.97252, -47.08495, -47.23206, 
        -47.41404, -47.63063, -47.87967, -48.15751, -48.45817, -48.77385, 
        -49.09643, -49.41796, -49.73202, -50.0334, -50.31828, -50.58707, 
        -50.83822, -51.07172, -51.28845, -51.49038, -51.6796, -51.85824, 
        -52.02803, -52.19044, -52.34612, -52.49556, -52.63907, -52.77713, 
        -52.9097, -53.03555, -53.1566, -53.27154, -53.38025, -53.48302, 
        -53.58061, -53.67378, -53.76377, -53.85124, -53.93659, -54.01978, 
        -54.10081, -54.17896, -54.25388, -54.32512, -54.39307, -54.45738, 
        -54.52058, -54.58269, -54.64467, -54.70699, -54.77046, -54.83538, 
        -54.90186, -54.96946, -55.03766, -55.10587, -55.17342, -55.23947, 
        -55.30392, -55.36712, -55.42946, -55.49096, -55.55072, -55.61053, 
        -55.66954, -55.72799, -55.78609, -55.84393, -55.90165, -55.95906, 
        -56.01643, -56.07375, -56.13137, -56.18952, -56.24816, -56.30714, 
        -56.36601, -56.42492, -56.48388, -56.54284, -56.60096, -56.66004, 
        -56.71893, -56.77761, -56.83574, -56.89341, -56.9504, -57.00647, 
        -57.06142, -57.11474, -57.16642, -57.21638, -57.26481, -57.31216, 
        -57.35866, -57.40498, -57.45152, -57.49893, -57.54811, -57.59888, 
        -57.65459, -57.71523, -57.78154, -57.85372, -57.93107, -58.01244, 
        -58.096, -58.18, -58.26298, -58.34358, -58.42121, -58.49542, 
        -58.56624, -58.63416, -58.69959, -58.76342, -58.826, -58.88729, 
        -58.94681, -59.00271, -59.05674, -59.10795, -59.1571, -59.20497, 
        -59.25195, -59.29847, -59.34468, -59.39083, -59.43718, -59.48388, 
        -59.53115, -59.57887, -59.62683, -59.67484, -59.7229, -59.77139, 
        -59.82078, -59.87133, -59.92288, -59.97497, -60.02709, -60.07778, 
        -60.12889, -60.17943, -60.22951, -60.27914, -60.32842, -60.37745, 
        -60.42641, -60.47549, -60.525, -60.57479, -60.62439, -60.6736, 
        -60.72255, -60.77163, -60.82114, -60.87121, -60.92182, -60.97296, 
        -61.02458, -61.07645, -61.12824, -61.17941, -61.22937, -61.27692, 
        -61.32387, -61.36898, -61.41192, -61.45231, -61.49003, -61.52514, 
        -61.55796, -61.58881, -61.61782, -61.645, -61.67018, -61.69334, 
        -61.7146, -61.7342, -61.75248, -61.7696, -61.7855, -61.80006, 
        -61.81298, -61.82394, -61.83261, -61.83874, -61.84209, -61.84243, 
        -61.83958, -61.83237, -61.82283, -61.81019, -61.79489, -61.77752, 
        -61.75865, -61.73874, -61.71812, -61.69678, -61.67437, -61.6503, 
        -61.62401, -61.59526, -61.56406, -61.53068, -61.49535, -61.45827, 
        -61.41966, -61.37966, -61.33867, -61.29702, -61.25486, -61.21202, 
        -61.16768, -61.1212, -61.07205, -61.02025, -60.96625, -60.9104, 
        -60.85303, -60.79421, -60.73304, -60.67179, -60.60967, -60.54688, 
        -60.48331, -60.4186, -60.35222, -60.28349, -60.2121, -60.13791, 
        -60.061, -59.98167, -59.90017, -59.81712, -59.73306, -59.64853, 
        -59.56383, -59.47888, -59.39363, -59.30813, -59.22281, -59.13825, 
        -59.05477, -58.97225, -58.89005, -58.80735, -58.72362, -58.63869, 
        -58.55276, -58.46611, -58.37892, -58.29147, -58.20413, -58.11748, 
        -58.03187, -57.9474, -57.864, -57.78051, -57.69876, -57.61758, 
        -57.53682, -57.45643, -57.37663, -57.29795, -57.22105, -57.1466, 
        -57.07506, -57.00661, -56.94105, -56.87793, -56.81668, -56.7567, 
        -56.6977, -56.63967, -56.58282, -56.52765, -56.47467, -56.42437, 
        -56.3769, -56.33214, -56.28976, -56.2494, -56.21094, -56.17439, 
        -56.13977, -56.10702, -56.07607, -56.04689, -56.01939, -55.99332, 
        -55.96818,
  -47.4047, -47.25433, -47.12117, -47.01077, -46.92882, -46.87854, 
        -46.86141, -46.87758, -46.92623, -47.00658, -47.11839, -47.26178, 
        -47.4374, -47.64614, -47.88766, -48.15967, -48.45657, -48.77293, 
        -49.09986, -49.4291, -49.75309, -50.0656, -50.36304, -50.64291, 
        -50.90451, -51.14756, -51.3731, -51.58301, -51.77989, -51.96585, 
        -52.14299, -52.31169, -52.4748, -52.63175, -52.78288, -52.92804, 
        -53.06756, -53.20082, -53.3279, -53.44864, -53.56312, -53.67148, 
        -53.77457, -53.87318, -53.96819, -54.06062, -54.15067, -54.23758, 
        -54.3225, -54.40461, -54.48339, -54.55842, -54.6304, -54.69952, 
        -54.76653, -54.83208, -54.89727, -54.96276, -55.02927, -55.09695, 
        -55.166, -55.23615, -55.30652, -55.37658, -55.44473, -55.51262, 
        -55.5789, -55.64398, -55.70786, -55.77148, -55.83423, -55.89605, 
        -55.95721, -56.01791, -56.0778, -56.13712, -56.19595, -56.2544, 
        -56.3129, -56.37154, -56.43079, -56.49046, -56.55003, -56.61104, 
        -56.67193, -56.73275, -56.7934, -56.85405, -56.91477, -56.97548, 
        -57.03612, -57.09708, -57.15797, -57.21864, -57.27903, -57.33857, 
        -57.39702, -57.45393, -57.50902, -57.56231, -57.61279, -57.66298, 
        -57.71219, -57.76076, -57.80906, -57.8577, -57.90786, -57.9601, 
        -58.0158, -58.07594, -58.14095, -58.21128, -58.28653, -58.36574, 
        -58.44743, -58.52999, -58.61185, -58.69182, -58.76913, -58.84303, 
        -58.91236, -58.97976, -59.04488, -59.10874, -59.17173, -59.23341, 
        -59.2935, -59.35131, -59.40656, -59.45872, -59.50913, -59.55816, 
        -59.60608, -59.65319, -59.69975, -59.74625, -59.79296, -59.84026, 
        -59.8886, -59.93766, -59.98713, -60.0357, -60.08559, -60.13599, 
        -60.18711, -60.23938, -60.2924, -60.34588, -60.39898, -60.45124, 
        -60.50272, -60.55352, -60.60395, -60.65368, -60.70317, -60.75243, 
        -60.80176, -60.8511, -60.90094, -60.95093, -61.0004, -61.04909, 
        -61.09705, -61.14455, -61.19085, -61.23801, -61.28516, -61.33232, 
        -61.37962, -61.42728, -61.47511, -61.52297, -61.56967, -61.61561, 
        -61.66023, -61.70337, -61.74441, -61.78339, -61.82028, -61.8548, 
        -61.88717, -61.91748, -61.94566, -61.97173, -61.99541, -62.01671, 
        -62.03571, -62.0532, -62.06964, -62.08423, -62.09822, -62.11082, 
        -62.12146, -62.12976, -62.13551, -62.13861, -62.13912, -62.13676, 
        -62.13157, -62.12342, -62.11267, -62.09935, -62.08366, -62.06598, 
        -62.04671, -62.02615, -62.00463, -61.9821, -61.95822, -61.93261, 
        -61.9048, -61.87475, -61.84249, -61.80827, -61.77219, -61.73462, 
        -61.69564, -61.65568, -61.61394, -61.57272, -61.53101, -61.4887, 
        -61.44498, -61.39917, -61.35085, -61.30006, -61.24748, -61.19355, 
        -61.13842, -61.08202, -61.02427, -60.96545, -60.90604, -60.84565, 
        -60.78477, -60.72258, -60.65851, -60.5921, -60.52277, -60.45077, 
        -60.37577, -60.29798, -60.21764, -60.13534, -60.0518, -59.96764, 
        -59.88299, -59.79775, -59.71184, -59.6256, -59.53941, -59.45396, 
        -59.36954, -59.28502, -59.20189, -59.11834, -59.03392, -58.94853, 
        -58.86219, -58.77501, -58.68707, -58.59874, -58.51059, -58.42319, 
        -58.33701, -58.25209, -58.16829, -58.08527, -58.00288, -57.92096, 
        -57.83931, -57.75816, -57.67741, -57.59797, -57.52034, -57.44501, 
        -57.37235, -57.30269, -57.2359, -57.17163, -57.10945, -57.04873, 
        -56.98911, -56.93061, -56.87334, -56.81798, -56.765, -56.71482, 
        -56.6675, -56.62289, -56.58066, -56.54038, -56.50182, -56.46486, 
        -56.42948, -56.39564, -56.36338, -56.33158, -56.30226, -56.27413, 
        -56.24702,
  -47.40077, -47.25337, -47.12498, -47.02199, -46.94915, -46.9086, 
        -46.90062, -46.92405, -46.97742, -47.05927, -47.16933, -47.30707, 
        -47.47551, -47.67596, -47.9095, -48.1748, -48.46872, -48.78468, 
        -49.11455, -49.44938, -49.78176, -50.10401, -50.4115, -50.70152, 
        -50.97258, -51.22452, -51.45763, -51.67577, -51.8806, -52.07436, 
        -52.25948, -52.43708, -52.60812, -52.77301, -52.93182, -53.08427, 
        -53.23067, -53.37041, -53.50351, -53.63017, -53.75042, -53.86478, 
        -53.97283, -54.07722, -54.17818, -54.27605, -54.37133, -54.46407, 
        -54.5539, -54.64009, -54.72263, -54.80151, -54.87735, -54.95039, 
        -55.02141, -55.09067, -55.15929, -55.22791, -55.29643, -55.36714, 
        -55.43892, -55.51143, -55.58391, -55.65557, -55.72615, -55.79541, 
        -55.86335, -55.92992, -55.99541, -56.06031, -56.1246, -56.18805, 
        -56.25074, -56.31297, -56.37416, -56.43374, -56.49363, -56.55327, 
        -56.61294, -56.67306, -56.73396, -56.79581, -56.85845, -56.9215, 
        -56.98448, -57.04722, -57.10994, -57.17205, -57.23401, -57.29589, 
        -57.3583, -57.42135, -57.48456, -57.54717, -57.61063, -57.67347, 
        -57.73542, -57.79592, -57.85428, -57.91085, -57.96553, -58.01873, 
        -58.07086, -58.12164, -58.17217, -58.22261, -58.27398, -58.32755, 
        -58.38391, -58.44396, -58.50836, -58.57753, -58.65011, -58.72726, 
        -58.80701, -58.88776, -58.96822, -59.04694, -59.12307, -59.19537, 
        -59.26461, -59.3311, -59.39583, -59.4595, -59.52273, -59.58537, 
        -59.64656, -59.70609, -59.76284, -59.81692, -59.86948, -59.92016, 
        -59.96914, -60.01614, -60.06313, -60.10971, -60.15683, -60.20489, 
        -60.25404, -60.30419, -60.35504, -60.40651, -60.45821, -60.51046, 
        -60.56332, -60.61693, -60.67129, -60.72551, -60.77918, -60.83184, 
        -60.88351, -60.93431, -60.98476, -61.03472, -61.08454, -61.13319, 
        -61.18278, -61.23248, -61.28232, -61.33196, -61.38084, -61.4287, 
        -61.4751, -61.52068, -61.56549, -61.60954, -61.65291, -61.69585, 
        -61.73857, -61.78138, -61.82438, -61.8675, -61.9103, -61.95246, 
        -61.99404, -62.0345, -62.07346, -62.1108, -62.14636, -62.1802, 
        -62.21127, -62.24119, -62.26899, -62.29464, -62.31755, -62.33751, 
        -62.35503, -62.37069, -62.38531, -62.3987, -62.41055, -62.42065, 
        -62.42868, -62.43398, -62.43641, -62.43643, -62.43359, -62.42853, 
        -62.42089, -62.41094, -62.39876, -62.38446, -62.36808, -62.34977, 
        -62.33002, -62.30834, -62.28583, -62.26097, -62.23561, -62.20857, 
        -62.17952, -62.14837, -62.11523, -62.08015, -62.04354, -62.00551, 
        -61.96637, -61.92634, -61.88557, -61.84434, -61.80273, -61.76042, 
        -61.71672, -61.67109, -61.62315, -61.57314, -61.52185, -61.46946, 
        -61.41603, -61.36137, -61.3058, -61.24907, -61.19144, -61.13352, 
        -61.07517, -61.01523, -60.95332, -60.88891, -60.82172, -60.75065, 
        -60.67777, -60.60187, -60.5233, -60.44246, -60.36016, -60.27685, 
        -60.19275, -60.10775, -60.02181, -59.93528, -59.84877, -59.76287, 
        -59.67784, -59.59355, -59.50954, -59.42524, -59.34025, -59.25441, 
        -59.16771, -59.08018, -58.99187, -58.90304, -58.81431, -58.72631, 
        -58.63953, -58.55408, -58.46984, -58.38656, -58.30373, -58.22125, 
        -58.13906, -58.05709, -57.97606, -57.89615, -57.8181, -57.74203, 
        -57.66841, -57.59756, -57.52961, -57.46334, -57.40013, -57.33867, 
        -57.27848, -57.21954, -57.16211, -57.10674, -57.05386, -57.00377, 
        -56.95649, -56.91185, -56.86949, -56.82902, -56.79018, -56.75278, 
        -56.71687, -56.68232, -56.64904, -56.61701, -56.58622, -56.5565, 
        -56.52782,
  -47.41873, -47.27568, -47.15327, -47.05885, -46.99487, -46.96251, 
        -46.96281, -46.99238, -47.0489, -47.13109, -47.23881, -47.37249, 
        -47.53389, -47.72574, -47.95033, -48.208, -48.49599, -48.80951, 
        -49.14054, -49.47923, -49.81661, -50.14686, -50.46302, -50.76162, 
        -51.04104, -51.30127, -51.54391, -51.7707, -51.98404, -52.18652, 
        -52.38024, -52.56625, -52.74557, -52.91868, -53.08516, -53.24517, 
        -53.39731, -53.54344, -53.6827, -53.81513, -53.94143, -54.06168, 
        -54.17683, -54.28764, -54.39462, -54.49858, -54.59962, -54.69785, 
        -54.79262, -54.88337, -54.97007, -55.05324, -55.13215, -55.20917, 
        -55.28415, -55.35741, -55.42961, -55.50158, -55.5741, -55.64762, 
        -55.72204, -55.79677, -55.87112, -55.94433, -56.01623, -56.08659, 
        -56.15584, -56.22373, -56.29042, -56.35533, -56.42066, -56.48508, 
        -56.54902, -56.61213, -56.67458, -56.73597, -56.79679, -56.85743, 
        -56.91836, -56.97993, -57.04278, -57.10675, -57.1718, -57.23703, 
        -57.30216, -57.36702, -57.43158, -57.49459, -57.55774, -57.62119, 
        -57.68465, -57.74929, -57.81499, -57.88105, -57.9476, -58.01349, 
        -58.07851, -58.14215, -58.20383, -58.26361, -58.32161, -58.3777, 
        -58.43257, -58.48618, -58.53908, -58.59087, -58.64386, -58.69876, 
        -58.75634, -58.81702, -58.88161, -58.94997, -59.02216, -59.09756, 
        -59.17556, -59.25454, -59.33315, -59.41007, -59.484, -59.55465, 
        -59.62199, -59.68694, -59.75084, -59.8144, -59.87821, -59.94089, 
        -60.00365, -60.06496, -60.12378, -60.18065, -60.23546, -60.28813, 
        -60.33893, -60.38792, -60.43569, -60.48286, -60.53038, -60.57911, 
        -60.62908, -60.68017, -60.73231, -60.78522, -60.83856, -60.89227, 
        -60.94666, -61.00165, -61.05672, -61.11057, -61.16457, -61.21739, 
        -61.26905, -61.31984, -61.36994, -61.41993, -61.46988, -61.51984, 
        -61.56982, -61.61972, -61.66925, -61.71795, -61.76578, -61.81198, 
        -61.85659, -61.89999, -61.94201, -61.98267, -62.02208, -62.0606, 
        -62.0985, -62.13604, -62.17364, -62.21034, -62.24817, -62.28603, 
        -62.32378, -62.36072, -62.39682, -62.43202, -62.46574, -62.49875, 
        -62.53086, -62.56089, -62.58899, -62.61446, -62.63689, -62.65621, 
        -62.67274, -62.6871, -62.69983, -62.71105, -62.72058, -62.72818, 
        -62.73282, -62.7349, -62.7342, -62.731, -62.72506, -62.71599, 
        -62.70592, -62.69405, -62.68044, -62.66502, -62.64785, -62.62871, 
        -62.60748, -62.58518, -62.56117, -62.53569, -62.50895, -62.48059, 
        -62.45041, -62.41835, -62.38447, -62.34887, -62.31179, -62.2735, 
        -62.23423, -62.19426, -62.15359, -62.11227, -62.0704, -62.02756, 
        -61.98345, -61.93753, -61.88972, -61.84018, -61.78951, -61.73705, 
        -61.68467, -61.63124, -61.57686, -61.52146, -61.46572, -61.40971, 
        -61.35312, -61.29493, -61.23468, -61.17199, -61.10674, -61.03863, 
        -60.96772, -60.89376, -60.81725, -60.73846, -60.65802, -60.5761, 
        -60.49295, -60.40856, -60.32318, -60.23707, -60.15098, -60.06521, 
        -59.98001, -59.89524, -59.81052, -59.72548, -59.63983, -59.5536, 
        -59.46671, -59.3791, -59.29074, -59.20181, -59.11279, -59.02326, 
        -58.93579, -58.84968, -58.76493, -58.68122, -58.59814, -58.5154, 
        -58.43293, -58.35096, -58.26984, -58.18998, -58.11167, -58.03521, 
        -57.96094, -57.88917, -57.82009, -57.7538, -57.68972, -57.62753, 
        -57.56676, -57.50742, -57.4498, -57.39442, -57.34159, -57.29141, 
        -57.24399, -57.19906, -57.15629, -57.11551, -57.07626, -57.03846, 
        -57.002, -56.96683, -56.93281, -56.89982, -56.8678, -56.83673, 
        -56.80659,
  -47.457, -47.31914, -47.20454, -47.11898, -47.06489, -47.04211, 
        -47.0496, -47.08474, -47.14391, -47.22597, -47.33085, -47.4589, 
        -47.61267, -47.79561, -48.01121, -48.25957, -48.5411, -48.85009, 
        -49.1799, -49.52027, -49.86226, -50.19762, -50.51995, -50.82531, 
        -51.11174, -51.37967, -51.63061, -51.86609, -52.08871, -52.30089, 
        -52.5033, -52.69884, -52.88717, -53.06864, -53.24315, -53.41043, 
        -53.5703, -53.72265, -53.86774, -54.00614, -54.13813, -54.26443, 
        -54.38583, -54.50293, -54.61658, -54.72676, -54.83295, -54.93692, 
        -55.03716, -55.13311, -55.22493, -55.31276, -55.39711, -55.47839, 
        -55.55731, -55.6345, -55.71036, -55.78573, -55.86116, -55.93722, 
        -56.0139, -56.09044, -56.16622, -56.24005, -56.31303, -56.38436, 
        -56.4544, -56.52339, -56.59117, -56.65784, -56.72377, -56.78889, 
        -56.85331, -56.91721, -56.9803, -57.04266, -57.10435, -57.16597, 
        -57.22827, -57.29172, -57.3556, -57.42184, -57.48898, -57.55651, 
        -57.62403, -57.69122, -57.75761, -57.82292, -57.88781, -57.95275, 
        -58.01788, -58.08431, -58.15174, -58.22043, -58.28952, -58.35828, 
        -58.42612, -58.49266, -58.55648, -58.61943, -58.68044, -58.73954, 
        -58.79706, -58.85368, -58.90932, -58.96427, -59.01943, -59.07558, 
        -59.1344, -59.19578, -59.26067, -59.3287, -59.39978, -59.47393, 
        -59.55007, -59.62717, -59.70376, -59.77813, -59.84878, -59.91709, 
        -59.98254, -60.04594, -60.10885, -60.17251, -60.23706, -60.30226, 
        -60.36695, -60.4304, -60.49232, -60.55217, -60.60974, -60.66488, 
        -60.71737, -60.76765, -60.8161, -60.86395, -60.91202, -60.96126, 
        -61.01185, -61.06285, -61.11594, -61.17004, -61.22469, -61.27975, 
        -61.3353, -61.39098, -61.44662, -61.50168, -61.55557, -61.60837, 
        -61.65992, -61.71057, -61.76029, -61.80989, -61.85954, -61.90916, 
        -61.95878, -62.00826, -62.05669, -62.1044, -62.15053, -62.19497, 
        -62.23662, -62.2776, -62.31665, -62.35398, -62.38953, -62.42352, 
        -62.45654, -62.48886, -62.52093, -62.55297, -62.58535, -62.61832, 
        -62.6517, -62.68504, -62.7182, -62.75084, -62.78276, -62.81489, 
        -62.84608, -62.87642, -62.90458, -62.92992, -62.95221, -62.97118, 
        -62.98704, -62.99931, -63.01059, -63.01959, -63.02657, -63.03114, 
        -63.03289, -63.03189, -63.02795, -63.02153, -63.01264, -63.00181, 
        -62.98924, -62.97527, -62.95984, -62.94295, -62.92404, -62.9035, 
        -62.88117, -62.85732, -62.83172, -62.80486, -62.77679, -62.74732, 
        -62.71638, -62.68371, -62.64941, -62.6136, -62.57639, -62.53806, 
        -62.49779, -62.45767, -62.41708, -62.37533, -62.3329, -62.28942, 
        -62.24464, -62.19842, -62.15053, -62.1013, -62.05113, -62.00029, 
        -61.94857, -61.89579, -61.84216, -61.78787, -61.73318, -61.67828, 
        -61.62261, -61.56552, -61.50621, -61.44455, -61.38052, -61.31367, 
        -61.24449, -61.17289, -61.0984, -61.02169, -60.9432, -60.86292, 
        -60.78118, -60.69783, -60.61349, -60.52747, -60.44213, -60.35687, 
        -60.27192, -60.18698, -60.10184, -60.01628, -59.93014, -59.84352, 
        -59.75644, -59.66886, -59.58063, -59.49181, -59.40279, -59.31405, 
        -59.22609, -59.13943, -59.05413, -58.9701, -58.88697, -58.8043, 
        -58.72204, -58.6404, -58.5596, -58.48002, -58.40183, -58.32513, 
        -58.25042, -58.17797, -58.10809, -58.04072, -57.97578, -57.91282, 
        -57.85152, -57.79185, -57.73411, -57.67865, -57.62563, -57.57535, 
        -57.52749, -57.48207, -57.43888, -57.39761, -57.35786, -57.31841, 
        -57.2814, -57.24558, -57.21091, -57.17717, -57.14434, -57.11236, 
        -57.08123,
  -47.51368, -47.38316, -47.27761, -47.20266, -47.15821, -47.14521, 
        -47.15996, -47.20018, -47.26182, -47.34392, -47.44471, -47.56763, 
        -47.7142, -47.88833, -48.09452, -48.33485, -48.60803, -48.91068, 
        -49.23624, -49.57527, -49.91805, -50.25594, -50.58212, -50.89229, 
        -51.18468, -51.45816, -51.71708, -51.96173, -52.19439, -52.41698, 
        -52.63081, -52.83673, -53.0349, -53.22549, -53.40816, -53.58284, 
        -53.74925, -53.90769, -54.05849, -54.20216, -54.3387, -54.47071, 
        -54.59809, -54.72149, -54.84167, -54.95861, -55.0723, -55.18245, 
        -55.28879, -55.39069, -55.48807, -55.58123, -55.6707, -55.75669, 
        -55.83979, -55.92085, -56.0002, -56.07789, -56.15634, -56.23466, 
        -56.31311, -56.39103, -56.46811, -56.54372, -56.61775, -56.69004, 
        -56.76079, -56.83045, -56.89876, -56.96611, -57.03218, -57.09774, 
        -57.16249, -57.22685, -57.28962, -57.35261, -57.41516, -57.47795, 
        -57.54171, -57.60691, -57.67377, -57.7422, -57.81166, -57.88151, 
        -57.95126, -58.02051, -58.0888, -58.15598, -58.22262, -58.28923, 
        -58.35642, -58.42463, -58.49332, -58.56419, -58.63545, -58.7066, 
        -58.77709, -58.84638, -58.91394, -58.97963, -59.04339, -59.10554, 
        -59.16615, -59.22534, -59.28362, -59.34076, -59.39779, -59.45578, 
        -59.51575, -59.57791, -59.64297, -59.71003, -59.78072, -59.85363, 
        -59.92818, -60.00338, -60.07761, -60.14964, -60.21863, -60.28452, 
        -60.34766, -60.40977, -60.47226, -60.53592, -60.60128, -60.66786, 
        -60.73472, -60.801, -60.86583, -60.92871, -60.98909, -61.04584, 
        -61.10052, -61.15255, -61.2022, -61.25072, -61.29927, -61.34904, 
        -61.40012, -61.4525, -61.5063, -61.56112, -61.61664, -61.67276, 
        -61.72895, -61.78509, -61.84061, -61.89546, -61.94922, -62.00196, 
        -62.05334, -62.10377, -62.15302, -62.20074, -62.24945, -62.29822, 
        -62.34679, -62.39496, -62.44202, -62.48792, -62.53223, -62.57473, 
        -62.61514, -62.6535, -62.68966, -62.72353, -62.75533, -62.78536, 
        -62.81376, -62.84094, -62.86741, -62.89381, -62.92045, -62.94822, 
        -62.97701, -63.00628, -63.03595, -63.06586, -63.09488, -63.12534, 
        -63.15592, -63.18548, -63.21344, -63.2388, -63.26105, -63.27962, 
        -63.29514, -63.30742, -63.31691, -63.32377, -63.32798, -63.32964, 
        -63.32837, -63.32421, -63.31745, -63.3081, -63.29658, -63.28319, 
        -63.26831, -63.25198, -63.23472, -63.21572, -63.19523, -63.17298, 
        -63.14904, -63.12254, -63.09546, -63.0671, -63.03773, -63.00729, 
        -62.97564, -62.94267, -62.90832, -62.87265, -62.83567, -62.79746, 
        -62.75838, -62.71842, -62.67756, -62.63571, -62.59269, -62.54842, 
        -62.50296, -62.45621, -62.4083, -62.35934, -62.30954, -62.25879, 
        -62.20717, -62.15476, -62.10136, -62.04765, -61.99358, -61.9389, 
        -61.88348, -61.82645, -61.76638, -61.70504, -61.64163, -61.57581, 
        -61.50781, -61.43779, -61.3653, -61.29043, -61.21391, -61.13548, 
        -61.05512, -60.97337, -60.89055, -60.807, -60.72301, -60.63866, 
        -60.55421, -60.46935, -60.38404, -60.2982, -60.21173, -60.12484, 
        -60.03751, -59.94992, -59.86206, -59.77372, -59.68514, -59.59653, 
        -59.5084, -59.42135, -59.33569, -59.25157, -59.16848, -59.08607, 
        -59.00437, -58.92326, -58.84332, -58.76445, -58.68679, -58.60942, 
        -58.53449, -58.46156, -58.39086, -58.32259, -58.25668, -58.19288, 
        -58.13108, -58.07112, -58.01326, -57.9577, -57.90445, -57.85348, 
        -57.80481, -57.75866, -57.71491, -57.67323, -57.63259, -57.59343, 
        -57.5557, -57.51909, -57.48382, -57.4496, -57.41629, -57.38376, 
        -57.35196,
  -47.58758, -47.46626, -47.37141, -47.3073, -47.27319, -47.26993, 
        -47.29214, -47.33725, -47.40128, -47.4831, -47.58218, -47.70037, 
        -47.84053, -48.00654, -48.20331, -48.43396, -48.69811, -48.99254, 
        -49.31136, -49.64482, -49.98516, -50.32232, -50.64947, -50.96211, 
        -51.25892, -51.53952, -51.80565, -52.05956, -52.30287, -52.53678, 
        -52.76223, -52.97948, -53.18843, -53.38875, -53.58002, -53.76106, 
        -53.93399, -54.09804, -54.25409, -54.40267, -54.54509, -54.68245, 
        -54.81551, -54.94494, -55.07138, -55.19504, -55.31557, -55.43254, 
        -55.54536, -55.65378, -55.75756, -55.85576, -55.95083, -56.04214, 
        -56.12987, -56.21484, -56.29762, -56.37922, -56.4603, -56.54078, 
        -56.62059, -56.6998, -56.77773, -56.85426, -56.9291, -57.00212, 
        -57.07358, -57.14246, -57.21111, -57.27833, -57.3448, -57.41041, 
        -57.47524, -57.53962, -57.60362, -57.66735, -57.73093, -57.79497, 
        -57.86026, -57.92731, -57.99604, -58.0666, -58.13811, -58.21017, 
        -58.28216, -58.35237, -58.42282, -58.49212, -58.56072, -58.62919, 
        -58.69836, -58.76878, -58.84053, -58.91339, -58.9868, -59.06018, 
        -59.13308, -59.20483, -59.27491, -59.34336, -59.40983, -59.47486, 
        -59.53824, -59.60007, -59.65971, -59.7191, -59.77812, -59.83772, 
        -59.8984, -59.9613, -60.0269, -60.09489, -60.16522, -60.23722, 
        -60.31044, -60.38357, -60.45559, -60.52522, -60.59181, -60.65525, 
        -60.71697, -60.77827, -60.84021, -60.90375, -60.96871, -61.03662, 
        -61.1055, -61.17424, -61.24183, -61.30769, -61.37082, -61.43135, 
        -61.48833, -61.54181, -61.59283, -61.64252, -61.69194, -61.742, 
        -61.79334, -61.84608, -61.90016, -61.95544, -62.0116, -62.06815, 
        -62.12451, -62.17947, -62.23466, -62.28886, -62.3423, -62.39464, 
        -62.44576, -62.49575, -62.5443, -62.59194, -62.63912, -62.6863, 
        -62.73305, -62.77913, -62.82426, -62.86803, -62.9103, -62.95078, 
        -62.98906, -63.02502, -63.05843, -63.08927, -63.11752, -63.14379, 
        -63.168, -63.18941, -63.21041, -63.23139, -63.25269, -63.27517, 
        -63.29892, -63.32399, -63.35, -63.37685, -63.40456, -63.43308, 
        -63.46182, -63.49019, -63.51716, -63.54177, -63.56345, -63.58144, 
        -63.5961, -63.60717, -63.61481, -63.61959, -63.62127, -63.62006, 
        -63.61599, -63.60905, -63.59961, -63.5868, -63.5728, -63.55708, 
        -63.53997, -63.52155, -63.502, -63.48093, -63.45834, -63.43417, 
        -63.40845, -63.38127, -63.3527, -63.32304, -63.2925, -63.26121, 
        -63.22906, -63.19598, -63.16184, -63.12659, -63.09006, -63.05204, 
        -63.01323, -62.9733, -62.93221, -62.89022, -62.84682, -62.80209, 
        -62.75607, -62.70889, -62.65982, -62.61082, -62.5612, -62.51074, 
        -62.45895, -62.40637, -62.35302, -62.29958, -62.24582, -62.19107, 
        -62.13517, -62.07785, -62.01845, -61.95695, -61.89343, -61.8279, 
        -61.76072, -61.69168, -61.62074, -61.54781, -61.47287, -61.39594, 
        -61.31723, -61.23721, -61.15613, -61.0743, -60.99176, -60.90856, 
        -60.82468, -60.74015, -60.65494, -60.56908, -60.4826, -60.39563, 
        -60.30822, -60.22083, -60.13222, -60.04462, -59.95668, -59.86869, 
        -59.78091, -59.69395, -59.60861, -59.52448, -59.44143, -59.35926, 
        -59.2781, -59.19778, -59.11862, -59.04057, -58.96372, -58.88792, 
        -58.81332, -58.74025, -58.66905, -58.60015, -58.53337, -58.46891, 
        -58.40668, -58.34661, -58.2887, -58.23289, -58.17896, -58.12728, 
        -58.07768, -58.0307, -57.98623, -57.94362, -57.90247, -57.86245, 
        -57.82375, -57.78635, -57.75045, -57.71552, -57.6818, -57.64899, 
        -57.61664,
  -47.67503, -47.56512, -47.48244, -47.43017, -47.40834, -47.41472, 
        -47.44534, -47.49542, -47.56216, -47.64368, -47.74052, -47.85469, 
        -47.98905, -48.14869, -48.33575, -48.55684, -48.81163, -49.09626, 
        -49.40592, -49.73278, -50.06757, -50.40091, -50.72636, -51.03969, 
        -51.339, -51.62442, -51.89773, -52.16073, -52.41467, -52.65947, 
        -52.89707, -53.12637, -53.34663, -53.55712, -53.75726, -53.94693, 
        -54.12603, -54.2957, -54.45641, -54.60956, -54.75636, -54.89841, 
        -55.03658, -55.17174, -55.30432, -55.4334, -55.56073, -55.68475, 
        -55.80482, -55.92035, -56.03099, -56.13689, -56.23845, -56.33532, 
        -56.42807, -56.5173, -56.60361, -56.68795, -56.77118, -56.85351, 
        -56.93475, -57.01385, -57.09262, -57.16994, -57.24548, -57.31907, 
        -57.39066, -57.46063, -57.52922, -57.59639, -57.66245, -57.72791, 
        -57.79271, -57.85722, -57.92165, -57.98579, -58.0504, -58.11559, 
        -58.18246, -58.2502, -58.32066, -58.39317, -58.46676, -58.54092, 
        -58.61481, -58.68799, -58.76039, -58.83189, -58.90258, -58.97321, 
        -59.04433, -59.11684, -59.19069, -59.2656, -59.34108, -59.41655, 
        -59.49175, -59.56477, -59.6375, -59.70841, -59.7776, -59.84524, 
        -59.91125, -59.97574, -60.03868, -60.10012, -60.16098, -60.22187, 
        -60.28368, -60.34719, -60.41293, -60.48108, -60.55112, -60.62257, 
        -60.6945, -60.76595, -60.83516, -60.90277, -60.96724, -61.029, 
        -61.08951, -61.14982, -61.21117, -61.27502, -61.34138, -61.41011, 
        -61.48042, -61.55105, -61.62086, -61.6891, -61.75484, -61.81756, 
        -61.87687, -61.93264, -61.98529, -62.03614, -62.08604, -62.13549, 
        -62.18702, -62.23973, -62.29385, -62.34925, -62.40548, -62.46194, 
        -62.51807, -62.57347, -62.62789, -62.68143, -62.73411, -62.78596, 
        -62.83666, -62.88584, -62.93343, -62.9798, -63.02535, -63.07049, 
        -63.11485, -63.15851, -63.20097, -63.24242, -63.28149, -63.31972, 
        -63.35596, -63.38961, -63.42059, -63.44872, -63.47401, -63.49673, 
        -63.51703, -63.53485, -63.55114, -63.56709, -63.58295, -63.60027, 
        -63.61906, -63.63958, -63.66156, -63.68491, -63.70989, -63.73596, 
        -63.76227, -63.78831, -63.81333, -63.83638, -63.85666, -63.87234, 
        -63.88546, -63.89497, -63.90108, -63.9036, -63.90295, -63.89907, 
        -63.89238, -63.88303, -63.8713, -63.85732, -63.84118, -63.82328, 
        -63.804, -63.78349, -63.76175, -63.73842, -63.71365, -63.68757, 
        -63.66007, -63.63135, -63.60142, -63.57057, -63.53896, -63.50694, 
        -63.47445, -63.44127, -63.40737, -63.37157, -63.33546, -63.29799, 
        -63.2593, -63.21947, -63.17846, -63.13625, -63.09262, -63.0477, 
        -63.00136, -62.95393, -62.90565, -62.85661, -62.80696, -62.7562, 
        -62.70448, -62.65189, -62.59894, -62.54534, -62.49115, -62.43606, 
        -62.37963, -62.32169, -62.26162, -62.19978, -62.13599, -62.07055, 
        -62.00374, -61.93528, -61.86521, -61.79332, -61.71953, -61.64384, 
        -61.56551, -61.48698, -61.40774, -61.32759, -61.24658, -61.16455, 
        -61.08168, -60.99765, -60.91277, -60.8272, -60.74096, -60.65416, 
        -60.56703, -60.47989, -60.39283, -60.30587, -60.21894, -60.13184, 
        -60.04488, -59.95855, -59.87332, -59.78935, -59.7064, -59.62455, 
        -59.54365, -59.46385, -59.38552, -59.30869, -59.23275, -59.1579, 
        -59.08384, -59.01101, -58.93979, -58.87054, -58.80352, -58.73869, 
        -58.67634, -58.61634, -58.55835, -58.50216, -58.44761, -58.39506, 
        -58.34368, -58.29572, -58.25041, -58.20721, -58.16527, -58.12437, 
        -58.08464, -58.04635, -58.00942, -57.97396, -57.93966, -57.90616, 
        -57.87337,
  -47.77569, -47.67884, -47.60964, -47.57043, -47.56054, -47.57685, 
        -47.615, -47.67039, -47.73879, -47.82096, -47.91655, -48.02799, 
        -48.15864, -48.31265, -48.4942, -48.70652, -48.95074, -49.22434, 
        -49.52365, -49.84058, -50.16702, -50.49438, -50.81577, -51.12655, 
        -51.42694, -51.71611, -51.99547, -52.26689, -52.53118, -52.78882, 
        -53.03885, -53.28038, -53.51215, -53.73306, -53.94216, -54.13932, 
        -54.32482, -54.49963, -54.66467, -54.82064, -54.97137, -55.11744, 
        -55.26024, -55.40043, -55.53875, -55.67519, -55.80926, -55.94045, 
        -56.06826, -56.1915, -56.30988, -56.42307, -56.53143, -56.63433, 
        -56.73229, -56.82458, -56.91429, -57.00116, -57.08638, -57.17023, 
        -57.25282, -57.33402, -57.41354, -57.49138, -57.56744, -57.64133, 
        -57.71302, -57.78274, -57.8509, -57.91781, -57.98361, -58.04891, 
        -58.11284, -58.17755, -58.24232, -58.30716, -58.37266, -58.43916, 
        -58.5071, -58.57714, -58.64945, -58.7236, -58.79882, -58.87455, 
        -58.95007, -59.02515, -59.09952, -59.17303, -59.24577, -59.31856, 
        -59.39075, -59.46526, -59.54093, -59.61786, -59.6954, -59.77304, 
        -59.85038, -59.9267, -60.00183, -60.07532, -60.14722, -60.21746, 
        -60.28599, -60.35277, -60.41776, -60.48133, -60.54399, -60.60614, 
        -60.66879, -60.73198, -60.79812, -60.86646, -60.93647, -61.00735, 
        -61.07827, -61.14861, -61.21724, -61.28313, -61.34626, -61.40735, 
        -61.46695, -61.52658, -61.58757, -61.65115, -61.71754, -61.78667, 
        -61.85771, -61.92948, -62.00067, -62.07051, -62.13716, -62.20197, 
        -62.26325, -62.32084, -62.37539, -62.42746, -62.47815, -62.52876, 
        -62.57992, -62.63242, -62.68633, -62.74162, -62.79773, -62.85383, 
        -62.90922, -62.96356, -63.01683, -63.06937, -63.12132, -63.17252, 
        -63.22253, -63.271, -63.31661, -63.36166, -63.40523, -63.44791, 
        -63.48947, -63.53023, -63.56993, -63.60867, -63.64624, -63.6823, 
        -63.71643, -63.74805, -63.77694, -63.80287, -63.82581, -63.84554, 
        -63.86185, -63.87576, -63.88822, -63.8992, -63.91034, -63.92282, 
        -63.93656, -63.95211, -63.96834, -63.98826, -64.00968, -64.03232, 
        -64.05541, -64.07851, -64.10074, -64.12118, -64.1389, -64.1535, 
        -64.1647, -64.17219, -64.17606, -64.17622, -64.17323, -64.16696, 
        -64.15781, -64.14622, -64.13261, -64.1168, -64.09887, -64.07921, 
        -64.05799, -64.03534, -64.01124, -63.98569, -63.9589, -63.92991, 
        -63.90078, -63.87057, -63.83942, -63.80744, -63.77505, -63.74231, 
        -63.70928, -63.67606, -63.64236, -63.60795, -63.57233, -63.53524, 
        -63.49665, -63.45689, -63.41593, -63.37383, -63.33028, -63.28531, 
        -63.23888, -63.19129, -63.14291, -63.09382, -63.0441, -62.99329, 
        -62.94158, -62.88914, -62.83611, -62.7827, -62.72833, -62.67254, 
        -62.61457, -62.55614, -62.49546, -62.43281, -62.36844, -62.30264, 
        -62.23564, -62.16728, -62.09754, -62.02618, -61.95309, -61.87829, 
        -61.80196, -61.7247, -61.64695, -61.56856, -61.48925, -61.40866, 
        -61.32686, -61.24381, -61.15969, -61.0747, -60.989, -60.90271, 
        -60.81604, -60.72937, -60.6428, -60.55643, -60.47032, -60.38433, 
        -60.29852, -60.21313, -60.12848, -60.04479, -59.96202, -59.88021, 
        -59.7995, -59.72031, -59.64185, -59.56589, -59.49096, -59.41684, 
        -59.34351, -59.27106, -59.20005, -59.13076, -59.06374, -58.99916, 
        -58.93728, -58.87765, -58.81989, -58.7635, -58.7081, -58.65474, 
        -58.60345, -58.55478, -58.50865, -58.46456, -58.4219, -58.38031, 
        -58.33975, -58.30061, -58.26287, -58.22655, -58.19147, -58.15725, 
        -58.12368,
  -47.88783, -47.80572, -47.75104, -47.72445, -47.72651, -47.7525, 
        -47.79782, -47.85819, -47.93043, -48.0137, -48.10906, -48.21912, 
        -48.34752, -48.49792, -48.67429, -48.87903, -49.11428, -49.37757, 
        -49.66412, -49.96988, -50.28609, -50.60508, -50.92052, -51.22929, 
        -51.52934, -51.82114, -52.10572, -52.38468, -52.65849, -52.92685, 
        -53.18852, -53.44151, -53.6842, -53.91403, -54.13172, -54.33631, 
        -54.52814, -54.70816, -54.87766, -55.03842, -55.19258, -55.34211, 
        -55.48882, -55.63352, -55.7771, -55.91937, -56.05999, -56.19849, 
        -56.33372, -56.46404, -56.59031, -56.7114, -56.82698, -56.93628, 
        -57.0396, -57.1372, -57.23036, -57.31989, -57.40693, -57.49207, 
        -57.57568, -57.65767, -57.73779, -57.81601, -57.89224, -57.96641, 
        -58.03723, -58.10674, -58.17457, -58.2412, -58.30721, -58.37239, 
        -58.43747, -58.50253, -58.56769, -58.63308, -58.6992, -58.76643, 
        -58.83537, -58.90642, -58.97976, -59.05518, -59.13182, -59.20903, 
        -59.28498, -59.36163, -59.43751, -59.51274, -59.58758, -59.66232, 
        -59.73751, -59.81379, -59.89141, -59.97023, -60.0498, -60.1295, 
        -60.2089, -60.28756, -60.3651, -60.44107, -60.51559, -60.58827, 
        -60.65828, -60.72736, -60.79419, -60.85962, -60.92379, -60.98742, 
        -61.05117, -61.11609, -61.18272, -61.25114, -61.32117, -61.39187, 
        -61.46233, -61.53188, -61.59963, -61.66486, -61.72737, -61.7879, 
        -61.84713, -61.90645, -61.96632, -62.02951, -62.09552, -62.16441, 
        -62.23526, -62.3072, -62.37894, -62.44947, -62.51804, -62.58411, 
        -62.64698, -62.70633, -62.76214, -62.81523, -62.86648, -62.91718, 
        -62.96807, -63.02026, -63.07375, -63.1286, -63.18433, -63.23864, 
        -63.29294, -63.346, -63.39801, -63.44938, -63.50039, -63.55071, 
        -63.59996, -63.64763, -63.69329, -63.73684, -63.77853, -63.81871, 
        -63.8575, -63.89526, -63.93213, -63.96806, -64.00296, -64.03649, 
        -64.06826, -64.09786, -64.12473, -64.14854, -64.1691, -64.18506, 
        -64.19866, -64.20924, -64.21743, -64.22441, -64.23119, -64.2389, 
        -64.24752, -64.25803, -64.27113, -64.28642, -64.304, -64.32294, 
        -64.34168, -64.36098, -64.37952, -64.39651, -64.41109, -64.42288, 
        -64.43139, -64.43636, -64.43767, -64.43555, -64.43007, -64.42161, 
        -64.40923, -64.39578, -64.38036, -64.36288, -64.34332, -64.32214, 
        -64.29903, -64.2744, -64.24839, -64.22101, -64.19239, -64.16256, 
        -64.13201, -64.10034, -64.06812, -64.03514, -64.00183, -63.96833, 
        -63.93488, -63.90131, -63.86742, -63.83292, -63.79738, -63.7605, 
        -63.72205, -63.68246, -63.64178, -63.59991, -63.55665, -63.5119, 
        -63.46458, -63.41696, -63.36863, -63.31944, -63.26939, -63.21861, 
        -63.16695, -63.11469, -63.06171, -63.00824, -62.95402, -62.89802, 
        -62.84068, -62.78145, -62.72023, -62.65718, -62.59235, -62.52611, 
        -62.45853, -62.38988, -62.31995, -62.24846, -62.17545, -62.1011, 
        -62.02569, -61.94942, -61.87288, -61.79605, -61.71823, -61.63934, 
        -61.55884, -61.47692, -61.39381, -61.30978, -61.22485, -61.13836, 
        -61.0525, -60.96667, -60.88081, -60.79525, -60.71009, -60.62518, 
        -60.54044, -60.4558, -60.37192, -60.28858, -60.20596, -60.12429, 
        -60.04387, -59.96511, -59.88823, -59.81291, -59.73881, -59.66543, 
        -59.5927, -59.52069, -59.45013, -59.38128, -59.31472, -59.25061, 
        -59.18905, -59.12983, -59.07232, -59.01588, -58.96046, -58.90649, 
        -58.85463, -58.80535, -58.75853, -58.71391, -58.67063, -58.62842, 
        -58.58723, -58.54734, -58.50875, -58.47143, -58.43522, -58.40019, 
        -58.36582,
  -48.01151, -47.9454, -47.90625, -47.89424, -47.90722, -47.9423, 
        -47.99409, -48.05869, -48.1338, -48.21901, -48.31538, -48.42543, 
        -48.55328, -48.70125, -48.87437, -49.07403, -49.30145, -49.5552, 
        -49.83157, -50.12553, -50.43052, -50.74007, -51.04836, -51.35292, 
        -51.65145, -51.94407, -52.23239, -52.51739, -52.79827, -53.07611, 
        -53.34791, -53.61107, -53.86336, -54.10312, -54.329, -54.54071, 
        -54.7387, -54.92392, -55.09789, -55.26246, -55.4198, -55.57241, 
        -55.72243, -55.87016, -56.01828, -56.16592, -56.31269, -56.45799, 
        -56.60051, -56.73962, -56.87397, -57.00305, -57.12552, -57.2412, 
        -57.34978, -57.45195, -57.54839, -57.64048, -57.72941, -57.81582, 
        -57.89937, -57.98207, -58.06281, -58.14143, -58.21767, -58.29161, 
        -58.36364, -58.43328, -58.50113, -58.56775, -58.63381, -58.69949, 
        -58.76462, -58.82997, -58.89566, -58.96162, -59.02837, -59.09529, 
        -59.16483, -59.23643, -59.31031, -59.38658, -59.46412, -59.54223, 
        -59.62045, -59.69828, -59.77534, -59.85195, -59.92848, -60.00513, 
        -60.08231, -60.16029, -60.23949, -60.32011, -60.40152, -60.48228, 
        -60.56381, -60.64453, -60.72428, -60.80296, -60.87988, -60.95489, 
        -61.02814, -61.09951, -61.16843, -61.23577, -61.3012, -61.36635, 
        -61.43138, -61.49713, -61.56413, -61.63275, -61.70269, -61.77342, 
        -61.84397, -61.91235, -61.97981, -62.04489, -62.10756, -62.16824, 
        -62.22774, -62.28721, -62.34772, -62.41039, -62.47568, -62.54367, 
        -62.61378, -62.68503, -62.75632, -62.82669, -62.89529, -62.96187, 
        -63.02553, -63.08569, -63.1425, -63.19622, -63.24686, -63.29751, 
        -63.34783, -63.39935, -63.45246, -63.50707, -63.56202, -63.61629, 
        -63.66935, -63.72093, -63.77145, -63.82164, -63.87143, -63.92088, 
        -63.96934, -64.01617, -64.06081, -64.10295, -64.14272, -64.18045, 
        -64.21664, -64.25149, -64.28445, -64.3175, -64.34947, -64.38023, 
        -64.40949, -64.43683, -64.46181, -64.48374, -64.50207, -64.51671, 
        -64.52751, -64.53506, -64.54002, -64.54342, -64.5462, -64.54931, 
        -64.55323, -64.55905, -64.56741, -64.57867, -64.5915, -64.60601, 
        -64.6206, -64.63544, -64.64935, -64.66078, -64.6714, -64.67958, 
        -64.68487, -64.68689, -64.68536, -64.68052, -64.67249, -64.6617, 
        -64.64844, -64.63315, -64.61632, -64.59736, -64.57635, -64.55327, 
        -64.52882, -64.50238, -64.47432, -64.4451, -64.41483, -64.38354, 
        -64.35153, -64.31875, -64.28542, -64.25164, -64.21755, -64.18345, 
        -64.14922, -64.11398, -64.07952, -64.04459, -64.00876, -63.97171, 
        -63.9335, -63.89403, -63.85351, -63.81184, -63.76881, -63.72422, 
        -63.67825, -63.63097, -63.58281, -63.5337, -63.48373, -63.43301, 
        -63.38179, -63.33002, -63.27773, -63.22425, -63.16999, -63.11407, 
        -63.05631, -62.99665, -62.93507, -62.8715, -62.80634, -62.7396, 
        -62.67164, -62.60246, -62.53193, -62.45897, -62.38583, -62.31164, 
        -62.23655, -62.161, -62.08532, -62.00951, -61.93314, -61.85569, 
        -61.77671, -61.69617, -61.61425, -61.53125, -61.44762, -61.36321, 
        -61.2784, -61.19341, -61.10818, -61.02341, -60.9392, -60.85531, 
        -60.77161, -60.68814, -60.60481, -60.52197, -60.43941, -60.35796, 
        -60.27755, -60.19906, -60.12263, -60.04794, -59.9743, -59.90124, 
        -59.82891, -59.75744, -59.6873, -59.61913, -59.55313, -59.48967, 
        -59.42868, -59.3698, -59.31149, -59.25529, -59.20007, -59.146, 
        -59.09409, -59.04452, -58.99734, -58.95226, -58.90845, -58.86624, 
        -58.82487, -58.78457, -58.74527, -58.70678, -58.66971, -58.6335, 
        -58.59813,
  -48.15039, -48.10073, -48.07646, -48.07739, -48.10099, -48.14367, 
        -48.2012, -48.26878, -48.34671, -48.43407, -48.53244, -48.64463, 
        -48.77376, -48.92311, -49.09513, -49.29146, -49.51338, -49.75925, 
        -50.02597, -50.30917, -50.60342, -50.9034, -51.20323, -51.50216, 
        -51.79808, -52.09097, -52.38166, -52.67081, -52.95829, -53.24282, 
        -53.52198, -53.79304, -54.05311, -54.30044, -54.53354, -54.75196, 
        -54.95599, -55.14659, -55.32421, -55.49272, -55.65347, -55.8091, 
        -55.96202, -56.11391, -56.26583, -56.41788, -56.56984, -56.72109, 
        -56.87047, -57.01689, -57.15891, -57.29508, -57.42443, -57.54609, 
        -57.65908, -57.76563, -57.86563, -57.9604, -58.05123, -58.13892, 
        -58.22424, -58.30745, -58.38843, -58.46736, -58.54374, -58.6177, 
        -58.68971, -58.75982, -58.82824, -58.89536, -58.96181, -59.02688, 
        -59.09274, -59.15845, -59.22446, -59.29096, -59.35811, -59.42643, 
        -59.49624, -59.5682, -59.64232, -59.71866, -59.7967, -59.87549, 
        -59.95439, -60.03281, -60.1109, -60.18854, -60.26628, -60.34352, 
        -60.42226, -60.50202, -60.58292, -60.66504, -60.74815, -60.83163, 
        -60.91505, -60.99778, -61.0795, -61.16024, -61.23943, -61.31684, 
        -61.39224, -61.4655, -61.53661, -61.60563, -61.67302, -61.73941, 
        -61.80469, -61.87137, -61.93912, -62.00805, -62.07819, -62.14887, 
        -62.21951, -62.28926, -62.35728, -62.42308, -62.48657, -62.54812, 
        -62.60831, -62.66817, -62.72849, -62.79035, -62.85453, -62.92118, 
        -62.98993, -63.05987, -63.12901, -63.19847, -63.2665, -63.33259, 
        -63.39612, -63.45651, -63.51356, -63.5677, -63.61953, -63.67007, 
        -63.72021, -63.77117, -63.82348, -63.87699, -63.93084, -63.98394, 
        -64.03546, -64.08553, -64.13465, -64.18341, -64.23226, -64.28083, 
        -64.32743, -64.37331, -64.41697, -64.45778, -64.49577, -64.53142, 
        -64.56499, -64.59717, -64.6282, -64.65815, -64.68712, -64.71497, 
        -64.7415, -64.76631, -64.78895, -64.8086, -64.82462, -64.83688, 
        -64.84518, -64.85006, -64.85213, -64.85246, -64.85189, -64.85094, 
        -64.84978, -64.8513, -64.85522, -64.86165, -64.87003, -64.87949, 
        -64.88942, -64.89917, -64.90823, -64.91613, -64.92233, -64.92653, 
        -64.92805, -64.92653, -64.92164, -64.9136, -64.90265, -64.88915, 
        -64.8738, -64.85679, -64.8381, -64.81778, -64.79552, -64.77119, 
        -64.745, -64.7169, -64.68644, -64.65578, -64.62408, -64.59164, 
        -64.55836, -64.52455, -64.49018, -64.4556, -64.42081, -64.38576, 
        -64.35068, -64.31549, -64.28012, -64.24432, -64.20798, -64.17081, 
        -64.13261, -64.09335, -64.05302, -64.01163, -63.96888, -63.92466, 
        -63.87899, -63.83206, -63.78421, -63.73529, -63.6855, -63.63514, 
        -63.58414, -63.53282, -63.48071, -63.42668, -63.37215, -63.31605, 
        -63.25818, -63.19852, -63.13712, -63.07385, -63.0087, -62.94191, 
        -62.87367, -62.80394, -62.73288, -62.66053, -62.58695, -62.5124, 
        -62.43726, -62.36181, -62.28653, -62.21133, -62.13591, -62.05971, 
        -61.98207, -61.90287, -61.82221, -61.74047, -61.65792, -61.57465, 
        -61.49096, -61.40691, -61.3229, -61.23925, -61.15612, -61.07352, 
        -60.99104, -60.90855, -60.82584, -60.74325, -60.65988, -60.57821, 
        -60.49781, -60.41945, -60.34322, -60.26867, -60.19539, -60.12283, 
        -60.05091, -59.97984, -59.91041, -59.84273, -59.77716, -59.71402, 
        -59.65319, -59.59434, -59.5371, -59.4809, -59.42585, -59.37203, 
        -59.32034, -59.27084, -59.22373, -59.17847, -59.13481, -59.09255, 
        -59.05123, -59.0108, -58.97118, -58.93226, -58.89437, -58.85743, 
        -58.82141,
  -48.30708, -48.27364, -48.26311, -48.27587, -48.30849, -48.35709, 
        -48.41893, -48.49055, -48.57081, -48.66056, -48.76168, -48.8767, 
        -49.00875, -49.16038, -49.33369, -49.52939, -49.74829, -49.98774, 
        -50.24685, -50.5208, -50.8053, -51.09609, -51.3896, -51.68279, 
        -51.97549, -52.26686, -52.55818, -52.8492, -53.13967, -53.42821, 
        -53.71211, -53.98841, -54.25322, -54.50648, -54.74586, -54.97026, 
        -55.1799, -55.37587, -55.55933, -55.73215, -55.89645, -56.05514, 
        -56.21066, -56.36528, -56.52014, -56.67574, -56.83201, -56.98822, 
        -57.14249, -57.29512, -57.4436, -57.58633, -57.72159, -57.84862, 
        -57.96709, -58.07767, -58.18121, -58.27864, -58.37155, -58.46071, 
        -58.54702, -58.63073, -58.71212, -58.79133, -58.86794, -58.9413, 
        -59.01342, -59.0841, -59.15322, -59.22145, -59.28876, -59.35564, 
        -59.42215, -59.48825, -59.55457, -59.62136, -59.68882, -59.75739, 
        -59.82729, -59.89917, -59.97329, -60.04951, -60.12641, -60.20543, 
        -60.28466, -60.36358, -60.44201, -60.52034, -60.59905, -60.67847, 
        -60.75878, -60.84008, -60.92252, -61.00611, -61.09051, -61.17548, 
        -61.26034, -61.3446, -61.42812, -61.51069, -61.59178, -61.67012, 
        -61.74751, -61.82304, -61.89621, -61.96736, -62.03662, -62.10479, 
        -62.1725, -62.24023, -62.30848, -62.37754, -62.44769, -62.51845, 
        -62.58932, -62.65951, -62.72854, -62.79562, -62.8606, -62.92368, 
        -62.98395, -63.04424, -63.10421, -63.16512, -63.22776, -63.29269, 
        -63.35959, -63.42779, -63.49645, -63.56435, -63.6314, -63.69651, 
        -63.75911, -63.8189, -63.87583, -63.93002, -63.98187, -64.03234, 
        -64.08216, -64.13254, -64.18388, -64.23614, -64.28764, -64.33921, 
        -64.38914, -64.43772, -64.48554, -64.53306, -64.58076, -64.62828, 
        -64.67508, -64.72016, -64.76279, -64.80238, -64.83884, -64.87246, 
        -64.90381, -64.93342, -64.96162, -64.98853, -65.01436, -65.0392, 
        -65.06274, -65.08487, -65.10486, -65.12081, -65.13423, -65.14388, 
        -65.14967, -65.15176, -65.15144, -65.14912, -65.14574, -65.1418, 
        -65.13804, -65.13564, -65.13529, -65.13706, -65.14068, -65.14525, 
        -65.15002, -65.15453, -65.15837, -65.16128, -65.16291, -65.16297, 
        -65.16035, -65.15485, -65.14628, -65.13472, -65.11951, -65.10333, 
        -65.0855, -65.06641, -65.04586, -65.02386, -65.00014, -64.97427, 
        -64.94658, -64.917, -64.88615, -64.85419, -64.82143, -64.78777, 
        -64.75342, -64.7187, -64.68357, -64.64825, -64.61273, -64.57686, 
        -64.5408, -64.50445, -64.46795, -64.43123, -64.39414, -64.35664, 
        -64.31839, -64.27919, -64.23892, -64.19652, -64.15406, -64.1099, 
        -64.06496, -64.01857, -63.97135, -63.92282, -63.8734, -63.82313, 
        -63.77254, -63.72135, -63.66951, -63.61636, -63.56156, -63.50544, 
        -63.44766, -63.38855, -63.32772, -63.26533, -63.20086, -63.1346, 
        -63.06645, -62.99638, -62.92483, -62.85173, -62.77735, -62.70235, 
        -62.62666, -62.55079, -62.47538, -62.40025, -62.3253, -62.24976, 
        -62.17339, -62.09555, -62.01518, -61.93478, -61.85334, -61.77121, 
        -61.68851, -61.60557, -61.52273, -61.44039, -61.35863, -61.27729, 
        -61.19575, -61.11414, -61.0321, -60.94984, -60.86746, -60.78558, 
        -60.70519, -60.62685, -60.55057, -60.47616, -60.40292, -60.33039, 
        -60.25877, -60.18821, -60.11916, -60.05212, -59.98721, -59.92419, 
        -59.86293, -59.8035, -59.74572, -59.68947, -59.63477, -59.58167, 
        -59.53054, -59.48163, -59.43469, -59.38988, -59.34673, -59.30484, 
        -59.2639, -59.22391, -59.18465, -59.14581, -59.10765, -59.06931, 
        -59.03315,
  -48.48259, -48.46478, -48.46812, -48.491, -48.5309, -48.58439, 
        -48.64891, -48.7229, -48.80534, -48.89769, -49.00205, -49.11999, 
        -49.25614, -49.41191, -49.58811, -49.78508, -50.00328, -50.24064, 
        -50.49453, -50.76157, -51.03826, -51.32151, -51.60817, -51.89616, 
        -52.1847, -52.47371, -52.76247, -53.05298, -53.34369, -53.63298, 
        -53.91845, -54.19731, -54.46671, -54.72435, -54.96889, -55.19886, 
        -55.41439, -55.61593, -55.80454, -55.98188, -56.14969, -56.31125, 
        -56.46812, -56.62474, -56.78165, -56.93956, -57.09889, -57.2589, 
        -57.41849, -57.57607, -57.72965, -57.87751, -58.01786, -58.14933, 
        -58.27187, -58.38598, -58.49252, -58.59257, -58.68736, -58.77703, 
        -58.86435, -58.94879, -59.03073, -59.11021, -59.18732, -59.26214, 
        -59.33504, -59.40635, -59.47641, -59.54558, -59.61407, -59.68202, 
        -59.74933, -59.81629, -59.88301, -59.95026, -60.01703, -60.08576, 
        -60.15587, -60.22742, -60.30107, -60.37696, -60.45454, -60.53337, 
        -60.61258, -60.6914, -60.76994, -60.84872, -60.92792, -61.00803, 
        -61.08932, -61.17176, -61.25539, -61.3401, -61.42448, -61.51053, 
        -61.59692, -61.68279, -61.76784, -61.8518, -61.93438, -62.01537, 
        -62.09461, -62.17207, -62.24739, -62.32079, -62.39223, -62.46253, 
        -62.53181, -62.60077, -62.66984, -62.73916, -62.80927, -62.87901, 
        -62.95005, -63.02089, -63.09081, -63.15924, -63.22577, -63.29021, 
        -63.3527, -63.41349, -63.4733, -63.53332, -63.59441, -63.65736, 
        -63.72203, -63.78812, -63.85468, -63.921, -63.98622, -64.04948, 
        -64.11083, -64.16967, -64.22514, -64.27915, -64.33118, -64.38165, 
        -64.43143, -64.48128, -64.53145, -64.58237, -64.63279, -64.68278, 
        -64.73123, -64.77824, -64.82475, -64.87096, -64.91762, -64.96419, 
        -65.01002, -65.05406, -65.09556, -65.13387, -65.16899, -65.2011, 
        -65.22964, -65.257, -65.28258, -65.30685, -65.32965, -65.35143, 
        -65.37194, -65.39105, -65.40802, -65.42214, -65.43282, -65.43964, 
        -65.44274, -65.4427, -65.43999, -65.43517, -65.42934, -65.42249, 
        -65.41557, -65.40937, -65.40482, -65.40205, -65.40072, -65.40049, 
        -65.4003, -65.39886, -65.39782, -65.39581, -65.39275, -65.38804, 
        -65.38123, -65.3714, -65.35859, -65.34321, -65.32556, -65.30611, 
        -65.28535, -65.26369, -65.24097, -65.2169, -65.19132, -65.16398, 
        -65.13477, -65.10396, -65.07201, -65.03903, -65.0052, -64.97074, 
        -64.93558, -64.90014, -64.8644, -64.8283, -64.79108, -64.75443, 
        -64.7173, -64.67992, -64.6424, -64.60481, -64.56709, -64.52925, 
        -64.49085, -64.45164, -64.41131, -64.36983, -64.32722, -64.28357, 
        -64.23895, -64.19328, -64.14635, -64.0982, -64.04873, -63.99863, 
        -63.94797, -63.89683, -63.8453, -63.79232, -63.73775, -63.68187, 
        -63.62484, -63.56659, -63.50682, -63.44539, -63.38184, -63.31589, 
        -63.2469, -63.17664, -63.10442, -63.03068, -62.95574, -62.8798, 
        -62.80335, -62.72698, -62.65107, -62.57578, -62.50097, -62.42623, 
        -62.35052, -62.27358, -62.1953, -62.11572, -62.03507, -61.95369, 
        -61.87192, -61.79002, -61.70855, -61.62758, -61.54721, -61.46709, 
        -61.38685, -61.30623, -61.22462, -61.14246, -61.06009, -60.97824, 
        -60.89774, -60.81918, -60.74254, -60.6678, -60.5944, -60.52195, 
        -60.45057, -60.38037, -60.31206, -60.24558, -60.18077, -60.11669, 
        -60.05478, -59.99458, -59.93629, -59.87958, -59.82485, -59.77221, 
        -59.72171, -59.67342, -59.62732, -59.58333, -59.54106, -59.5001, 
        -59.46017, -59.42106, -59.38234, -59.34384, -59.30613, -59.26917, 
        -59.23341,
  -48.67912, -48.67568, -48.69016, -48.72136, -48.76666, -48.82331, 
        -48.88882, -48.96412, -49.0484, -49.14339, -49.25132, -49.37482, 
        -49.5161, -49.6769, -49.85757, -50.05791, -50.27729, -50.51385, 
        -50.76481, -51.02747, -51.29871, -51.57471, -51.85566, -52.13861, 
        -52.42272, -52.70811, -52.99487, -53.28275, -53.57099, -53.85839, 
        -54.14275, -54.42183, -54.69296, -54.95361, -55.20221, -55.43765, 
        -55.65786, -55.86499, -56.0588, -56.24076, -56.41256, -56.57684, 
        -56.73664, -56.89469, -57.0528, -57.21219, -57.37326, -57.53556, 
        -57.69803, -57.85894, -58.0162, -58.16759, -58.31153, -58.44542, 
        -58.57099, -58.68786, -58.79694, -58.89916, -58.99606, -59.08816, 
        -59.17646, -59.26169, -59.34412, -59.42421, -59.50188, -59.57748, 
        -59.65136, -59.72354, -59.79465, -59.86486, -59.93349, -60.00258, 
        -60.07104, -60.13891, -60.20656, -60.27427, -60.3424, -60.41144, 
        -60.48158, -60.55302, -60.62634, -60.70156, -60.77866, -60.85693, 
        -60.93566, -61.01448, -61.0929, -61.17049, -61.24971, -61.33004, 
        -61.41179, -61.49487, -61.57919, -61.66468, -61.75115, -61.83836, 
        -61.92569, -62.013, -62.09937, -62.18465, -62.26849, -62.35078, 
        -62.4316, -62.51093, -62.58853, -62.6641, -62.73699, -62.80944, 
        -62.88057, -62.95109, -63.02101, -63.09098, -63.16132, -63.23205, 
        -63.30308, -63.37411, -63.4446, -63.51398, -63.58168, -63.64739, 
        -63.71078, -63.77206, -63.83179, -63.89101, -63.95066, -64.01164, 
        -64.07301, -64.13647, -64.20054, -64.26438, -64.32755, -64.38911, 
        -64.44874, -64.50647, -64.56221, -64.61615, -64.66828, -64.71884, 
        -64.76839, -64.81753, -64.86698, -64.91624, -64.96506, -65.01297, 
        -65.05971, -65.10555, -65.15072, -65.19566, -65.2402, -65.28559, 
        -65.33018, -65.37312, -65.4133, -65.45042, -65.48438, -65.51514, 
        -65.54329, -65.56889, -65.59251, -65.61427, -65.63441, -65.65323, 
        -65.67065, -65.68661, -65.70062, -65.71161, -65.71924, -65.72314, 
        -65.72368, -65.72095, -65.71507, -65.70818, -65.69952, -65.69028, 
        -65.68029, -65.67045, -65.66182, -65.65462, -65.64848, -65.64352, 
        -65.63867, -65.63363, -65.62778, -65.6211, -65.61342, -65.60391, 
        -65.5922, -65.57769, -65.56041, -65.54086, -65.51936, -65.49641, 
        -65.47253, -65.44779, -65.42234, -65.39584, -65.3681, -65.3379, 
        -65.30722, -65.27528, -65.24224, -65.20842, -65.17384, -65.13861, 
        -65.10291, -65.06693, -65.03071, -64.99424, -64.95741, -64.92027, 
        -64.88255, -64.84428, -64.80595, -64.76768, -64.72956, -64.69124, 
        -64.65257, -64.61301, -64.57245, -64.53086, -64.48812, -64.44463, 
        -64.40022, -64.35474, -64.30817, -64.26015, -64.20983, -64.15987, 
        -64.10928, -64.05849, -64.00706, -63.9545, -63.90062, -63.84517, 
        -63.78898, -63.73154, -63.6727, -63.61198, -63.54903, -63.48336, 
        -63.41525, -63.34489, -63.27233, -63.1981, -63.12246, -63.04586, 
        -62.96884, -62.89177, -62.81533, -62.73981, -62.66511, -62.59062, 
        -62.51569, -62.43958, -62.36212, -62.28316, -62.20304, -62.12197, 
        -62.04073, -61.95966, -61.87897, -61.7992, -61.72003, -61.64109, 
        -61.5618, -61.48088, -61.39992, -61.31783, -61.23542, -61.1535, 
        -61.07274, -60.99374, -60.9166, -60.84127, -60.76744, -60.69491, 
        -60.62365, -60.55399, -60.48621, -60.42023, -60.35545, -60.29201, 
        -60.22968, -60.1686, -60.10952, -60.0526, -59.99794, -59.94573, 
        -59.89605, -59.84857, -59.8034, -59.76046, -59.7193, -59.67966, 
        -59.64106, -59.60304, -59.56537, -59.52783, -59.4909, -59.45471, 
        -59.41964,
  -48.89365, -48.90207, -48.92626, -48.96365, -49.01254, -49.07115, 
        -49.13853, -49.21476, -49.30064, -49.39834, -49.51027, -49.6389, 
        -49.7865, -49.95327, -50.13953, -50.34412, -50.56477, -50.80205, 
        -51.0518, -51.31171, -51.57907, -51.85162, -52.12785, -52.40604, 
        -52.68552, -52.96652, -53.24902, -53.53289, -53.8168, -54.10046, 
        -54.38214, -54.65872, -54.93, -55.1928, -55.44487, -55.68499, 
        -55.91181, -56.12466, -56.3238, -56.51036, -56.68594, -56.853, 
        -57.01452, -57.17346, -57.3322, -57.49213, -57.65394, -57.81626, 
        -57.98007, -58.14272, -58.30177, -58.4551, -58.60089, -58.73786, 
        -58.86542, -58.98428, -59.09529, -59.19946, -59.29784, -59.39135, 
        -59.48077, -59.56686, -59.64996, -59.72957, -59.80801, -59.88432, 
        -59.95914, -60.03256, -60.10484, -60.17619, -60.24697, -60.31731, 
        -60.387, -60.45601, -60.52451, -60.5929, -60.66168, -60.73096, 
        -60.80123, -60.8727, -60.94567, -61.0195, -61.09595, -61.17365, 
        -61.2519, -61.33015, -61.40836, -61.48663, -61.56567, -61.64589, 
        -61.72745, -61.81053, -61.89524, -61.98121, -62.06836, -62.1563, 
        -62.2448, -62.33314, -62.42073, -62.50625, -62.59131, -62.67509, 
        -62.75725, -62.83836, -62.91801, -62.99592, -63.07235, -63.14697, 
        -63.22004, -63.29229, -63.36349, -63.43417, -63.50476, -63.57536, 
        -63.6461, -63.7169, -63.78741, -63.85715, -63.92559, -63.99084, 
        -64.05486, -64.11646, -64.17607, -64.2347, -64.29315, -64.35232, 
        -64.41232, -64.47303, -64.53416, -64.59545, -64.65612, -64.71565, 
        -64.77384, -64.83046, -64.88552, -64.93904, -64.99102, -65.04163, 
        -65.09096, -65.13933, -65.18662, -65.23416, -65.28111, -65.32742, 
        -65.37283, -65.4174, -65.46152, -65.50549, -65.5496, -65.59348, 
        -65.6366, -65.67815, -65.71729, -65.75338, -65.78634, -65.81624, 
        -65.84327, -65.86771, -65.88962, -65.90922, -65.92699, -65.94305, 
        -65.9567, -65.96964, -65.98042, -65.98824, -65.99286, -65.99402, 
        -65.99169, -65.98633, -65.97863, -65.96922, -65.95826, -65.94563, 
        -65.93267, -65.9194, -65.90678, -65.89536, -65.88509, -65.87576, 
        -65.86673, -65.85733, -65.84728, -65.83611, -65.82355, -65.80903, 
        -65.79222, -65.77184, -65.74998, -65.72587, -65.7002, -65.67344, 
        -65.64609, -65.61813, -65.58952, -65.56043, -65.53029, -65.49921, 
        -65.46668, -65.43334, -65.39887, -65.36401, -65.32858, -65.29274, 
        -65.25652, -65.22024, -65.18398, -65.14751, -65.1106, -65.07323, 
        -65.03526, -64.99687, -64.95825, -64.91943, -64.88079, -64.84097, 
        -64.80189, -64.762, -64.72126, -64.67946, -64.63652, -64.5928, 
        -64.54819, -64.50269, -64.45596, -64.40796, -64.35904, -64.30937, 
        -64.25917, -64.20886, -64.1577, -64.10532, -64.05186, -63.99727, 
        -63.94154, -63.88466, -63.82636, -63.76617, -63.70344, -63.63796, 
        -63.56985, -63.49925, -63.42671, -63.35214, -63.27601, -63.19883, 
        -63.12109, -63.04343, -62.9666, -62.88979, -62.81508, -62.74087, 
        -62.66648, -62.59103, -62.51407, -62.4355, -62.35559, -62.27486, 
        -62.19381, -62.1131, -62.03321, -61.95428, -61.87617, -61.79805, 
        -61.71933, -61.63975, -61.55887, -61.47699, -61.39447, -61.31225, 
        -61.23111, -61.15147, -61.0736, -60.99748, -60.92304, -60.85015, 
        -60.77888, -60.70954, -60.64206, -60.57635, -60.51181, -60.44811, 
        -60.38532, -60.32397, -60.26458, -60.20762, -60.15328, -60.10155, 
        -60.05257, -60.00608, -59.96228, -59.92065, -59.88099, -59.8426, 
        -59.80427, -59.76735, -59.73101, -59.6949, -59.65918, -59.6238, 
        -59.59025,
  -49.12113, -49.14173, -49.17397, -49.2164, -49.26763, -49.32713, 
        -49.39489, -49.47175, -49.55933, -49.65992, -49.77529, -49.90958, 
        -50.06318, -50.23633, -50.42869, -50.6383, -50.86321, -51.1019, 
        -51.35151, -51.60973, -51.87447, -52.14338, -52.41518, -52.68907, 
        -52.96416, -53.23951, -53.51716, -53.79589, -54.07512, -54.35413, 
        -54.63209, -54.90736, -55.17804, -55.44207, -55.69719, -55.94153, 
        -56.17356, -56.39186, -56.59631, -56.78737, -56.96663, -57.13539, 
        -57.29863, -57.45832, -57.61715, -57.77698, -57.93862, -58.10168, 
        -58.26542, -58.42791, -58.58703, -58.7408, -58.88707, -59.0246, 
        -59.15332, -59.27314, -59.38534, -59.49001, -59.58976, -59.68439, 
        -59.77475, -59.86153, -59.94542, -60.02671, -60.10569, -60.18281, 
        -60.25853, -60.33322, -60.40685, -60.47951, -60.55135, -60.62272, 
        -60.69354, -60.76379, -60.83224, -60.90152, -60.97088, -61.04059, 
        -61.11116, -61.18274, -61.25583, -61.33032, -61.40637, -61.48348, 
        -61.56115, -61.63892, -61.71679, -61.79475, -61.8732, -61.9527, 
        -62.03376, -62.1166, -62.20117, -62.2865, -62.37423, -62.46293, 
        -62.5523, -62.64162, -62.73034, -62.81797, -62.90419, -62.98904, 
        -63.07268, -63.15515, -63.23688, -63.31726, -63.39589, -63.47274, 
        -63.54813, -63.62213, -63.69471, -63.76632, -63.83618, -63.90652, 
        -63.9767, -64.04684, -64.11675, -64.18623, -64.25455, -64.321, 
        -64.38523, -64.4471, -64.5069, -64.56503, -64.62254, -64.67996, 
        -64.73739, -64.7953, -64.85334, -64.91159, -64.96979, -65.02731, 
        -65.08306, -65.13861, -65.19286, -65.24599, -65.29758, -65.34784, 
        -65.39679, -65.44453, -65.49134, -65.53732, -65.5827, -65.62737, 
        -65.67159, -65.71522, -65.75831, -65.80143, -65.84404, -65.88614, 
        -65.9276, -65.96753, -66.00561, -66.03992, -66.07232, -66.10172, 
        -66.12806, -66.15167, -66.17242, -66.19057, -66.20632, -66.22005, 
        -66.23188, -66.24173, -66.2494, -66.25429, -66.25571, -66.25364, 
        -66.24812, -66.23975, -66.22881, -66.21612, -66.20212, -66.1867, 
        -66.17014, -66.1536, -66.13772, -66.12167, -66.10772, -66.09467, 
        -66.08179, -66.06853, -66.05459, -66.03914, -66.02186, -66.00231, 
        -65.98032, -65.95587, -65.92909, -65.90043, -65.87047, -65.83967, 
        -65.80859, -65.77724, -65.74537, -65.71287, -65.67999, -65.64651, 
        -65.61204, -65.57681, -65.54105, -65.50481, -65.46832, -65.43185, 
        -65.39431, -65.35802, -65.32178, -65.28577, -65.24924, -65.21217, 
        -65.17445, -65.13628, -65.09762, -65.05878, -65.01997, -64.98093, 
        -64.94138, -64.90124, -64.86005, -64.81766, -64.77428, -64.72992, 
        -64.68488, -64.63895, -64.59209, -64.54427, -64.49556, -64.44645, 
        -64.3968, -64.34672, -64.29585, -64.24381, -64.19086, -64.13657, 
        -64.08113, -64.02446, -63.9653, -63.90512, -63.8424, -63.77701, 
        -63.70884, -63.63826, -63.56556, -63.49089, -63.41433, -63.33643, 
        -63.25804, -63.17976, -63.10231, -63.02635, -62.95166, -62.87767, 
        -62.80366, -62.72873, -62.65204, -62.5737, -62.49383, -62.41314, 
        -62.3324, -62.2521, -62.17271, -62.0943, -62.01659, -61.93901, 
        -61.86076, -61.7813, -61.70041, -61.61839, -61.53569, -61.453, 
        -61.37124, -61.29065, -61.2119, -61.13497, -61.05894, -60.98561, 
        -60.91514, -60.8447, -60.77726, -60.71144, -60.64687, -60.58314, 
        -60.52037, -60.45914, -60.39992, -60.34319, -60.28936, -60.23852, 
        -60.1906, -60.1455, -60.10298, -60.06277, -60.02441, -59.98754, 
        -59.95159, -59.91591, -59.88058, -59.84593, -59.81176, -59.77824, 
        -59.74579,
  -49.35693, -49.38748, -49.42629, -49.47278, -49.52589, -49.58494, 
        -49.65302, -49.731, -49.82074, -49.92487, -50.0462, -50.18634, 
        -50.34651, -50.52626, -50.7244, -50.93863, -51.16671, -51.40674, 
        -51.65633, -51.91304, -52.17408, -52.43973, -52.70778, -52.97762, 
        -53.24841, -53.5202, -53.79321, -54.0671, -54.34154, -54.61627, 
        -54.89053, -55.16339, -55.43326, -55.69828, -55.95584, -56.20304, 
        -56.4396, -56.66288, -56.87212, -57.06758, -57.25034, -57.4226, 
        -57.58747, -57.74815, -57.90707, -58.06623, -58.22679, -58.3886, 
        -58.55078, -58.71177, -58.86956, -59.02094, -59.16632, -59.30341, 
        -59.43201, -59.55245, -59.6653, -59.7717, -59.87239, -59.9679, 
        -60.05903, -60.14655, -60.23085, -60.31271, -60.39228, -60.47021, 
        -60.54677, -60.62235, -60.69617, -60.77018, -60.84313, -60.91554, 
        -60.98731, -61.05871, -61.12952, -61.19963, -61.2696, -61.33979, 
        -61.41066, -61.48269, -61.55592, -61.63048, -61.70636, -61.78305, 
        -61.86036, -61.93783, -62.01433, -62.09175, -62.16962, -62.24838, 
        -62.32862, -62.41074, -62.4952, -62.58165, -62.66994, -62.75941, 
        -62.84951, -62.93956, -63.029, -63.11752, -63.20469, -63.29064, 
        -63.37571, -63.45985, -63.54348, -63.62463, -63.70541, -63.78447, 
        -63.86157, -63.93764, -64.01195, -64.08452, -64.1556, -64.22563, 
        -64.29498, -64.36407, -64.43304, -64.50173, -64.56921, -64.63524, 
        -64.6993, -64.76136, -64.82106, -64.87888, -64.93569, -64.99043, 
        -65.04585, -65.10095, -65.1561, -65.21158, -65.26743, -65.32316, 
        -65.37824, -65.43275, -65.48618, -65.5384, -65.58932, -65.63888, 
        -65.68707, -65.734, -65.77958, -65.82405, -65.86798, -65.91137, 
        -65.95467, -65.99669, -66.03913, -66.08093, -66.12183, -66.16209, 
        -66.20149, -66.23962, -66.27666, -66.31154, -66.34379, -66.37298, 
        -66.3993, -66.42248, -66.44246, -66.45972, -66.47388, -66.48547, 
        -66.49462, -66.50159, -66.50611, -66.50764, -66.50592, -66.50049, 
        -66.49079, -66.47909, -66.4649, -66.44865, -66.43098, -66.41204, 
        -66.39246, -66.37291, -66.35354, -66.33532, -66.31796, -66.30138, 
        -66.28507, -66.26831, -66.25038, -66.2307, -66.2088, -66.18444, 
        -66.15746, -66.12799, -66.09637, -66.06311, -66.02879, -65.99382, 
        -65.95879, -65.9236, -65.88745, -65.8518, -65.81568, -65.77918, 
        -65.74244, -65.70506, -65.66727, -65.62994, -65.59267, -65.55551, 
        -65.51868, -65.48239, -65.4468, -65.41114, -65.37521, -65.33892, 
        -65.30198, -65.26445, -65.22633, -65.18762, -65.14861, -65.10925, 
        -65.06933, -65.02858, -64.98701, -64.94432, -64.9005, -64.85562, 
        -64.80975, -64.76316, -64.71503, -64.66722, -64.6189, -64.57009, 
        -64.52099, -64.47131, -64.42068, -64.36892, -64.31583, -64.26157, 
        -64.20595, -64.14912, -64.09065, -64.0301, -63.96703, -63.90141, 
        -63.83321, -63.76279, -63.6902, -63.61534, -63.53842, -63.45998, 
        -63.38071, -63.30167, -63.22375, -63.14753, -63.07296, -62.99906, 
        -62.92517, -62.85028, -62.77382, -62.69558, -62.61587, -62.53535, 
        -62.45477, -62.37375, -62.29483, -62.21687, -62.13951, -62.06208, 
        -61.98399, -61.90439, -61.82334, -61.74099, -61.6578, -61.57462, 
        -61.49199, -61.41042, -61.33047, -61.25248, -61.17651, -61.10269, 
        -61.03094, -60.96124, -60.8934, -60.82729, -60.76255, -60.69897, 
        -60.63643, -60.57569, -60.51736, -60.46164, -60.40888, -60.3593, 
        -60.31261, -60.26872, -60.22757, -60.18873, -60.1518, -60.1162, 
        -60.08172, -60.04769, -60.01411, -59.98087, -59.94799, -59.91594, 
        -59.88485,
  -49.5916, -49.6306, -49.67539, -49.72542, -49.78069, -49.84185, 
        -49.91121, -49.99113, -50.08401, -50.19271, -50.31961, -50.4662, 
        -50.63269, -50.81857, -51.02185, -51.23889, -51.46917, -51.7098, 
        -51.9586, -52.21339, -52.47258, -52.73459, -52.99884, -53.26487, 
        -53.53167, -53.79949, -54.06863, -54.33864, -54.60928, -54.88039, 
        -55.15073, -55.4217, -55.69116, -55.95708, -56.21693, -56.46827, 
        -56.70869, -56.93622, -57.14949, -57.3487, -57.53453, -57.70942, 
        -57.87607, -58.0375, -58.19649, -58.35498, -58.5132, -58.67304, 
        -58.83273, -58.99094, -59.14591, -59.29584, -59.43901, -59.57469, 
        -59.70238, -59.82238, -59.93531, -60.04227, -60.14345, -60.23943, 
        -60.33103, -60.41877, -60.50253, -60.58472, -60.66491, -60.74339, 
        -60.82085, -60.89738, -60.97321, -61.04823, -61.12238, -61.19589, 
        -61.2684, -61.34091, -61.41262, -61.48381, -61.55441, -61.62526, 
        -61.69672, -61.76819, -61.84171, -61.91673, -61.99261, -62.06945, 
        -62.14654, -62.22382, -62.30092, -62.37788, -62.45519, -62.53311, 
        -62.61274, -62.69409, -62.77802, -62.86457, -62.95321, -63.04338, 
        -63.13413, -63.22471, -63.31371, -63.40283, -63.49075, -63.57778, 
        -63.66422, -63.74995, -63.83484, -63.91881, -64.0013, -64.08199, 
        -64.16136, -64.23911, -64.31488, -64.38851, -64.45979, -64.52934, 
        -64.59775, -64.6656, -64.73212, -64.79916, -64.86536, -64.93061, 
        -64.99416, -65.05613, -65.11585, -65.17373, -65.22984, -65.28442, 
        -65.33804, -65.39095, -65.44389, -65.49706, -65.55058, -65.60466, 
        -65.6584, -65.71187, -65.76428, -65.81554, -65.86543, -65.91287, 
        -65.95982, -66.00542, -66.04958, -66.0929, -66.13581, -66.17839, 
        -66.22123, -66.26401, -66.30582, -66.34624, -66.38534, -66.42352, 
        -66.46095, -66.49773, -66.53355, -66.56785, -66.59994, -66.62916, 
        -66.65536, -66.67843, -66.6981, -66.71445, -66.72643, -66.73615, 
        -66.74303, -66.74734, -66.74875, -66.74722, -66.74232, -66.73387, 
        -66.7216, -66.70665, -66.68918, -66.66954, -66.64818, -66.62571, 
        -66.60297, -66.58004, -66.5576, -66.53597, -66.51543, -66.49568, 
        -66.47598, -66.45576, -66.43402, -66.41008, -66.38367, -66.35345, 
        -66.32171, -66.28756, -66.2513, -66.21351, -66.17477, -66.13559, 
        -66.09657, -66.05771, -66.01881, -65.97987, -65.94055, -65.90101, 
        -65.8614, -65.8215, -65.78176, -65.74265, -65.70412, -65.66624, 
        -65.62906, -65.5928, -65.55753, -65.52271, -65.48792, -65.45267, 
        -65.41682, -65.3801, -65.3426, -65.3031, -65.26384, -65.22391, 
        -65.18337, -65.14239, -65.10069, -65.05794, -65.01395, -64.96848, 
        -64.9217, -64.87424, -64.82648, -64.77847, -64.73034, -64.68211, 
        -64.63346, -64.58409, -64.53338, -64.48138, -64.42797, -64.37316, 
        -64.31714, -64.25964, -64.20036, -64.13915, -64.07561, -64.00969, 
        -63.94167, -63.87133, -63.79877, -63.72381, -63.64643, -63.56739, 
        -63.48639, -63.40668, -63.32821, -63.25161, -63.17667, -63.10271, 
        -63.02879, -62.95378, -62.87723, -62.79902, -62.7196, -62.63944, 
        -62.55931, -62.47985, -62.4015, -62.32401, -62.2467, -62.16922, 
        -62.09093, -62.01101, -61.92953, -61.84658, -61.76294, -61.67902, 
        -61.59546, -61.51291, -61.43167, -61.35236, -61.27541, -61.20074, 
        -61.12845, -61.05805, -60.98963, -60.92302, -60.85821, -60.79465, 
        -60.73293, -60.67336, -60.61624, -60.56208, -60.51086, -60.46194, 
        -60.41676, -60.37397, -60.33384, -60.29614, -60.26038, -60.22624, 
        -60.19335, -60.16095, -60.12914, -60.09757, -60.06654, -60.0362, 
        -60.00647,
  -49.81953, -49.86659, -49.91719, -49.97107, -50.02938, -50.09337, 
        -50.16532, -50.24843, -50.34566, -50.45872, -50.59185, -50.7448, 
        -50.91745, -51.1086, -51.31587, -51.53644, -51.76777, -52.00803, 
        -52.25483, -52.50665, -52.76219, -53.02059, -53.28102, -53.54306, 
        -53.80534, -54.07045, -54.33661, -54.60392, -54.87202, -55.14093, 
        -55.41076, -55.6809, -55.95033, -56.21724, -56.47919, -56.73317, 
        -56.97661, -57.20721, -57.42348, -57.62545, -57.81296, -57.98992, 
        -58.15824, -58.32087, -58.4801, -58.63811, -58.79571, -58.95317, 
        -59.10981, -59.26435, -59.41552, -59.56176, -59.70187, -59.83501, 
        -59.96097, -60.08003, -60.19177, -60.29843, -60.39977, -60.49603, 
        -60.5879, -60.67601, -60.7608, -60.84325, -60.9238, -61.00275, 
        -61.08087, -61.15836, -61.23524, -61.31133, -61.38667, -61.46092, 
        -61.53452, -61.60675, -61.67926, -61.75116, -61.82265, -61.89434, 
        -61.96638, -62.0393, -62.11335, -62.18888, -62.2653, -62.34243, 
        -62.41953, -62.49644, -62.57328, -62.64996, -62.72691, -62.80465, 
        -62.88371, -62.96379, -63.04746, -63.13401, -63.22265, -63.31301, 
        -63.40397, -63.49478, -63.58504, -63.67456, -63.7632, -63.85105, 
        -63.93844, -64.02524, -64.11137, -64.19653, -64.28046, -64.36319, 
        -64.44437, -64.52296, -64.60012, -64.67455, -64.74599, -64.81502, 
        -64.88249, -64.94899, -65.01503, -65.0802, -65.14497, -65.20898, 
        -65.27175, -65.33306, -65.39235, -65.4501, -65.5057, -65.55932, 
        -65.61161, -65.66293, -65.71397, -65.76535, -65.81625, -65.86869, 
        -65.9213, -65.97359, -66.02518, -66.07557, -66.12452, -66.17181, 
        -66.21782, -66.26219, -66.30556, -66.34783, -66.38963, -66.43195, 
        -66.47414, -66.51611, -66.55703, -66.59624, -66.63415, -66.67077, 
        -66.70657, -66.74068, -66.77528, -66.80879, -66.84028, -66.8694, 
        -66.89568, -66.91872, -66.93798, -66.95367, -66.96546, -66.97353, 
        -66.97809, -66.97971, -66.97821, -66.97363, -66.96574, -66.95411, 
        -66.93895, -66.92078, -66.90021, -66.87735, -66.85245, -66.82697, 
        -66.80109, -66.77449, -66.74911, -66.7244, -66.70064, -66.67746, 
        -66.65437, -66.63039, -66.60464, -66.57652, -66.54564, -66.51208, 
        -66.47577, -66.43723, -66.39662, -66.35455, -66.31145, -66.26817, 
        -66.22504, -66.18246, -66.14001, -66.09749, -66.05487, -66.01205, 
        -65.96927, -65.92667, -65.88464, -65.84373, -65.80284, -65.76411, 
        -65.72661, -65.69028, -65.65519, -65.6209, -65.58679, -65.55254, 
        -65.51756, -65.48163, -65.44437, -65.406, -65.36646, -65.32616, 
        -65.28523, -65.24414, -65.20258, -65.15974, -65.11527, -65.06907, 
        -65.02153, -64.97341, -64.92502, -64.87665, -64.82864, -64.78066, 
        -64.73212, -64.68256, -64.63157, -64.57908, -64.52491, -64.46848, 
        -64.4116, -64.35318, -64.29317, -64.23115, -64.16739, -64.10154, 
        -64.03353, -63.96334, -63.89079, -63.81562, -63.73799, -63.65841, 
        -63.57761, -63.49692, -63.41773, -63.34027, -63.26456, -63.18983, 
        -63.1153, -63.04007, -62.96354, -62.88562, -62.80659, -62.72692, 
        -62.64739, -62.5685, -62.49047, -62.41315, -62.3361, -62.2583, 
        -62.17974, -62.09945, -62.01739, -61.93409, -61.84983, -61.76513, 
        -61.6807, -61.59601, -61.51349, -61.43317, -61.3551, -61.27945, 
        -61.2061, -61.13488, -61.06567, -60.99843, -60.93337, -60.87034, 
        -60.80952, -60.75117, -60.69571, -60.64332, -60.59404, -60.54784, 
        -60.50368, -60.46226, -60.42327, -60.38672, -60.3523, -60.31981, 
        -60.28868, -60.25835, -60.22848, -60.19878, -60.16953, -60.1408, 
        -60.11269,
  -50.03341, -50.0878, -50.1447, -50.2038, -50.26534, -50.33352, 
        -50.41008, -50.49832, -50.60142, -50.72177, -50.8615, -51.02078, 
        -51.199, -51.39456, -51.60456, -51.82658, -52.05769, -52.29579, 
        -52.53967, -52.7865, -53.03796, -53.29203, -53.54847, -53.80682, 
        -54.06775, -54.33014, -54.59455, -54.86048, -55.12774, -55.39616, 
        -55.66579, -55.93624, -56.20646, -56.47466, -56.73731, -56.99334, 
        -57.2387, -57.47113, -57.68919, -57.89285, -58.08319, -58.26189, 
        -58.43179, -58.59543, -58.7551, -58.91266, -59.06876, -59.22376, 
        -59.37709, -59.52761, -59.67348, -59.81548, -59.95164, -60.08162, 
        -60.2053, -60.32293, -60.43465, -60.54082, -60.64198, -60.73812, 
        -60.8301, -60.91822, -61.00312, -61.08553, -61.16609, -61.2455, 
        -61.32418, -61.40143, -61.47921, -61.55629, -61.63283, -61.70825, 
        -61.78282, -61.85654, -61.92975, -62.00257, -62.07486, -62.14727, 
        -62.22009, -62.29382, -62.36859, -62.44461, -62.52154, -62.5989, 
        -62.67613, -62.75219, -62.82894, -62.90553, -62.98232, -63.06006, 
        -63.13905, -63.21989, -63.30348, -63.38977, -63.47827, -63.56845, 
        -63.65935, -63.75027, -63.84045, -63.93001, -64.01906, -64.10746, 
        -64.19454, -64.28228, -64.36931, -64.4555, -64.54076, -64.62493, 
        -64.7079, -64.78886, -64.86745, -64.94254, -65.01449, -65.08321, 
        -65.14986, -65.21522, -65.27956, -65.34305, -65.40593, -65.46827, 
        -65.52975, -65.59022, -65.64846, -65.70565, -65.7604, -65.8134, 
        -65.86476, -65.9149, -65.96468, -66.01463, -66.06525, -66.11653, 
        -66.16825, -66.21964, -66.27032, -66.31971, -66.36771, -66.41427, 
        -66.4594, -66.50328, -66.54592, -66.58783, -66.62945, -66.66988, 
        -66.71131, -66.75238, -66.79237, -66.8307, -66.86716, -66.90234, 
        -66.93674, -66.97054, -67.00388, -67.03643, -67.06728, -67.09596, 
        -67.12196, -67.14455, -67.16346, -67.17833, -67.18905, -67.19544, 
        -67.1981, -67.197, -67.19232, -67.18477, -67.17419, -67.15897, 
        -67.14112, -67.12029, -67.09702, -67.07141, -67.04375, -67.01543, 
        -66.98689, -66.9586, -66.93044, -66.9028, -66.87571, -66.84905, 
        -66.82217, -66.79434, -66.76453, -66.73225, -66.69713, -66.65922, 
        -66.61868, -66.57577, -66.53101, -66.48471, -66.43759, -66.39016, 
        -66.3422, -66.2957, -66.24952, -66.20338, -66.15733, -66.1111, 
        -66.06496, -66.01947, -65.97517, -65.93234, -65.89128, -65.85187, 
        -65.81419, -65.77787, -65.74272, -65.70865, -65.67459, -65.6406, 
        -65.60616, -65.57045, -65.53353, -65.49481, -65.4549, -65.41429, 
        -65.37333, -65.33203, -65.29026, -65.24714, -65.2023, -65.15462, 
        -65.10656, -65.05745, -65.00822, -64.95959, -64.91129, -64.86313, 
        -64.81427, -64.76439, -64.71291, -64.65971, -64.60483, -64.5485, 
        -64.49076, -64.43155, -64.37083, -64.30836, -64.24434, -64.1784, 
        -64.11083, -64.04086, -63.96841, -63.89293, -63.81497, -63.7347, 
        -63.65316, -63.57153, -63.49109, -63.41229, -63.33524, -63.25932, 
        -63.18399, -63.10814, -63.03144, -62.95385, -62.87435, -62.79541, 
        -62.71658, -62.63824, -62.56076, -62.48357, -62.4062, -62.32822, 
        -62.24907, -62.16856, -62.08605, -62.00219, -61.91727, -61.8318, 
        -61.74646, -61.66174, -61.57828, -61.49669, -61.41741, -61.34055, 
        -61.26616, -61.19399, -61.12403, -61.05634, -60.99118, -60.92854, 
        -60.86873, -60.81188, -60.75826, -60.70778, -60.6604, -60.61581, 
        -60.57329, -60.53289, -60.49488, -60.45918, -60.42624, -60.39554, 
        -60.36653, -60.33829, -60.3104, -60.2827, -60.25526, -60.22816, 
        -60.20192,
  -50.22653, -50.28865, -50.35238, -50.41823, -50.4872, -50.5616, 
        -50.64447, -50.73957, -50.84975, -50.97718, -51.1235, -51.28873, 
        -51.47175, -51.66977, -51.88194, -52.10413, -52.33366, -52.56886, 
        -52.80875, -53.05209, -53.29885, -53.54846, -53.80102, -54.05639, 
        -54.3148, -54.57581, -54.83929, -55.10479, -55.37257, -55.64096, 
        -55.91172, -56.18344, -56.45512, -56.72482, -56.98978, -57.2468, 
        -57.493, -57.72596, -57.94453, -58.14895, -58.34015, -58.52013, 
        -58.69124, -58.85585, -59.015, -59.17217, -59.3271, -59.47979, 
        -59.6297, -59.77627, -59.91859, -60.05592, -60.1879, -60.31427, 
        -60.43523, -60.55103, -60.66147, -60.76684, -60.86742, -60.96342, 
        -61.05512, -61.14212, -61.22683, -61.3091, -61.38959, -61.46918, 
        -61.54825, -61.62719, -61.70582, -61.78404, -61.86144, -61.93782, 
        -62.01331, -62.08789, -62.16197, -62.23563, -62.30876, -62.38103, 
        -62.45475, -62.52926, -62.60483, -62.68138, -62.75874, -62.83664, 
        -62.91428, -62.99152, -63.06828, -63.14502, -63.22196, -63.29968, 
        -63.37888, -63.46, -63.54354, -63.62953, -63.71746, -63.80613, 
        -63.8964, -63.98691, -64.07719, -64.16685, -64.25591, -64.3448, 
        -64.43324, -64.52122, -64.60885, -64.69587, -64.78238, -64.86813, 
        -64.95227, -65.03472, -65.11427, -65.1902, -65.2625, -65.33144, 
        -65.3978, -65.46124, -65.52414, -65.58598, -65.64711, -65.70764, 
        -65.7679, -65.82722, -65.88549, -65.94189, -65.99625, -66.04847, 
        -66.09917, -66.14886, -66.19791, -66.24702, -66.29666, -66.34692, 
        -66.39784, -66.44839, -66.49804, -66.54658, -66.59253, -66.63844, 
        -66.68313, -66.72691, -66.76974, -66.81164, -66.85329, -66.89445, 
        -66.93526, -66.97528, -67.01411, -67.0512, -67.08671, -67.12088, 
        -67.15406, -67.18631, -67.21806, -67.2491, -67.27878, -67.30647, 
        -67.33147, -67.35361, -67.37093, -67.38512, -67.39456, -67.39931, 
        -67.40011, -67.39685, -67.38979, -67.37959, -67.36636, -67.34991, 
        -67.32969, -67.30637, -67.28073, -67.25279, -67.2232, -67.19294, 
        -67.16228, -67.13175, -67.10121, -67.07069, -67.0404, -67.01011, 
        -66.97921, -66.94714, -66.91316, -66.87525, -66.83585, -66.79388, 
        -66.74932, -66.70272, -66.65411, -66.60358, -66.55218, -66.50072, 
        -66.44991, -66.39974, -66.34985, -66.30009, -66.25028, -66.20034, 
        -66.15105, -66.10242, -66.05557, -66.01081, -65.96837, -65.92831, 
        -65.89027, -65.85389, -65.81872, -65.78438, -65.75027, -65.71594, 
        -65.68105, -65.64413, -65.60677, -65.56783, -65.5279, -65.48706, 
        -65.4459, -65.40443, -65.36217, -65.31856, -65.2731, -65.22562, 
        -65.17659, -65.12679, -65.07726, -65.02813, -64.97914, -64.93031, 
        -64.88105, -64.83057, -64.77841, -64.72443, -64.66882, -64.61191, 
        -64.55357, -64.49374, -64.43235, -64.36961, -64.30549, -64.24, 
        -64.17261, -64.10276, -64.03036, -63.95383, -63.8755, -63.79456, 
        -63.71225, -63.62971, -63.54773, -63.46709, -63.38813, -63.31055, 
        -63.23408, -63.15753, -63.08066, -63.0031, -62.9249, -62.84654, 
        -62.76834, -62.69062, -62.6133, -62.53596, -62.45858, -62.38034, 
        -62.30085, -62.21986, -62.13708, -62.05288, -61.96742, -61.88127, 
        -61.79508, -61.70939, -61.62487, -61.54207, -61.46147, -61.38334, 
        -61.30779, -61.23469, -61.16411, -61.09638, -61.03157, -60.96972, 
        -60.91099, -60.85552, -60.80256, -60.75398, -60.70842, -60.66528, 
        -60.62416, -60.58489, -60.54781, -60.51351, -60.48214, -60.45319, 
        -60.4263, -60.40029, -60.37454, -60.34863, -60.32312, -60.29794, 
        -60.27354,
  -50.39724, -50.46782, -50.53951, -50.61306, -50.69001, -50.77259, 
        -50.86393, -50.96724, -51.08432, -51.21933, -51.37217, -51.54283, 
        -51.72992, -51.93156, -52.14443, -52.36582, -52.59319, -52.82499, 
        -53.06075, -53.29974, -53.54194, -53.78758, -54.03675, -54.28843, 
        -54.54522, -54.80535, -55.06867, -55.33507, -55.60416, -55.87545, 
        -56.14826, -56.42189, -56.69522, -56.96595, -57.23154, -57.48866, 
        -57.73437, -57.96681, -58.18482, -58.38786, -58.57927, -58.75988, 
        -58.93166, -59.0969, -59.25732, -59.4143, -59.56807, -59.7187, 
        -59.8657, -60.00842, -60.14647, -60.27943, -60.4072, -60.53009, 
        -60.64816, -60.76084, -60.86976, -60.9742, -61.07419, -61.16991, 
        -61.26124, -61.34879, -61.4331, -61.51502, -61.5953, -61.67487, 
        -61.75406, -61.83331, -61.91264, -61.99162, -62.07014, -62.14672, 
        -62.22325, -62.29879, -62.37377, -62.4482, -62.52211, -62.59614, 
        -62.67078, -62.74631, -62.82283, -62.89999, -62.97784, -63.05601, 
        -63.1339, -63.21141, -63.28859, -63.36549, -63.44275, -63.52017, 
        -63.59988, -63.68144, -63.76494, -63.8505, -63.93787, -64.02654, 
        -64.11595, -64.20573, -64.2956, -64.38505, -64.47429, -64.56284, 
        -64.65145, -64.73953, -64.82747, -64.9152, -65.00278, -65.0895, 
        -65.174, -65.25731, -65.33775, -65.41461, -65.48745, -65.5567, 
        -65.62331, -65.68738, -65.74962, -65.81023, -65.8699, -65.92921, 
        -65.98817, -66.04652, -66.10371, -66.15929, -66.21298, -66.26466, 
        -66.31495, -66.3641, -66.41156, -66.46004, -66.50884, -66.55836, 
        -66.60838, -66.65794, -66.70683, -66.75474, -66.80156, -66.84718, 
        -66.89201, -66.93616, -66.97926, -67.02168, -67.06319, -67.10399, 
        -67.1441, -67.18306, -67.22053, -67.25638, -67.29069, -67.32396, 
        -67.35497, -67.3858, -67.41589, -67.44506, -67.47303, -67.49928, 
        -67.52293, -67.54379, -67.56094, -67.57439, -67.58298, -67.58666, 
        -67.58597, -67.58089, -67.57211, -67.55978, -67.54433, -67.52552, 
        -67.50306, -67.47765, -67.44965, -67.41969, -67.38831, -67.35623, 
        -67.32302, -67.29102, -67.25846, -67.2257, -67.19254, -67.15897, 
        -67.12437, -67.08841, -67.0503, -67.00907, -66.96531, -66.91908, 
        -66.87065, -66.82029, -66.76763, -66.71343, -66.65835, -66.60284, 
        -66.54784, -66.49354, -66.43969, -66.38595, -66.33247, -66.2791, 
        -66.22645, -66.17507, -66.12463, -66.07771, -66.03375, -65.99226, 
        -65.95317, -65.91595, -65.88033, -65.84547, -65.81053, -65.77574, 
        -65.74032, -65.70372, -65.66602, -65.62691, -65.58673, -65.54573, 
        -65.50429, -65.46232, -65.41947, -65.3751, -65.32863, -65.28027, 
        -65.23056, -65.18017, -65.12991, -65.07995, -65.03038, -64.98087, 
        -64.93082, -64.87954, -64.82664, -64.77106, -64.71497, -64.65742, 
        -64.59873, -64.53862, -64.47702, -64.41425, -64.3503, -64.28511, 
        -64.21808, -64.14864, -64.07625, -64.00046, -63.92178, -63.84018, 
        -63.75694, -63.67284, -63.58919, -63.50677, -63.42587, -63.34677, 
        -63.26884, -63.19156, -63.11427, -63.03642, -62.95829, -62.87993, 
        -62.80161, -62.72384, -62.64631, -62.56879, -62.49078, -62.41201, 
        -62.33246, -62.2514, -62.16884, -62.08466, -61.99807, -61.91162, 
        -61.8249, -61.73829, -61.6527, -61.56859, -61.48655, -61.40691, 
        -61.33011, -61.25635, -61.18552, -61.11821, -61.0542, -60.99335, 
        -60.93597, -60.88197, -60.83152, -60.78441, -60.74035, -60.69879, 
        -60.6589, -60.62104, -60.5854, -60.55249, -60.52255, -60.49547, 
        -60.47044, -60.4461, -60.4223, -60.39867, -60.37527, -60.35245, 
        -60.32991,
  -50.54191, -50.62176, -50.70222, -50.78378, -50.87004, -50.96223, 
        -51.06332, -51.17604, -51.30284, -51.44549, -51.60472, -51.78001, 
        -51.97054, -52.1739, -52.38715, -52.60728, -52.83217, -53.0606, 
        -53.2916, -53.52657, -53.76493, -54.00721, -54.25372, -54.50445, 
        -54.76007, -55.02021, -55.28417, -55.55205, -55.82334, -56.09706, 
        -56.3725, -56.64826, -56.92303, -57.19339, -57.45849, -57.71447, 
        -57.95864, -58.1892, -58.40558, -58.60842, -58.79919, -58.97964, 
        -59.15174, -59.31731, -59.4779, -59.63451, -59.78745, -59.93629, 
        -60.08075, -60.21927, -60.35351, -60.48258, -60.60674, -60.72634, 
        -60.84174, -60.95327, -61.06085, -61.16421, -61.26339, -61.35841, 
        -61.44925, -61.53617, -61.61996, -61.7014, -61.78131, -61.85944, 
        -61.93854, -62.01794, -62.09764, -62.17727, -62.2568, -62.33556, 
        -62.4131, -62.48959, -62.56533, -62.6404, -62.71542, -62.79042, 
        -62.86623, -62.94274, -63.02028, -63.09823, -63.17548, -63.25389, 
        -63.33212, -63.41002, -63.48772, -63.56539, -63.6435, -63.72271, 
        -63.80295, -63.88517, -63.96872, -64.05388, -64.14036, -64.22786, 
        -64.31602, -64.40464, -64.49362, -64.5826, -64.67139, -64.75894, 
        -64.84741, -64.93573, -65.02393, -65.11236, -65.20068, -65.28818, 
        -65.37425, -65.45821, -65.53931, -65.61691, -65.6904, -65.76054, 
        -65.82748, -65.89187, -65.95396, -66.01414, -66.07326, -66.1316, 
        -66.18919, -66.2453, -66.30148, -66.35632, -66.4095, -66.46066, 
        -66.51054, -66.55914, -66.60705, -66.65487, -66.70294, -66.75178, 
        -66.80102, -66.84997, -66.89851, -66.94601, -66.993, -67.03887, 
        -67.08413, -67.12894, -67.17248, -67.21527, -67.25598, -67.29652, 
        -67.33583, -67.37357, -67.40977, -67.44441, -67.47762, -67.50967, 
        -67.54026, -67.56993, -67.59852, -67.62595, -67.65192, -67.67634, 
        -67.69858, -67.71787, -67.73375, -67.74564, -67.75327, -67.75595, 
        -67.75408, -67.74796, -67.73776, -67.7228, -67.7054, -67.68446, 
        -67.66013, -67.63269, -67.60255, -67.5711, -67.53834, -67.50499, 
        -67.47158, -67.43803, -67.40414, -67.36904, -67.33315, -67.2966, 
        -67.2585, -67.21894, -67.17716, -67.13223, -67.08456, -67.03476, 
        -66.98266, -66.92828, -66.87185, -66.81353, -66.75354, -66.69434, 
        -66.63548, -66.5771, -66.51908, -66.4612, -66.40394, -66.34715, 
        -66.29141, -66.23719, -66.18523, -66.13619, -66.09, -66.04666, 
        -66.00591, -65.96717, -65.93, -65.89377, -65.85774, -65.82173, 
        -65.78532, -65.74823, -65.71019, -65.67094, -65.63058, -65.58929, 
        -65.54745, -65.50468, -65.46084, -65.41431, -65.36683, -65.31776, 
        -65.26723, -65.21633, -65.16529, -65.11465, -65.06413, -65.01356, 
        -64.9626, -64.91041, -64.85683, -64.80175, -64.74529, -64.68752, 
        -64.62852, -64.56816, -64.50679, -64.44413, -64.38045, -64.31548, 
        -64.24879, -64.17958, -64.10709, -64.03137, -63.95204, -63.86975, 
        -63.78543, -63.70013, -63.61487, -63.53046, -63.44773, -63.367, 
        -63.28782, -63.20868, -63.13049, -63.05205, -62.9733, -62.89461, 
        -62.81599, -62.73751, -62.65922, -62.581, -62.50232, -62.42312, 
        -62.34327, -62.26235, -62.18022, -62.09651, -62.01122, -61.92461, 
        -61.83751, -61.75044, -61.66385, -61.57853, -61.49497, -61.41401, 
        -61.3362, -61.26186, -61.19124, -61.12471, -61.06198, -61.00289, 
        -60.94719, -60.89484, -60.84578, -60.8001, -60.75726, -60.71687, 
        -60.67846, -60.64188, -60.60757, -60.57616, -60.54776, -60.52238, 
        -60.49863, -60.47633, -60.45471, -60.4334, -60.41077, -60.39027, 
        -60.3705,
  -50.65763, -50.74757, -50.83794, -50.93007, -51.02643, -51.12919, 
        -51.24059, -51.36316, -51.49903, -51.6493, -51.81456, -51.99451, 
        -52.18639, -52.39089, -52.60403, -52.82299, -53.04566, -53.27132, 
        -53.50027, -53.73247, -53.96826, -54.20837, -54.45321, -54.70301, 
        -54.95832, -55.21912, -55.4845, -55.75338, -56.02731, -56.30377, 
        -56.58158, -56.85919, -57.13485, -57.40593, -57.6695, -57.92323, 
        -58.16448, -58.39209, -58.60593, -58.80685, -58.99631, -59.17602, 
        -59.3468, -59.5124, -59.67302, -59.82921, -59.98125, -60.12872, 
        -60.27108, -60.40791, -60.53912, -60.6651, -60.78625, -60.9031, 
        -61.01632, -61.12596, -61.23217, -61.33467, -61.43309, -61.52627, 
        -61.61634, -61.70259, -61.78547, -61.86624, -61.94558, -62.02412, 
        -62.10291, -62.18225, -62.26227, -62.34242, -62.42241, -62.502, 
        -62.58041, -62.65778, -62.7342, -62.81013, -62.88519, -62.9615, 
        -63.03852, -63.11638, -63.19469, -63.27344, -63.35223, -63.431, 
        -63.50968, -63.58827, -63.66689, -63.74557, -63.82476, -63.90505, 
        -63.98659, -64.06918, -64.15308, -64.23782, -64.32216, -64.40833, 
        -64.49493, -64.58198, -64.66978, -64.75789, -64.8463, -64.93473, 
        -65.02296, -65.11156, -65.20036, -65.28931, -65.37779, -65.46555, 
        -65.55186, -65.63592, -65.71745, -65.7956, -65.86998, -65.94016, 
        -66.00789, -66.07286, -66.13537, -66.19582, -66.25466, -66.31217, 
        -66.36898, -66.4249, -66.4802, -66.53448, -66.58717, -66.63811, 
        -66.6875, -66.73566, -66.78309, -66.83037, -66.87798, -66.92604, 
        -66.97476, -67.02369, -67.07143, -67.11941, -67.16692, -67.2134, 
        -67.25939, -67.30482, -67.34936, -67.39243, -67.43413, -67.47425, 
        -67.51266, -67.54921, -67.58419, -67.61759, -67.65003, -67.68091, 
        -67.71053, -67.73865, -67.76571, -67.79148, -67.81555, -67.83816, 
        -67.85748, -67.87478, -67.88892, -67.89923, -67.90539, -67.90698, 
        -67.90392, -67.89676, -67.88541, -67.87006, -67.85092, -67.82806, 
        -67.80169, -67.77235, -67.74093, -67.70802, -67.67434, -67.64034, 
        -67.60597, -67.57104, -67.53527, -67.49816, -67.45999, -67.42066, 
        -67.37976, -67.33585, -67.2905, -67.24236, -67.19147, -67.13845, 
        -67.08312, -67.02512, -66.96511, -66.90311, -66.84033, -66.77721, 
        -66.71432, -66.6519, -66.58999, -66.52858, -66.46772, -66.40762, 
        -66.34885, -66.29164, -66.23694, -66.18503, -66.13628, -66.09058, 
        -66.04745, -66.00659, -65.96739, -65.92908, -65.8903, -65.85284, 
        -65.81519, -65.7774, -65.73875, -65.69909, -65.6585, -65.6169, 
        -65.57433, -65.53064, -65.48567, -65.43877, -65.39019, -65.33993, 
        -65.28885, -65.23739, -65.18597, -65.13461, -65.08299, -65.0312, 
        -64.9791, -64.92592, -64.87158, -64.81595, -64.75911, -64.70125, 
        -64.64205, -64.58183, -64.52044, -64.45796, -64.39463, -64.33002, 
        -64.26252, -64.19336, -64.12081, -64.04462, -63.96481, -63.88172, 
        -63.7965, -63.70977, -63.62313, -63.53736, -63.45324, -63.37099, 
        -63.29047, -63.21112, -63.13201, -63.05268, -62.973, -62.89331, 
        -62.81387, -62.73444, -62.6549, -62.57543, -62.49574, -62.416, 
        -62.33598, -62.25536, -62.1736, -62.09026, -62.0054, -61.91903, 
        -61.8318, -61.74437, -61.65714, -61.57098, -61.4865, -61.4046, 
        -61.32612, -61.25164, -61.18174, -61.11636, -61.05437, -60.99721, 
        -60.94346, -60.89299, -60.84563, -60.80148, -60.76004, -60.72101, 
        -60.68373, -60.64857, -60.61563, -60.58541, -60.5582, -60.53374, 
        -60.51149, -60.49075, -60.47086, -60.45181, -60.433, -60.41473, 
        -60.39747,
  -50.74575, -50.84604, -50.94658, -51.04889, -51.15512, -51.26838, 
        -51.39031, -51.52187, -51.66684, -51.82468, -51.99583, -52.17985, 
        -52.37505, -52.58027, -52.79305, -53.01108, -53.23223, -53.45624, 
        -53.68336, -53.91396, -54.1487, -54.3883, -54.63192, -54.88235, 
        -55.13848, -55.40079, -55.66827, -55.94043, -56.2168, -56.49553, 
        -56.77532, -57.05417, -57.32989, -57.59956, -57.86064, -58.11077, 
        -58.34823, -58.57108, -58.78176, -58.98019, -59.16776, -59.34615, 
        -59.51714, -59.68216, -59.84233, -59.99821, -60.14954, -60.29594, 
        -60.43648, -60.57128, -60.70021, -60.82389, -60.94283, -61.05673, 
        -61.16801, -61.27637, -61.38148, -61.48309, -61.58074, -61.67427, 
        -61.76355, -61.84885, -61.93076, -62.0106, -62.08918, -62.16752, 
        -62.24619, -62.3253, -62.40504, -62.4852, -62.56447, -62.64445, 
        -62.72334, -62.80119, -62.87811, -62.95504, -63.03228, -63.11, 
        -63.18844, -63.26747, -63.34693, -63.42645, -63.50592, -63.58535, 
        -63.66486, -63.74432, -63.82409, -63.90417, -63.98409, -64.0657, 
        -64.14848, -64.23201, -64.31616, -64.40054, -64.48485, -64.56934, 
        -64.65426, -64.73977, -64.82605, -64.91318, -65.00099, -65.08932, 
        -65.1778, -65.26663, -65.35588, -65.4451, -65.53267, -65.62021, 
        -65.70621, -65.79019, -65.87175, -65.95036, -66.02563, -66.09776, 
        -66.16647, -66.23235, -66.29572, -66.35652, -66.41531, -66.47249, 
        -66.52885, -66.58417, -66.63881, -66.69268, -66.74542, -66.79633, 
        -66.84495, -66.89309, -66.94045, -66.98718, -67.03444, -67.08235, 
        -67.13099, -67.18015, -67.22952, -67.27862, -67.32671, -67.37424, 
        -67.42059, -67.46686, -67.51208, -67.55532, -67.59682, -67.63633, 
        -67.67369, -67.70932, -67.74313, -67.77548, -67.80608, -67.83631, 
        -67.86536, -67.89265, -67.91818, -67.942, -67.96404, -67.9844, 
        -68.00252, -68.01774, -68.02975, -68.03808, -68.04261, -68.04288, 
        -68.03859, -68.03009, -68.01733, -68.00085, -67.98022, -67.95554, 
        -67.92735, -67.89627, -67.86358, -67.82987, -67.79467, -67.76001, 
        -67.72462, -67.68845, -67.65104, -67.61191, -67.57166, -67.5297, 
        -67.4863, -67.44075, -67.39259, -67.34163, -67.2881, -67.23219, 
        -67.17366, -67.11233, -67.04886, -66.98335, -66.91683, -66.84997, 
        -66.78307, -66.71664, -66.65103, -66.58618, -66.52234, -66.45959, 
        -66.39697, -66.33707, -66.27938, -66.22443, -66.17239, -66.12347, 
        -66.07712, -66.03326, -65.99115, -65.95058, -65.91106, -65.87196, 
        -65.83318, -65.79434, -65.75494, -65.71462, -65.67326, -65.63069, 
        -65.58705, -65.54231, -65.49599, -65.44779, -65.39803, -65.34689, 
        -65.29507, -65.243, -65.19096, -65.13889, -65.0864, -65.03351, 
        -64.9791, -64.92478, -64.8697, -64.81339, -64.75603, -64.69775, 
        -64.63856, -64.57853, -64.51725, -64.45511, -64.39188, -64.3274, 
        -64.26093, -64.19173, -64.11884, -64.04208, -63.96141, -63.87763, 
        -63.79154, -63.70379, -63.61605, -63.52921, -63.44403, -63.36079, 
        -63.27887, -63.19806, -63.11756, -63.0371, -62.95653, -62.87577, 
        -62.79494, -62.71406, -62.63311, -62.55215, -62.4713, -62.3909, 
        -62.31041, -62.22884, -62.14741, -62.06444, -61.97982, -61.89376, 
        -61.80681, -61.71934, -61.63208, -61.54568, -61.46093, -61.37886, 
        -61.30051, -61.22661, -61.15774, -61.09393, -61.0348, -60.97978, 
        -60.92821, -60.87971, -60.83419, -60.7917, -60.75199, -60.71469, 
        -60.67902, -60.64524, -60.61367, -60.58451, -60.55788, -60.53388, 
        -60.51252, -60.4929, -60.47475, -60.4577, -60.4414, -60.42567, 
        -60.41097,
  -50.80431, -50.91506, -51.0246, -51.13708, -51.25344, -51.37632, 
        -51.50848, -51.65083, -51.80447, -51.96952, -52.14617, -52.33381, 
        -52.53139, -52.73743, -52.95021, -53.16784, -53.38855, -53.6109, 
        -53.83767, -54.06826, -54.3035, -54.54396, -54.79025, -55.04251, 
        -55.30093, -55.56575, -55.83603, -56.11073, -56.38928, -56.66999, 
        -56.95104, -57.22912, -57.50384, -57.77113, -58.02853, -58.27431, 
        -58.5072, -58.72673, -58.93364, -59.12904, -59.31418, -59.49073, 
        -59.66045, -59.82458, -59.98415, -60.13952, -60.29016, -60.43452, 
        -60.57392, -60.70704, -60.83436, -60.95621, -61.07365, -61.18709, 
        -61.2974, -61.40469, -61.50917, -61.61023, -61.70731, -61.7998, 
        -61.88811, -61.97257, -62.05392, -62.133, -62.21005, -62.28796, 
        -62.36622, -62.44509, -62.52452, -62.60436, -62.6843, -62.76398, 
        -62.8432, -62.92119, -62.99858, -63.07617, -63.15447, -63.2336, 
        -63.31384, -63.39434, -63.47508, -63.55474, -63.63503, -63.71523, 
        -63.79571, -63.87635, -63.95752, -64.03955, -64.12231, -64.20575, 
        -64.28989, -64.37449, -64.45915, -64.5434, -64.62701, -64.71017, 
        -64.79358, -64.87761, -64.96237, -65.04739, -65.13445, -65.22253, 
        -65.31148, -65.40063, -65.49005, -65.57921, -65.66785, -65.75522, 
        -65.84054, -65.92404, -66.00546, -66.08413, -66.16029, -66.23304, 
        -66.30273, -66.36944, -66.43354, -66.49532, -66.55434, -66.61043, 
        -66.66655, -66.72199, -66.77716, -66.83125, -66.88445, -66.936, 
        -66.98586, -67.03487, -67.08251, -67.12975, -67.17734, -67.22529, 
        -67.27442, -67.32401, -67.37362, -67.42319, -67.47205, -67.52058, 
        -67.56777, -67.61404, -67.65849, -67.70174, -67.74298, -67.78157, 
        -67.81783, -67.85211, -67.88488, -67.91679, -67.94743, -67.97697, 
        -68.00515, -68.03155, -68.05611, -68.07856, -68.09892, -68.11709, 
        -68.13293, -68.14616, -68.15575, -68.16206, -68.16449, -68.16311, 
        -68.15768, -68.14686, -68.13283, -68.1147, -68.09254, -68.06667, 
        -68.03642, -68.00372, -67.96962, -67.93511, -67.90057, -67.86506, 
        -67.82871, -67.79128, -67.7523, -67.71207, -67.6699, -67.62629, 
        -67.58041, -67.53246, -67.4822, -67.42904, -67.37313, -67.31446, 
        -67.25312, -67.18895, -67.12124, -67.05239, -66.98229, -66.91182, 
        -66.84133, -66.77116, -66.70203, -66.63402, -66.56735, -66.50216, 
        -66.43805, -66.37572, -66.31516, -66.25687, -66.20153, -66.14868, 
        -66.09834, -66.05043, -66.0049, -65.96155, -65.91977, -65.87894, 
        -65.83877, -65.79888, -65.75864, -65.71735, -65.67472, -65.63091, 
        -65.58586, -65.53839, -65.49036, -65.44072, -65.38976, -65.33798, 
        -65.2858, -65.23329, -65.1806, -65.12756, -65.07403, -65.02004, 
        -64.96538, -64.90993, -64.85365, -64.79653, -64.73875, -64.67999, 
        -64.62065, -64.56046, -64.49955, -64.43774, -64.37465, -64.31011, 
        -64.24332, -64.17357, -64.10032, -64.02287, -63.94142, -63.85675, 
        -63.76978, -63.68146, -63.59277, -63.50506, -63.41889, -63.33344, 
        -63.25039, -63.16795, -63.08596, -63.00406, -62.92223, -62.84042, 
        -62.75826, -62.67596, -62.59344, -62.51118, -62.42939, -62.34797, 
        -62.26694, -62.18589, -62.10426, -62.02144, -61.93695, -61.85112, 
        -61.76444, -61.67751, -61.59102, -61.50523, -61.4213, -61.34006, 
        -61.26269, -61.19011, -61.12266, -61.06064, -61.00365, -60.95096, 
        -60.90171, -60.8555, -60.81224, -60.77193, -60.73415, -60.69901, 
        -60.66499, -60.63287, -60.60246, -60.57374, -60.54742, -60.5235, 
        -60.50114, -60.48201, -60.46506, -60.44971, -60.43557, -60.42223, 
        -60.40974,
  -50.832, -50.95263, -51.07342, -51.19552, -51.32169, -51.45398, 
        -51.59504, -51.74633, -51.90797, -52.07987, -52.26162, -52.4518, 
        -52.65167, -52.85905, -53.07227, -53.29011, -53.51131, -53.73531, 
        -53.96314, -54.1953, -54.4326, -54.6758, -54.92514, -55.18071, 
        -55.44279, -55.71104, -55.98344, -56.26094, -56.54165, -56.82384, 
        -57.10529, -57.38362, -57.65623, -57.92022, -58.17327, -58.41416, 
        -58.64194, -58.85684, -59.05968, -59.25148, -59.43379, -59.60724, 
        -59.77539, -59.93847, -60.09702, -60.25161, -60.40174, -60.54605, 
        -60.68429, -60.8163, -60.94229, -61.06309, -61.1794, -61.29208, 
        -61.40191, -61.50886, -61.61274, -61.71346, -61.80874, -61.90073, 
        -61.98825, -62.07188, -62.15265, -62.2314, -62.30904, -62.38636, 
        -62.46442, -62.54292, -62.62186, -62.70128, -62.78049, -62.85957, 
        -62.93817, -63.01606, -63.09357, -63.1707, -63.25013, -63.33084, 
        -63.4127, -63.49514, -63.57732, -63.65925, -63.74085, -63.822, 
        -63.90358, -63.98568, -64.06881, -64.15305, -64.23784, -64.32339, 
        -64.40921, -64.49505, -64.58055, -64.66392, -64.74736, -64.82973, 
        -64.91209, -64.99494, -65.07841, -65.16328, -65.24955, -65.33735, 
        -65.42647, -65.51604, -65.60559, -65.69476, -65.78316, -65.87002, 
        -65.95489, -66.03783, -66.11873, -66.19736, -66.27232, -66.34545, 
        -66.41594, -66.48386, -66.54872, -66.61146, -66.67118, -66.72896, 
        -66.78537, -66.84132, -66.89721, -66.95207, -67.00564, -67.05793, 
        -67.1089, -67.15891, -67.20761, -67.25602, -67.30436, -67.35329, 
        -67.40178, -67.45159, -67.50183, -67.55166, -67.60138, -67.65036, 
        -67.69798, -67.74468, -67.7898, -67.83282, -67.87351, -67.91129, 
        -67.94682, -67.98045, -68.01293, -68.04453, -68.07438, -68.10297, 
        -68.13002, -68.15547, -68.1789, -68.19968, -68.21828, -68.23348, 
        -68.24711, -68.258, -68.26545, -68.26963, -68.27015, -68.26714, 
        -68.26044, -68.24926, -68.2339, -68.21428, -68.19054, -68.16277, 
        -68.13107, -68.0969, -68.06156, -68.02589, -67.99018, -67.9536, 
        -67.9162, -67.87769, -67.83772, -67.79643, -67.75328, -67.70729, 
        -67.65983, -67.61017, -67.55786, -67.50242, -67.44457, -67.38354, 
        -67.31967, -67.25282, -67.18336, -67.1116, -67.03848, -66.96488, 
        -66.8912, -66.81779, -66.74564, -66.67496, -66.60598, -66.53855, 
        -66.4723, -66.40742, -66.3441, -66.28268, -66.2234, -66.16611, 
        -66.1114, -66.05931, -66.00899, -65.96206, -65.91718, -65.87401, 
        -65.83199, -65.7905, -65.74893, -65.70629, -65.6624, -65.61674, 
        -65.56977, -65.5213, -65.47128, -65.42004, -65.36805, -65.31558, 
        -65.26308, -65.21027, -65.1572, -65.10334, -65.0488, -64.99353, 
        -64.93743, -64.88083, -64.82372, -64.76592, -64.70743, -64.64806, 
        -64.58834, -64.528, -64.46695, -64.40523, -64.34107, -64.27612, 
        -64.20888, -64.13831, -64.06425, -63.98587, -63.90371, -63.8182, 
        -63.73043, -63.64123, -63.55173, -63.4632, -63.37604, -63.29041, 
        -63.20588, -63.12173, -63.03815, -62.95466, -62.87144, -62.78834, 
        -62.70497, -62.62149, -62.53796, -62.45466, -62.37191, -62.28961, 
        -62.20778, -62.12605, -62.04386, -61.96082, -61.87636, -61.79097, 
        -61.70501, -61.6191, -61.53385, -61.44971, -61.36742, -61.28796, 
        -61.21244, -61.14075, -61.07533, -61.01547, -60.96079, -60.91056, 
        -60.86403, -60.82048, -60.77986, -60.74176, -60.70641, -60.67334, 
        -60.64144, -60.611, -60.58176, -60.55381, -60.52746, -60.50305, 
        -60.48117, -60.46213, -60.44571, -60.43161, -60.419, -60.40757, 
        -60.39702,
  -50.83028, -50.96061, -51.09079, -51.22245, -51.35743, -51.49773, 
        -51.6471, -51.80615, -51.97469, -52.15285, -52.33948, -52.53402, 
        -52.73629, -52.94518, -53.15959, -53.3784, -53.60115, -53.82729, 
        -54.05744, -54.29277, -54.53259, -54.77984, -55.03356, -55.2937, 
        -55.56016, -55.83247, -56.10949, -56.39003, -56.6728, -56.95592, 
        -57.2372, -57.51395, -57.78364, -58.04365, -58.29214, -58.52776, 
        -58.74936, -58.9595, -59.1579, -59.34614, -59.52557, -59.69773, 
        -59.86404, -60.02567, -60.18326, -60.3368, -60.48584, -60.62903, 
        -60.76633, -60.89735, -61.02246, -61.14252, -61.25724, -61.36963, 
        -61.47927, -61.58627, -61.69013, -61.79035, -61.8863, -61.97763, 
        -62.06475, -62.14812, -62.22843, -62.30695, -62.38441, -62.46153, 
        -62.53919, -62.61722, -62.69569, -62.77327, -62.85168, -62.92979, 
        -63.00733, -63.08478, -63.16234, -63.24091, -63.3213, -63.40338, 
        -63.48676, -63.57103, -63.65516, -63.73849, -63.82119, -63.90405, 
        -63.98751, -64.07169, -64.15585, -64.24202, -64.32919, -64.41694, 
        -64.50504, -64.59251, -64.67889, -64.76395, -64.8476, -64.93007, 
        -65.01176, -65.09367, -65.17637, -65.26048, -65.34615, -65.43336, 
        -65.52193, -65.61155, -65.70147, -65.78977, -65.87784, -65.96413, 
        -66.04843, -66.13074, -66.2112, -66.28926, -66.3651, -66.43849, 
        -66.50984, -66.5784, -66.64442, -66.7076, -66.76841, -66.82698, 
        -66.8845, -66.94123, -66.99704, -67.05284, -67.10769, -67.16032, 
        -67.21259, -67.26353, -67.314, -67.36383, -67.41358, -67.46362, 
        -67.51377, -67.56412, -67.61452, -67.66498, -67.715, -67.76418, 
        -67.81251, -67.85954, -67.90481, -67.94772, -67.98776, -68.02547, 
        -68.06094, -68.09489, -68.12606, -68.1565, -68.18589, -68.21363, 
        -68.23969, -68.26374, -68.28522, -68.30443, -68.32093, -68.33515, 
        -68.34633, -68.35455, -68.35976, -68.36166, -68.36053, -68.35579, 
        -68.34718, -68.33481, -68.31823, -68.29769, -68.27264, -68.24321, 
        -68.21046, -68.17522, -68.13784, -68.10094, -68.06358, -68.02573, 
        -67.98705, -67.94745, -67.9066, -67.86439, -67.82054, -67.7747, 
        -67.72662, -67.67582, -67.6218, -67.56478, -67.50493, -67.44157, 
        -67.37489, -67.30556, -67.23354, -67.15934, -67.08392, -67.00776, 
        -66.93144, -66.85586, -66.7816, -66.70909, -66.63727, -66.56798, 
        -66.49996, -66.43276, -66.36674, -66.30183, -66.23833, -66.17697, 
        -66.11777, -66.06103, -66.00723, -65.95607, -65.90739, -65.86084, 
        -65.81593, -65.77197, -65.72805, -65.68343, -65.63741, -65.58981, 
        -65.54055, -65.48971, -65.43793, -65.38513, -65.33199, -65.27898, 
        -65.22601, -65.17301, -65.1196, -65.06532, -65.00901, -64.95264, 
        -64.89556, -64.83762, -64.77934, -64.72069, -64.66143, -64.60178, 
        -64.54155, -64.48089, -64.41946, -64.35721, -64.29363, -64.228, 
        -64.15951, -64.08791, -64.01252, -63.93307, -63.84983, -63.76338, 
        -63.67467, -63.58466, -63.49432, -63.4048, -63.31651, -63.22939, 
        -63.143, -63.0573, -62.97186, -62.88701, -62.80249, -62.71785, 
        -62.63367, -62.54943, -62.46532, -62.38139, -62.29692, -62.21398, 
        -62.13129, -62.04883, -61.96604, -61.88254, -61.79837, -61.71352, 
        -61.62872, -61.54436, -61.46087, -61.37887, -61.29896, -61.2221, 
        -61.14914, -61.08083, -61.0179, -60.96052, -60.9085, -60.86107, 
        -60.8173, -60.77672, -60.73905, -60.70388, -60.67106, -60.64029, 
        -60.6106, -60.58198, -60.55386, -60.5265, -60.50012, -60.47528, 
        -60.45308, -60.43356, -60.41736, -60.40394, -60.39236, -60.38235, 
        -60.37344,
  -50.7973, -50.93651, -51.07555, -51.2159, -51.35939, -51.50882, 
        -51.66579, -51.83162, -52.00648, -52.18992, -52.38112, -52.57914, 
        -52.78389, -52.99455, -53.21072, -53.43065, -53.65578, -53.88502, 
        -54.11913, -54.35879, -54.6044, -54.85671, -55.11578, -55.3812, 
        -55.65265, -55.9293, -56.2101, -56.49376, -56.7784, -57.06235, 
        -57.3419, -57.61674, -57.88317, -58.13901, -58.38271, -58.61323, 
        -58.83084, -59.03622, -59.23022, -59.41484, -59.5914, -59.7613, 
        -59.9259, -60.0861, -60.24239, -60.39457, -60.54102, -60.68309, 
        -60.81923, -60.94947, -61.07384, -61.19338, -61.30891, -61.42125, 
        -61.53104, -61.6382, -61.74205, -61.84209, -61.93782, -62.02898, 
        -62.11598, -62.19923, -62.27868, -62.35726, -62.43477, -62.51192, 
        -62.58918, -62.66681, -62.74457, -62.82207, -62.89948, -62.97622, 
        -63.05285, -63.12979, -63.20723, -63.28619, -63.36727, -63.45069, 
        -63.53576, -63.62181, -63.70676, -63.79193, -63.87657, -63.96139, 
        -64.04663, -64.13291, -64.2202, -64.30891, -64.39857, -64.48876, 
        -64.57912, -64.6684, -64.75615, -64.84241, -64.92699, -65.00993, 
        -65.0918, -65.17326, -65.25453, -65.33768, -65.42269, -65.50935, 
        -65.59757, -65.68694, -65.7765, -65.86562, -65.95352, -66.03916, 
        -66.12286, -66.20441, -66.28445, -66.36217, -66.43789, -66.51172, 
        -66.58374, -66.65327, -66.72006, -66.78407, -66.84455, -66.90404, 
        -66.96212, -67.01949, -67.07655, -67.1333, -67.18921, -67.2441, 
        -67.29775, -67.35034, -67.40271, -67.45424, -67.50541, -67.55652, 
        -67.60744, -67.65882, -67.71008, -67.7611, -67.8114, -67.86115, 
        -67.9102, -67.95648, -68.00204, -68.04491, -68.08518, -68.12319, 
        -68.15916, -68.19324, -68.22527, -68.25555, -68.28417, -68.31077, 
        -68.33537, -68.35754, -68.37714, -68.39431, -68.40871, -68.42041, 
        -68.4292, -68.43485, -68.43789, -68.43772, -68.43442, -68.42638, 
        -68.41602, -68.40235, -68.38458, -68.36279, -68.33674, -68.30665, 
        -68.27316, -68.23737, -68.20031, -68.16245, -68.12397, -68.08495, 
        -68.04506, -68.00429, -67.96233, -67.91892, -67.87437, -67.82808, 
        -67.7793, -67.72755, -67.67259, -67.61455, -67.55299, -67.48788, 
        -67.41781, -67.34587, -67.27152, -67.1951, -67.11774, -67.0396, 
        -66.96145, -66.88421, -66.80861, -66.73499, -66.66307, -66.59261, 
        -66.52323, -66.45411, -66.38517, -66.3168, -66.24973, -66.18417, 
        -66.12064, -66.05923, -66.00033, -65.94402, -65.89072, -65.84001, 
        -65.79134, -65.74358, -65.69621, -65.64843, -65.59937, -65.5477, 
        -65.49574, -65.44252, -65.38902, -65.33494, -65.28088, -65.22713, 
        -65.17381, -65.12047, -65.06666, -65.01202, -64.95626, -64.89913, 
        -64.84109, -64.78226, -64.723, -64.66337, -64.60338, -64.54338, 
        -64.48261, -64.42134, -64.35919, -64.29614, -64.23144, -64.16454, 
        -64.09459, -64.02108, -63.94386, -63.86291, -63.7785, -63.69088, 
        -63.60114, -63.51005, -63.41743, -63.32658, -63.23682, -63.14801, 
        -63.05993, -62.97261, -62.88569, -62.79925, -62.71338, -62.62808, 
        -62.54324, -62.45874, -62.37446, -62.29029, -62.20652, -62.12323, 
        -62.04018, -61.95721, -61.87383, -61.79031, -61.70651, -61.62265, 
        -61.53925, -61.45668, -61.37546, -61.29608, -61.21902, -61.14503, 
        -61.07489, -61.00956, -60.94942, -60.89484, -60.84564, -60.80108, 
        -60.76043, -60.72305, -60.68853, -60.65654, -60.62667, -60.59844, 
        -60.57125, -60.5443, -60.51657, -60.4899, -60.46365, -60.43867, 
        -60.41586, -60.39645, -60.38027, -60.36705, -60.35612, -60.34704, 
        -60.33945,
  -50.7348, -50.88265, -51.02964, -51.1777, -51.32924, -51.48602, 
        -51.65006, -51.82223, -52.0028, -52.19109, -52.38578, -52.58723, 
        -52.79457, -53.00752, -53.22607, -53.44955, -53.67794, -53.91122, 
        -54.15007, -54.39483, -54.64599, -54.90419, -55.1692, -55.4403, 
        -55.71706, -55.99744, -56.28219, -56.56902, -56.85568, -57.14009, 
        -57.41991, -57.69271, -57.95595, -58.20774, -58.44702, -58.6726, 
        -58.88525, -59.08598, -59.27596, -59.45706, -59.62978, -59.79749, 
        -59.96022, -60.11886, -60.27363, -60.42433, -60.57023, -60.71091, 
        -60.84586, -60.97504, -61.09889, -61.21814, -61.33363, -61.44609, 
        -61.55599, -61.6633, -61.76623, -61.86635, -61.96191, -62.05291, 
        -62.13987, -62.22348, -62.30429, -62.38319, -62.46103, -62.53857, 
        -62.61597, -62.6933, -62.77053, -62.847, -62.92311, -62.99879, 
        -63.07451, -63.14993, -63.22722, -63.30667, -63.38866, -63.47307, 
        -63.55957, -63.64719, -63.73497, -63.82212, -63.90894, -63.99549, 
        -64.0828, -64.17155, -64.26167, -64.35272, -64.44492, -64.53747, 
        -64.62994, -64.7204, -64.81023, -64.89809, -64.98386, -65.06796, 
        -65.15059, -65.2322, -65.31403, -65.39671, -65.48094, -65.56715, 
        -65.65472, -65.74364, -65.83264, -65.92111, -66.00839, -66.09377, 
        -66.17677, -66.25797, -66.33749, -66.41439, -66.49035, -66.56472, 
        -66.63741, -66.7076, -66.77515, -66.83985, -66.90203, -66.9621, 
        -67.02099, -67.07914, -67.13677, -67.19406, -67.25063, -67.30675, 
        -67.36206, -67.41642, -67.47031, -67.52365, -67.57671, -67.62861, 
        -67.68114, -67.73333, -67.7856, -67.83739, -67.88844, -67.93861, 
        -67.98824, -68.03587, -68.0817, -68.12537, -68.16653, -68.20525, 
        -68.24176, -68.27624, -68.30878, -68.33892, -68.36678, -68.39209, 
        -68.41504, -68.43513, -68.45261, -68.46666, -68.47882, -68.48826, 
        -68.4947, -68.49812, -68.4987, -68.49619, -68.49063, -68.48167, 
        -68.46927, -68.45367, -68.43449, -68.41162, -68.38486, -68.35417, 
        -68.3204, -68.28411, -68.2468, -68.20869, -68.16977, -68.12981, 
        -68.0889, -68.04723, -68.00441, -67.95932, -67.91383, -67.86655, 
        -67.8169, -67.7646, -67.70911, -67.65015, -67.58737, -67.5209, 
        -67.45079, -67.3773, -67.30103, -67.22253, -67.14302, -67.06316, 
        -66.98383, -66.90569, -66.8293, -66.75478, -66.68226, -66.6109, 
        -66.54022, -66.46919, -66.39829, -66.32745, -66.25687, -66.18739, 
        -66.11823, -66.05197, -65.9882, -65.92693, -65.86834, -65.81224, 
        -65.75817, -65.7057, -65.65367, -65.60097, -65.54776, -65.4935, 
        -65.43834, -65.38247, -65.32681, -65.27122, -65.21649, -65.16231, 
        -65.1084, -65.05467, -65.0004, -64.94525, -64.88886, -64.83123, 
        -64.77245, -64.71292, -64.65299, -64.59266, -64.53203, -64.47123, 
        -64.40998, -64.3471, -64.2842, -64.21983, -64.15366, -64.08487, 
        -64.01292, -63.93729, -63.85789, -63.77475, -63.68804, -63.59893, 
        -63.50776, -63.41512, -63.32212, -63.22974, -63.13823, -63.04771, 
        -62.95782, -62.8688, -62.78035, -62.69283, -62.6063, -62.52057, 
        -62.43577, -62.35138, -62.26748, -62.1838, -62.10026, -62.01694, 
        -61.93369, -61.85059, -61.7675, -61.68415, -61.60108, -61.51849, 
        -61.43687, -61.35647, -61.27772, -61.20108, -61.12602, -61.05527, 
        -60.98836, -60.92596, -60.86884, -60.81709, -60.77068, -60.72909, 
        -60.6915, -60.65733, -60.62612, -60.59748, -60.57085, -60.54545, 
        -60.52075, -60.49596, -60.47069, -60.44503, -60.41916, -60.39433, 
        -60.37154, -60.35191, -60.33571, -60.32258, -60.31194, -60.30325, 
        -60.29638,
  -50.64224, -50.79809, -50.95263, -51.10806, -51.26575, -51.42949, 
        -51.60006, -51.77826, -51.96415, -52.15723, -52.35674, -52.56213, 
        -52.77245, -52.98812, -53.20946, -53.4362, -53.66841, -53.90613, 
        -54.15002, -54.39951, -54.65664, -54.92092, -55.19197, -55.46894, 
        -55.75116, -56.03749, -56.32656, -56.6164, -56.90513, -57.19042, 
        -57.46946, -57.74027, -58.00065, -58.24882, -58.48383, -58.70425, 
        -58.91249, -59.10883, -59.29491, -59.47256, -59.64359, -59.80923, 
        -59.97014, -60.12737, -60.28046, -60.42949, -60.57374, -60.71277, 
        -60.84638, -60.97457, -61.09781, -61.2158, -61.33121, -61.44379, 
        -61.55368, -61.66101, -61.76498, -61.86479, -61.96027, -62.05119, 
        -62.13832, -62.22232, -62.30375, -62.38342, -62.46207, -62.54028, 
        -62.61816, -62.69433, -62.77108, -62.84693, -62.92224, -62.99712, 
        -63.07227, -63.1483, -63.22578, -63.30562, -63.38861, -63.47412, 
        -63.56179, -63.6506, -63.74005, -63.82927, -63.91795, -64.00689, 
        -64.0967, -64.18689, -64.27965, -64.37339, -64.46812, -64.56312, 
        -64.65791, -64.75179, -64.84357, -64.93318, -65.02045, -65.10596, 
        -65.18974, -65.27202, -65.35379, -65.43637, -65.52024, -65.60547, 
        -65.69195, -65.77982, -65.86699, -65.95473, -66.04134, -66.1263, 
        -66.20943, -66.29063, -66.37056, -66.44911, -66.52594, -66.6009, 
        -66.67388, -66.74465, -66.81271, -66.87749, -66.93987, -67.00031, 
        -67.05949, -67.11818, -67.17585, -67.23244, -67.2896, -67.34658, 
        -67.40342, -67.45952, -67.51537, -67.57088, -67.62617, -67.68113, 
        -67.73518, -67.78864, -67.8415, -67.89429, -67.94621, -67.99724, 
        -68.04694, -68.09531, -68.1423, -68.18729, -68.22926, -68.26888, 
        -68.30633, -68.34052, -68.37347, -68.40327, -68.43043, -68.45438, 
        -68.47569, -68.49438, -68.50994, -68.52271, -68.53279, -68.53994, 
        -68.54433, -68.54535, -68.5437, -68.53918, -68.53139, -68.52059, 
        -68.50626, -68.48858, -68.46775, -68.44388, -68.41632, -68.38489, 
        -68.34978, -68.3134, -68.27614, -68.23811, -68.19881, -68.15842, 
        -68.11701, -68.07475, -68.03157, -67.9866, -67.94028, -67.89215, 
        -67.84184, -67.78886, -67.73251, -67.67303, -67.60979, -67.5429, 
        -67.47231, -67.39783, -67.32052, -67.24088, -67.15988, -67.07877, 
        -66.9983, -66.91941, -66.84126, -66.76637, -66.69331, -66.6209, 
        -66.549, -66.47712, -66.40469, -66.33187, -66.25867, -66.18567, 
        -66.1133, -66.04219, -65.97331, -65.90678, -65.84254, -65.7807, 
        -65.72076, -65.66213, -65.60405, -65.54575, -65.48692, -65.42783, 
        -65.36838, -65.30977, -65.2516, -65.19444, -65.13837, -65.0833, 
        -65.02863, -64.97416, -64.91832, -64.8626, -64.80578, -64.74747, 
        -64.68803, -64.62784, -64.5672, -64.5064, -64.44522, -64.38379, 
        -64.32201, -64.25937, -64.1955, -64.12965, -64.06144, -63.9903, 
        -63.91584, -63.83739, -63.75504, -63.66917, -63.58018, -63.4887, 
        -63.39548, -63.30112, -63.20651, -63.11216, -63.01881, -62.92646, 
        -62.83495, -62.74435, -62.65483, -62.5666, -62.47988, -62.39447, 
        -62.3102, -62.22572, -62.14291, -62.06017, -61.97743, -61.89473, 
        -61.812, -61.72931, -61.64677, -61.56438, -61.48249, -61.40138, 
        -61.3217, -61.24355, -61.16728, -61.09338, -61.02239, -60.95477, 
        -60.89114, -60.83206, -60.77786, -60.72885, -60.68533, -60.64658, 
        -60.61187, -60.5808, -60.55292, -60.52771, -60.5045, -60.48229, 
        -60.46031, -60.43783, -60.41441, -60.38999, -60.36485, -60.34035, 
        -60.31785, -60.29829, -60.28205, -60.26878, -60.25827, -60.25002, 
        -60.24398,
  -50.52039, -50.68335, -50.84515, -51.00729, -51.17244, -51.34288, 
        -51.51961, -51.70356, -51.89466, -52.09238, -52.29597, -52.50515, 
        -52.71915, -52.93808, -53.16159, -53.39191, -53.62816, -53.87086, 
        -54.11998, -54.37631, -54.63931, -54.90966, -55.18669, -55.46956, 
        -55.75744, -56.04891, -56.34228, -56.63535, -56.92613, -57.21118, 
        -57.48979, -57.75898, -58.01708, -58.26205, -58.49352, -58.71116, 
        -58.91558, -59.10811, -59.29069, -59.46526, -59.63349, -59.79686, 
        -59.95617, -60.11175, -60.26336, -60.40963, -60.55231, -60.68976, 
        -60.82201, -60.94905, -61.07133, -61.18972, -61.3047, -61.41699, 
        -61.52672, -61.63372, -61.73739, -61.83691, -61.9321, -62.02306, 
        -62.1102, -62.19367, -62.27602, -62.35695, -62.43685, -62.51586, 
        -62.59422, -62.67173, -62.74819, -62.82385, -62.89878, -62.97333, 
        -63.04839, -63.12463, -63.20269, -63.28353, -63.36714, -63.45355, 
        -63.5422, -63.63132, -63.72225, -63.81318, -63.90419, -63.99556, 
        -64.08789, -64.18179, -64.27721, -64.37367, -64.4711, -64.56887, 
        -64.66608, -64.76195, -64.85584, -64.94756, -65.03673, -65.12353, 
        -65.20849, -65.29086, -65.37322, -65.45532, -65.53832, -65.62261, 
        -65.70818, -65.79476, -65.88184, -65.96886, -66.05494, -66.13999, 
        -66.22337, -66.30553, -66.38617, -66.46539, -66.54305, -66.6188, 
        -66.69228, -66.76302, -66.82961, -66.89429, -66.95644, -67.01687, 
        -67.07597, -67.13421, -67.19196, -67.24976, -67.30759, -67.36539, 
        -67.42361, -67.48177, -67.53979, -67.59801, -67.65558, -67.71243, 
        -67.76812, -67.82286, -67.87705, -67.93044, -67.98305, -68.03391, 
        -68.08493, -68.13476, -68.18274, -68.22849, -68.27158, -68.31264, 
        -68.35143, -68.38719, -68.42009, -68.44957, -68.47583, -68.49892, 
        -68.51885, -68.53605, -68.54993, -68.56079, -68.56898, -68.57392, 
        -68.57607, -68.57514, -68.57148, -68.56488, -68.55421, -68.54131, 
        -68.5251, -68.50577, -68.48344, -68.45808, -68.4295, -68.39765, 
        -68.36354, -68.32738, -68.28982, -68.25172, -68.2125, -68.17233, 
        -68.13119, -68.08875, -68.04497, -67.9995, -67.95238, -67.90365, 
        -67.85258, -67.79901, -67.74233, -67.6824, -67.61809, -67.55091, 
        -67.48014, -67.40582, -67.32835, -67.24853, -67.1671, -67.08549, 
        -67.00442, -66.92481, -66.84708, -66.77152, -66.69749, -66.62408, 
        -66.55141, -66.47865, -66.40521, -66.33107, -66.25589, -66.18022, 
        -66.10445, -66.02924, -65.9552, -65.88293, -65.81272, -65.74465, 
        -65.6782, -65.61282, -65.54688, -65.48177, -65.41646, -65.35152, 
        -65.28753, -65.225, -65.16387, -65.10469, -65.04681, -64.99007, 
        -64.93401, -64.87824, -64.82234, -64.76585, -64.70831, -64.64944, 
        -64.58929, -64.52831, -64.46677, -64.40522, -64.34362, -64.28184, 
        -64.21951, -64.15601, -64.0908, -64.02317, -63.95266, -63.87882, 
        -63.80116, -63.71943, -63.6338, -63.54464, -63.45269, -63.35735, 
        -63.26166, -63.16537, -63.06874, -62.97262, -62.87719, -62.78302, 
        -62.69013, -62.59844, -62.50825, -62.41981, -62.33334, -62.24862, 
        -62.16574, -62.08393, -62.0027, -61.92175, -61.84051, -61.75912, 
        -61.67766, -61.59604, -61.51461, -61.43353, -61.3532, -61.27406, 
        -61.19628, -61.12017, -61.04632, -60.97511, -60.90712, -60.84272, 
        -60.7824, -60.72652, -60.67547, -60.62951, -60.58852, -60.55231, 
        -60.52023, -60.49208, -60.46745, -60.4457, -60.42595, -60.40606, 
        -60.38706, -60.36699, -60.34541, -60.32235, -60.29829, -60.27443, 
        -60.25237, -60.23299, -60.21663, -60.20321, -60.19268, -60.18495, 
        -60.17991,
  -50.37358, -50.54274, -50.711, -50.87942, -51.05056, -51.22709, 
        -51.40973, -51.59924, -51.79546, -51.99697, -52.20507, -52.41814, 
        -52.63643, -52.85924, -53.08741, -53.32162, -53.56248, -53.81015, 
        -54.06447, -54.32638, -54.5954, -54.87176, -55.15482, -55.44361, 
        -55.73615, -56.03247, -56.32975, -56.62576, -56.91853, -57.20557, 
        -57.48413, -57.75225, -58.00831, -58.25086, -58.4794, -58.69405, 
        -58.89545, -59.08488, -59.26451, -59.43523, -59.60101, -59.76225, 
        -59.91964, -60.07335, -60.2233, -60.36893, -60.50985, -60.64578, 
        -60.77662, -60.90244, -61.02365, -61.14098, -61.25521, -61.3667, 
        -61.47571, -61.581, -61.68394, -61.78315, -61.87798, -61.96888, 
        -62.05619, -62.14099, -62.22422, -62.30626, -62.3871, -62.46722, 
        -62.54637, -62.62441, -62.70113, -62.77684, -62.85185, -62.9268, 
        -63.00156, -63.07864, -63.15779, -63.23942, -63.32397, -63.41126, 
        -63.50076, -63.59212, -63.68456, -63.7775, -63.87083, -63.96454, 
        -64.05946, -64.15585, -64.25423, -64.35385, -64.45409, -64.55471, 
        -64.6534, -64.75173, -64.84805, -64.94168, -65.03252, -65.12097, 
        -65.20715, -65.29124, -65.3738, -65.45549, -65.53787, -65.62097, 
        -65.70554, -65.79111, -65.87704, -65.96331, -66.0494, -66.13471, 
        -66.21887, -66.30095, -66.38261, -66.46287, -66.5415, -66.61752, 
        -66.69078, -66.76086, -66.82797, -66.89201, -66.95351, -67.01339, 
        -67.07177, -67.12974, -67.18744, -67.24535, -67.30349, -67.36235, 
        -67.42197, -67.48223, -67.54249, -67.60185, -67.66157, -67.72061, 
        -67.77846, -67.83474, -67.88997, -67.94459, -67.99868, -68.05231, 
        -68.10479, -68.15566, -68.20467, -68.25188, -68.29665, -68.33874, 
        -68.37817, -68.41433, -68.44708, -68.47639, -68.50198, -68.52422, 
        -68.54302, -68.55785, -68.57054, -68.57972, -68.58591, -68.58896, 
        -68.58923, -68.58648, -68.58063, -68.57193, -68.56018, -68.54572, 
        -68.52812, -68.50721, -68.48329, -68.45644, -68.42706, -68.39509, 
        -68.36086, -68.32474, -68.28731, -68.24925, -68.21024, -68.17038, 
        -68.12929, -68.08601, -68.04238, -67.99713, -67.94986, -67.90044, 
        -67.84843, -67.79411, -67.7374, -67.67751, -67.6143, -67.54709, 
        -67.47667, -67.40302, -67.32599, -67.24673, -67.16596, -67.08473, 
        -67.00394, -66.92429, -66.84644, -66.76994, -66.69462, -66.6203, 
        -66.54643, -66.47267, -66.39819, -66.3227, -66.24497, -66.16705, 
        -66.08844, -66.00976, -65.93158, -65.85426, -65.77825, -65.70373, 
        -65.63032, -65.55762, -65.48531, -65.41299, -65.34081, -65.2695, 
        -65.19997, -65.13261, -65.06767, -65.00526, -64.94472, -64.88564, 
        -64.82747, -64.76965, -64.71195, -64.65394, -64.59507, -64.53509, 
        -64.47405, -64.41201, -64.34949, -64.28721, -64.22515, -64.1618, 
        -64.09896, -64.03445, -63.96775, -63.89793, -63.82476, -63.7477, 
        -63.66646, -63.58105, -63.49171, -63.39902, -63.30373, -63.20652, 
        -63.10849, -63.00995, -62.91151, -62.81323, -62.71622, -62.62054, 
        -62.5265, -62.43396, -62.34337, -62.25508, -62.16933, -62.08611, 
        -62.00484, -61.92516, -61.84638, -61.76778, -61.68907, -61.60986, 
        -61.53019, -61.45034, -61.37054, -61.29122, -61.21259, -61.13521, 
        -61.05944, -60.98477, -60.91355, -60.84507, -60.78008, -60.71885, 
        -60.66186, -60.60931, -60.56141, -60.5182, -60.47967, -60.44577, 
        -60.41624, -60.39088, -60.36917, -60.35049, -60.33381, -60.31778, 
        -60.30156, -60.28386, -60.26408, -60.24247, -60.21975, -60.19688, 
        -60.17525, -60.15604, -60.13969, -60.12628, -60.11589, -60.10882, 
        -60.1049,
  -50.20399, -50.37875, -50.5527, -50.72615, -50.90302, -51.08497, 
        -51.27331, -51.46805, -51.66927, -51.87654, -52.0893, -52.30681, 
        -52.52918, -52.7566, -52.98896, -53.22765, -53.4734, -53.72576, 
        -53.98445, -54.25179, -54.5267, -54.80896, -55.09803, -55.39249, 
        -55.69117, -55.99201, -56.29281, -56.59159, -56.88602, -57.17406, 
        -57.45298, -57.72054, -57.97521, -58.21511, -58.4416, -58.65392, 
        -58.85314, -59.0404, -59.21772, -59.38711, -59.55071, -59.70963, 
        -59.86483, -60.01646, -60.16447, -60.30823, -60.44755, -60.58196, 
        -60.71149, -60.83506, -60.95503, -61.07109, -61.18406, -61.29419, 
        -61.40178, -61.50665, -61.60853, -61.70682, -61.80109, -61.8917, 
        -61.9791, -62.06423, -62.14814, -62.23095, -62.31268, -62.3937, 
        -62.47272, -62.55146, -62.62871, -62.70525, -62.78127, -62.85733, 
        -62.93453, -63.01293, -63.09327, -63.17599, -63.26159, -63.34977, 
        -63.44023, -63.53268, -63.62671, -63.72148, -63.81705, -63.91328, 
        -64.00981, -64.10931, -64.21078, -64.31368, -64.41696, -64.52048, 
        -64.62326, -64.72432, -64.82298, -64.91888, -65.01147, -65.10149, 
        -65.18851, -65.27327, -65.35571, -65.43725, -65.51893, -65.60116, 
        -65.68327, -65.76743, -65.85255, -65.93829, -66.02422, -66.1102, 
        -66.19528, -66.27926, -66.36234, -66.44344, -66.52256, -66.59842, 
        -66.67124, -66.74073, -66.80682, -66.86972, -66.93011, -66.98877, 
        -67.04663, -67.10387, -67.16032, -67.21782, -67.27646, -67.33617, 
        -67.39711, -67.459, -67.52117, -67.58352, -67.6456, -67.70673, 
        -67.76657, -67.82476, -67.88197, -67.9389, -67.99503, -68.05048, 
        -68.10433, -68.15675, -68.20763, -68.25635, -68.30241, -68.34399, 
        -68.38378, -68.42033, -68.45316, -68.48227, -68.50727, -68.52876, 
        -68.54671, -68.56147, -68.57291, -68.58072, -68.58549, -68.58716, 
        -68.58572, -68.58123, -68.57335, -68.56259, -68.54916, -68.53299, 
        -68.51395, -68.49155, -68.46648, -68.4389, -68.40786, -68.37572, 
        -68.34115, -68.30509, -68.26828, -68.23029, -68.19144, -68.15141, 
        -68.11067, -68.06886, -68.02542, -67.98024, -67.93262, -67.8828, 
        -67.83062, -67.7761, -67.71908, -67.6589, -67.59591, -67.52982, 
        -67.46009, -67.38736, -67.31144, -67.23333, -67.15385, -67.07375, 
        -66.99305, -66.91392, -66.83572, -66.75867, -66.68272, -66.60755, 
        -66.5326, -66.45763, -66.38168, -66.30492, -66.22682, -66.14686, 
        -66.06609, -65.98444, -65.90264, -65.82102, -65.73972, -65.65889, 
        -65.57876, -65.49883, -65.41895, -65.33894, -65.2593, -65.1816, 
        -65.10581, -65.03282, -64.96298, -64.89626, -64.83211, -64.76874, 
        -64.70767, -64.64688, -64.58659, -64.52611, -64.46491, -64.40315, 
        -64.34033, -64.27708, -64.21355, -64.15033, -64.08755, -64.02448, 
        -63.96052, -63.89486, -63.82624, -63.75407, -63.67783, -63.59731, 
        -63.51254, -63.42312, -63.33014, -63.23356, -63.13497, -63.03495, 
        -62.93434, -62.83366, -62.73326, -62.63363, -62.53537, -62.43861, 
        -62.34373, -62.25065, -62.16016, -62.07249, -61.98694, -61.90528, 
        -61.82608, -61.74896, -61.67315, -61.59781, -61.52225, -61.44592, 
        -61.36908, -61.29166, -61.21405, -61.13673, -61.05992, -60.98446, 
        -60.91094, -60.8398, -60.77138, -60.70591, -60.64406, -60.58609, 
        -60.53248, -60.48322, -60.43826, -60.39779, -60.36176, -60.33012, 
        -60.30286, -60.27984, -60.26064, -60.2446, -60.23027, -60.2165, 
        -60.20195, -60.18605, -60.16822, -60.14805, -60.12642, -60.10443, 
        -60.08347, -60.0647, -60.04855, -60.03541, -60.02567, -60.01962, 
        -60.01734,
  -50.01351, -50.19386, -50.37297, -50.55284, -50.73529, -50.92214, 
        -51.11549, -51.3154, -51.52139, -51.73355, -51.95098, -52.17316, 
        -52.39997, -52.6312, -52.86872, -53.11208, -53.36251, -53.62025, 
        -53.88519, -54.1578, -54.4381, -54.72594, -55.02035, -55.3201, 
        -55.62358, -55.92846, -56.23248, -56.53361, -56.82871, -57.1179, 
        -57.39742, -57.66491, -57.91903, -58.15887, -58.38402, -58.59496, 
        -58.79261, -58.97829, -59.15393, -59.32163, -59.48319, -59.64001, 
        -59.793, -59.94252, -60.08749, -60.22928, -60.36687, -60.49982, 
        -60.62792, -60.75117, -60.86981, -60.98449, -61.0956, -61.20373, 
        -61.30937, -61.41225, -61.51233, -61.6091, -61.70247, -61.79234, 
        -61.87822, -61.96336, -62.04753, -62.13091, -62.21354, -62.29497, 
        -62.37563, -62.45525, -62.53368, -62.61161, -62.68932, -62.76738, 
        -62.84636, -62.92656, -63.00847, -63.09239, -63.17882, -63.26709, 
        -63.35866, -63.45236, -63.54778, -63.6445, -63.74232, -63.84128, 
        -63.94191, -64.04449, -64.14952, -64.2558, -64.36263, -64.46938, 
        -64.57515, -64.67915, -64.78053, -64.87883, -64.97353, -65.0647, 
        -65.15147, -65.23694, -65.32015, -65.40158, -65.48212, -65.563, 
        -65.64481, -65.72758, -65.81158, -65.89667, -65.98267, -66.06919, 
        -66.15533, -66.24062, -66.32446, -66.40627, -66.48564, -66.56114, 
        -66.63316, -66.70025, -66.76488, -66.82639, -66.88542, -66.94305, 
        -66.99978, -67.05629, -67.11315, -67.17067, -67.22945, -67.28941, 
        -67.3511, -67.41406, -67.47762, -67.54171, -67.60564, -67.66899, 
        -67.73105, -67.79197, -67.85219, -67.91161, -67.96893, -68.02638, 
        -68.08246, -68.13692, -68.18926, -68.23911, -68.28601, -68.32975, 
        -68.37041, -68.4072, -68.44022, -68.46906, -68.49356, -68.51427, 
        -68.53142, -68.54533, -68.55573, -68.56275, -68.5664, -68.56668, 
        -68.5639, -68.55786, -68.54754, -68.53533, -68.51999, -68.50201, 
        -68.4812, -68.45769, -68.43159, -68.40313, -68.37286, -68.34061, 
        -68.30642, -68.27052, -68.2334, -68.19555, -68.15715, -68.11754, 
        -68.07681, -68.03488, -67.99145, -67.94621, -67.89869, -67.84881, 
        -67.79646, -67.74199, -67.68518, -67.62452, -67.56216, -67.49665, 
        -67.42823, -67.35693, -67.2828, -67.20665, -67.12871, -67.04998, 
        -66.97131, -66.89297, -66.81518, -66.73799, -66.66156, -66.58528, 
        -66.50922, -66.43314, -66.35618, -66.27814, -66.19846, -66.11697, 
        -66.034, -65.95007, -65.8652, -65.78001, -65.69423, -65.60806, 
        -65.52025, -65.43307, -65.34575, -65.25803, -65.1713, -65.08651, 
        -65.00399, -64.92499, -64.84952, -64.77769, -64.70885, -64.64224, 
        -64.57693, -64.51243, -64.44833, -64.38426, -64.31993, -64.25523, 
        -64.19009, -64.12486, -64.05984, -63.99548, -63.93141, -63.86719, 
        -63.80186, -63.73442, -63.66377, -63.58897, -63.50959, -63.42561, 
        -63.33684, -63.24356, -63.14678, -63.04584, -62.94406, -62.84127, 
        -62.73827, -62.63566, -62.53385, -62.43303, -62.33368, -62.23624, 
        -62.14103, -62.04823, -61.95822, -61.87159, -61.78867, -61.70903, 
        -61.63246, -61.55829, -61.48588, -61.41415, -61.34232, -61.26989, 
        -61.19646, -61.12221, -61.04726, -60.97235, -60.89774, -60.82455, 
        -60.75343, -60.68494, -60.61945, -60.55722, -60.49874, -60.44433, 
        -60.39403, -60.34806, -60.30622, -60.26846, -60.2348, -60.20528, 
        -60.18006, -60.15802, -60.14103, -60.1267, -60.1136, -60.1008, 
        -60.08745, -60.07256, -60.05565, -60.03643, -60.01595, -59.99488, 
        -59.97486, -59.95682, -59.94148, -59.92928, -59.92079, -59.91641, 
        -59.91616,
  -49.80815, -49.99351, -50.17785, -50.36255, -50.54985, -50.7413, 
        -50.93906, -51.14351, -51.35292, -51.56955, -51.79162, -52.01862, 
        -52.25054, -52.48764, -52.73044, -52.97899, -53.23431, -53.49701, 
        -53.76706, -54.04479, -54.33021, -54.62322, -54.92284, -55.22647, 
        -55.5342, -55.84264, -56.14957, -56.45282, -56.75044, -57.04077, 
        -57.32119, -57.5891, -57.84316, -58.08269, -58.30724, -58.51748, 
        -58.71425, -58.89924, -59.07287, -59.23942, -59.39954, -59.55448, 
        -59.70558, -59.853, -59.99677, -60.13685, -60.27279, -60.40428, 
        -60.53094, -60.65274, -60.76976, -60.88236, -60.99113, -61.09671, 
        -61.19872, -61.29907, -61.39668, -61.49126, -61.58291, -61.67165, 
        -61.75797, -61.84233, -61.92651, -62.00957, -62.09238, -62.17422, 
        -62.25555, -62.33615, -62.41609, -62.49599, -62.57566, -62.65497, 
        -62.73569, -62.81768, -62.90121, -62.98654, -63.07416, -63.16447, 
        -63.25746, -63.35269, -63.44967, -63.5482, -63.64853, -63.75063, 
        -63.85484, -63.96112, -64.06979, -64.17989, -64.29063, -64.40015, 
        -64.50962, -64.61691, -64.72093, -64.8213, -64.91805, -65.01113, 
        -65.10054, -65.18665, -65.27029, -65.35165, -65.4314, -65.51079, 
        -65.59075, -65.67189, -65.75468, -65.83936, -65.92545, -66.01249, 
        -66.0985, -66.18481, -66.26966, -66.35169, -66.43031, -66.50503, 
        -66.57555, -66.64194, -66.70469, -66.76427, -66.8218, -66.87818, 
        -66.93401, -66.98994, -67.0461, -67.10334, -67.16212, -67.22227, 
        -67.28432, -67.34772, -67.41158, -67.47716, -67.5428, -67.60827, 
        -67.67299, -67.73716, -67.80042, -67.86251, -67.92333, -67.98299, 
        -68.04121, -68.0976, -68.15138, -68.20258, -68.2506, -68.29514, 
        -68.33624, -68.37344, -68.40656, -68.43533, -68.45953, -68.47993, 
        -68.49548, -68.50851, -68.51801, -68.5242, -68.52717, -68.52656, 
        -68.52265, -68.51511, -68.50436, -68.49068, -68.47399, -68.4545, 
        -68.43207, -68.40718, -68.3802, -68.35113, -68.32057, -68.28815, 
        -68.25408, -68.21886, -68.18224, -68.1444, -68.10552, -68.06567, 
        -68.02405, -67.9819, -67.93826, -67.89265, -67.84505, -67.79542, 
        -67.74339, -67.68926, -67.6328, -67.5739, -67.51257, -67.4483, 
        -67.38129, -67.31176, -67.23986, -67.16589, -67.09019, -67.01341, 
        -66.93587, -66.85827, -66.78128, -66.7044, -66.62763, -66.55077, 
        -66.4738, -66.39659, -66.31732, -66.23805, -66.15688, -66.07402, 
        -65.98926, -65.90313, -65.81589, -65.72744, -65.63777, -65.54691, 
        -65.45492, -65.3616, -65.26722, -65.17257, -65.07879, -64.98667, 
        -64.89742, -64.81157, -64.72978, -64.65212, -64.57757, -64.50544, 
        -64.43488, -64.36539, -64.29659, -64.22796, -64.15942, -64.09092, 
        -64.02247, -63.95452, -63.88732, -63.82007, -63.75423, -63.68822, 
        -63.62091, -63.55102, -63.47771, -63.3999, -63.31722, -63.22965, 
        -63.13713, -63.04013, -62.93949, -62.83633, -62.73169, -62.62645, 
        -62.52146, -62.41747, -62.31446, -62.21314, -62.11359, -62.01614, 
        -61.92104, -61.82888, -61.74041, -61.6555, -61.57436, -61.49711, 
        -61.42331, -61.35259, -61.28377, -61.21616, -61.14876, -61.08083, 
        -61.01199, -60.94166, -60.8701, -60.79793, -60.72488, -60.65411, 
        -60.58566, -60.5201, -60.45775, -60.39883, -60.34399, -60.29325, 
        -60.2467, -60.20424, -60.16554, -60.13038, -60.099, -60.07163, 
        -60.04818, -60.02884, -60.01309, -59.99955, -59.98709, -59.97463, 
        -59.96115, -59.94613, -59.92914, -59.91041, -59.89058, -59.87058, 
        -59.85161, -59.83456, -59.82048, -59.80978, -59.80313, -59.80098, 
        -59.80346,
  -49.59059, -49.78035, -49.96921, -50.15747, -50.34888, -50.54456, 
        -50.74604, -50.95422, -51.16904, -51.38975, -51.61631, -51.84812, 
        -52.08502, -52.32721, -52.57512, -52.82932, -53.08963, -53.35638, 
        -53.63146, -53.91402, -54.20432, -54.50175, -54.80571, -55.11443, 
        -55.42571, -55.73721, -56.04673, -56.352, -56.65134, -56.94304, 
        -57.22459, -57.49328, -57.74688, -57.98651, -58.21107, -58.42138, 
        -58.61807, -58.80297, -58.9774, -59.14341, -59.30279, -59.45673, 
        -59.6065, -59.7523, -59.89437, -60.03267, -60.16692, -60.29686, 
        -60.42088, -60.54087, -60.65577, -60.76594, -60.87191, -60.97444, 
        -61.07417, -61.17122, -61.26577, -61.35749, -61.44658, -61.53326, 
        -61.61809, -61.7017, -61.78452, -61.86703, -61.94915, -62.03006, 
        -62.112, -62.19375, -62.27557, -62.35756, -62.43947, -62.52184, 
        -62.60481, -62.68863, -62.77381, -62.86034, -62.94926, -63.04094, 
        -63.13512, -63.23153, -63.33005, -63.43094, -63.53377, -63.63847, 
        -63.74657, -63.85743, -63.9701, -64.08464, -64.1998, -64.31448, 
        -64.42765, -64.53837, -64.64555, -64.74899, -64.8485, -64.94386, 
        -65.03522, -65.12274, -65.20678, -65.28803, -65.36698, -65.44389, 
        -65.52178, -65.60126, -65.68279, -65.76635, -65.85198, -65.93912, 
        -66.02664, -66.11336, -66.19848, -66.28039, -66.35806, -66.4312, 
        -66.49982, -66.56424, -66.62495, -66.68269, -66.73853, -66.79366, 
        -66.84846, -66.90317, -66.95901, -67.01603, -67.07455, -67.13483, 
        -67.19708, -67.26091, -67.32642, -67.393, -67.4603, -67.52819, 
        -67.59564, -67.66253, -67.72875, -67.79356, -67.85703, -67.91909, 
        -67.97953, -68.03783, -68.09334, -68.14591, -68.19367, -68.23892, 
        -68.28071, -68.31824, -68.35152, -68.38023, -68.40418, -68.42401, 
        -68.43991, -68.4524, -68.46124, -68.46672, -68.46885, -68.46741, 
        -68.46263, -68.45413, -68.44241, -68.42754, -68.4095, -68.38866, 
        -68.36494, -68.33872, -68.31068, -68.27991, -68.24906, -68.21677, 
        -68.18295, -68.14788, -68.11133, -68.07368, -68.03462, -67.99441, 
        -67.95308, -67.91042, -67.8664, -67.82066, -67.77309, -67.72359, 
        -67.67194, -67.61852, -67.56297, -67.50507, -67.44496, -67.38242, 
        -67.31728, -67.24957, -67.1798, -67.10834, -67.034, -66.95936, 
        -66.88353, -66.80723, -66.73093, -66.65417, -66.57742, -66.50023, 
        -66.42255, -66.34435, -66.26506, -66.18439, -66.10194, -66.01766, 
        -65.93182, -65.84406, -65.7549, -65.66344, -65.57035, -65.47527, 
        -65.378, -65.27921, -65.17892, -65.07823, -64.97803, -64.87946, 
        -64.78373, -64.69103, -64.60236, -64.5166, -64.43555, -64.35697, 
        -64.28022, -64.20487, -64.13023, -64.05609, -63.98251, -63.90932, 
        -63.83672, -63.76529, -63.69487, -63.62561, -63.55712, -63.48861, 
        -63.41859, -63.34596, -63.26962, -63.18859, -63.10258, -63.01133, 
        -62.9151, -62.81463, -62.71066, -62.60456, -62.49757, -62.39034, 
        -62.28377, -62.1784, -62.07477, -61.97302, -61.87378, -61.77699, 
        -61.68288, -61.59122, -61.50465, -61.42207, -61.34382, -61.26947, 
        -61.19925, -61.13224, -61.06752, -61.00437, -60.94177, -60.87865, 
        -60.81446, -60.74861, -60.68099, -60.61231, -60.54324, -60.47549, 
        -60.41006, -60.34773, -60.2888, -60.23347, -60.18227, -60.13534, 
        -60.09272, -60.05377, -60.01813, -59.98583, -59.95681, -59.93131, 
        -59.90957, -59.89149, -59.87624, -59.86275, -59.84986, -59.83649, 
        -59.82196, -59.80592, -59.78826, -59.76931, -59.74976, -59.73058, 
        -59.71286, -59.69739, -59.6852, -59.6766, -59.67166, -59.67244, 
        -59.67821,
  -49.36135, -49.55561, -49.74847, -49.94146, -50.13681, -50.33605, 
        -50.54083, -50.7521, -50.97044, -51.19503, -51.42568, -51.66209, 
        -51.90291, -52.15024, -52.40321, -52.66278, -52.9284, -53.2008, 
        -53.48069, -53.76787, -54.06226, -54.36349, -54.67093, -54.98293, 
        -55.29731, -55.61149, -55.92333, -56.22976, -56.53089, -56.82406, 
        -57.10694, -57.377, -57.63252, -57.87296, -58.09838, -58.30941, 
        -58.50691, -58.69244, -58.86757, -59.03406, -59.19366, -59.34763, 
        -59.49668, -59.64053, -59.78126, -59.91812, -60.05075, -60.17893, 
        -60.30198, -60.41956, -60.53198, -60.639, -60.74181, -60.84066, 
        -60.93658, -61.02972, -61.12034, -61.20834, -61.29401, -61.3769, 
        -61.45947, -61.54122, -61.62255, -61.70369, -61.78502, -61.86656, 
        -61.9488, -62.03172, -62.11509, -62.19884, -62.28281, -62.36715, 
        -62.45203, -62.5377, -62.62426, -62.71241, -62.80169, -62.89438, 
        -62.98929, -63.08691, -63.1871, -63.29016, -63.39634, -63.50569, 
        -63.6185, -63.73405, -63.85225, -63.97165, -64.09149, -64.21072, 
        -64.32802, -64.44296, -64.55432, -64.66139, -64.76335, -64.86185, 
        -64.95565, -65.04489, -65.12984, -65.21111, -65.28913, -65.36555, 
        -65.4416, -65.51904, -65.59854, -65.68063, -65.7655, -65.8522, 
        -65.93961, -66.02629, -66.1106, -66.19121, -66.26743, -66.33854, 
        -66.40408, -66.46601, -66.52448, -66.58041, -66.63466, -66.68858, 
        -66.74291, -66.798, -66.85412, -66.91129, -66.96981, -67.02992, 
        -67.09229, -67.15662, -67.22253, -67.29, -67.35887, -67.42882, 
        -67.49885, -67.56818, -67.63599, -67.70354, -67.76991, -67.8345, 
        -67.89683, -67.95672, -68.0136, -68.06731, -68.11739, -68.16342, 
        -68.2056, -68.24325, -68.27655, -68.30511, -68.32874, -68.34809, 
        -68.3634, -68.37518, -68.38354, -68.38837, -68.38983, -68.38776, 
        -68.38139, -68.37238, -68.35977, -68.34377, -68.32446, -68.30238, 
        -68.27742, -68.25008, -68.22103, -68.19064, -68.15938, -68.1272, 
        -68.09351, -68.05835, -68.02148, -67.98342, -67.94426, -67.90364, 
        -67.86176, -67.81829, -67.77372, -67.7279, -67.6804, -67.63156, 
        -67.58041, -67.5266, -67.47238, -67.41581, -67.35728, -67.2963, 
        -67.23321, -67.16811, -67.10052, -67.03123, -66.96031, -66.88788, 
        -66.81425, -66.73947, -66.66396, -66.58764, -66.5108, -66.43353, 
        -66.35557, -66.27665, -66.19643, -66.11465, -66.03111, -65.94582, 
        -65.85881, -65.76981, -65.6785, -65.58517, -65.48791, -65.38889, 
        -65.28708, -65.18326, -65.07803, -64.97185, -64.8663, -64.76198, 
        -64.66012, -64.56111, -64.46548, -64.3735, -64.28481, -64.19899, 
        -64.11513, -64.03268, -63.95133, -63.87096, -63.79134, -63.71283, 
        -63.6354, -63.55934, -63.48487, -63.41187, -63.33974, -63.26768, 
        -63.19424, -63.11816, -63.03833, -62.95399, -62.86434, -62.76955, 
        -62.6688, -62.5651, -62.45823, -62.34965, -62.24043, -62.13148, 
        -62.02368, -61.91734, -61.8132, -61.71154, -61.613, -61.51741, 
        -61.42525, -61.33696, -61.25293, -61.17349, -61.09877, -61.02858, 
        -60.96238, -60.89964, -60.8395, -60.78107, -60.72339, -60.66535, 
        -60.6061, -60.54497, -60.48199, -60.41737, -60.35226, -60.28803, 
        -60.22615, -60.16745, -60.11224, -60.06077, -60.01335, -59.97025, 
        -59.93124, -59.89553, -59.86313, -59.83366, -59.80611, -59.7825, 
        -59.76218, -59.74465, -59.72939, -59.71523, -59.70116, -59.68624, 
        -59.66999, -59.65215, -59.63306, -59.61329, -59.59364, -59.57506, 
        -59.55862, -59.54502, -59.53516, -59.52967, -59.5287, -59.53294, 
        -59.54238,
  -49.12476, -49.32315, -49.51941, -49.71573, -49.91404, -50.11634, 
        -50.32404, -50.53708, -50.75813, -50.98612, -51.22049, -51.46099, 
        -51.70752, -51.96002, -52.21798, -52.48216, -52.75279, -53.03017, 
        -53.314, -53.60506, -53.90319, -54.20768, -54.51693, -54.83151, 
        -55.1481, -55.46441, -55.77842, -56.08796, -56.39116, -56.68611, 
        -56.9706, -57.24222, -57.49927, -57.74137, -57.96845, -58.18105, 
        -58.38023, -58.56644, -58.74335, -58.91159, -59.07248, -59.22715, 
        -59.37644, -59.52094, -59.66091, -59.79657, -59.92762, -60.0537, 
        -60.1743, -60.28915, -60.39833, -60.50197, -60.60094, -60.69485, 
        -60.78645, -60.87501, -60.96101, -61.04476, -61.12643, -61.20682, 
        -61.28647, -61.36567, -61.44498, -61.52435, -61.60418, -61.68511, 
        -61.7676, -61.85109, -61.93542, -62.02052, -62.10465, -62.19059, 
        -62.27674, -62.36349, -62.45154, -62.54093, -62.6319, -62.72531, 
        -62.82149, -62.92033, -63.02232, -63.1278, -63.23716, -63.35081, 
        -63.46888, -63.59022, -63.71394, -63.83875, -63.96266, -64.08707, 
        -64.2094, -64.32909, -64.44526, -64.55717, -64.66464, -64.76685, 
        -64.86375, -64.95538, -65.04171, -65.12337, -65.20101, -65.27585, 
        -65.34998, -65.42505, -65.50229, -65.58243, -65.66572, -65.75024, 
        -65.8367, -65.92232, -66.0051, -66.08364, -66.15733, -66.22604, 
        -66.28987, -66.34931, -66.4052, -66.45912, -66.51207, -66.56512, 
        -66.61902, -66.67431, -66.73073, -66.78825, -66.8472, -66.90775, 
        -66.97032, -67.03379, -67.1002, -67.16898, -67.23917, -67.31039, 
        -67.38212, -67.45398, -67.52568, -67.59609, -67.66463, -67.73096, 
        -67.79517, -67.85664, -67.91483, -67.96969, -68.02056, -68.06731, 
        -68.10965, -68.14726, -68.18018, -68.20808, -68.23033, -68.24929, 
        -68.26432, -68.27557, -68.28342, -68.28772, -68.28879, -68.28627, 
        -68.28006, -68.27017, -68.25664, -68.23973, -68.21933, -68.19585, 
        -68.16974, -68.14137, -68.11147, -68.08073, -68.04901, -68.01663, 
        -67.98283, -67.94766, -67.9106, -67.87192, -67.83079, -67.7894, 
        -67.74702, -67.70332, -67.65857, -67.61278, -67.56568, -67.51729, 
        -67.46746, -67.41551, -67.36208, -67.30701, -67.25036, -67.19157, 
        -67.13049, -67.06743, -67.00242, -66.93567, -66.86689, -66.79676, 
        -66.72514, -66.65205, -66.57777, -66.50224, -66.42561, -66.34831, 
        -66.26881, -66.18963, -66.10905, -66.02673, -65.94225, -65.85592, 
        -65.76764, -65.67722, -65.58437, -65.48882, -65.38974, -65.28775, 
        -65.18244, -65.07455, -64.96446, -64.85384, -64.74346, -64.63387, 
        -64.52618, -64.42114, -64.31894, -64.2199, -64.12364, -64.02998, 
        -63.93796, -63.84785, -63.75898, -63.67164, -63.58554, -63.50087, 
        -63.41674, -63.33579, -63.2564, -63.17876, -63.10217, -63.02563, 
        -62.94808, -62.86802, -62.78423, -62.69598, -62.60269, -62.50436, 
        -62.40143, -62.29469, -62.1852, -62.07425, -61.9632, -61.85308, 
        -61.74394, -61.63681, -61.53273, -61.43157, -61.33405, -61.24024, 
        -61.15059, -61.06542, -60.98502, -60.9094, -60.83873, -60.7731, 
        -60.71175, -60.65376, -60.59847, -60.5451, -60.49251, -60.43974, 
        -60.38584, -60.329, -60.27098, -60.21128, -60.15075, -60.09104, 
        -60.03331, -59.97872, -59.92762, -59.88028, -59.83665, -59.79709, 
        -59.76138, -59.72905, -59.69962, -59.67283, -59.64852, -59.62675, 
        -59.60735, -59.59014, -59.57438, -59.55904, -59.54322, -59.52603, 
        -59.50723, -59.48705, -59.466, -59.44509, -59.42507, -59.40702, 
        -59.39188, -59.38046, -59.37337, -59.37107, -59.37399, -59.38185, 
        -59.39531,
  -48.88103, -49.08317, -49.28144, -49.48052, -49.68127, -49.88588, 
        -50.09565, -50.31187, -50.53521, -50.76586, -51.00375, -51.24807, 
        -51.49863, -51.75547, -52.01821, -52.28662, -52.56032, -52.8417, 
        -53.12966, -53.42379, -53.72501, -54.03233, -54.34455, -54.66113, 
        -54.97953, -55.29783, -55.61368, -55.92534, -56.23071, -56.52772, 
        -56.8142, -57.087, -57.34655, -57.59106, -57.82071, -58.03601, 
        -58.23792, -58.42801, -58.60769, -58.77856, -58.94181, -59.09822, 
        -59.24865, -59.39349, -59.53309, -59.66768, -59.79694, -59.91956, 
        -60.03752, -60.14915, -60.25449, -60.35414, -60.44895, -60.5394, 
        -60.62617, -60.70974, -60.79085, -60.8698, -60.94711, -61.02356, 
        -61.09986, -61.17625, -61.25302, -61.3305, -61.40786, -61.4877, 
        -61.56936, -61.65265, -61.73715, -61.8226, -61.90826, -61.9945, 
        -62.08142, -62.16901, -62.25773, -62.34768, -62.43921, -62.53349, 
        -62.63074, -62.7309, -62.83468, -62.94164, -63.05471, -63.17301, 
        -63.29612, -63.4232, -63.55264, -63.68316, -63.81399, -63.94394, 
        -64.07198, -64.19735, -64.31955, -64.43712, -64.55009, -64.65725, 
        -64.75847, -64.85333, -64.94178, -65.02424, -65.10052, -65.17413, 
        -65.24622, -65.31882, -65.39344, -65.4712, -65.55209, -65.63543, 
        -65.72002, -65.80315, -65.88318, -65.95898, -66.02978, -66.09531, 
        -66.15603, -66.21245, -66.26601, -66.31815, -66.36987, -66.42155, 
        -66.47558, -66.5311, -66.58814, -66.64654, -66.70624, -66.7674, 
        -66.83014, -66.89513, -66.96246, -67.03187, -67.10313, -67.17577, 
        -67.24941, -67.32356, -67.39738, -67.46975, -67.54, -67.60847, 
        -67.6739, -67.7366, -67.79492, -67.85052, -67.90192, -67.94894, 
        -67.9912, -68.02853, -68.06072, -68.08815, -68.11091, -68.1293, 
        -68.14391, -68.15495, -68.16254, -68.16641, -68.16681, -68.16349, 
        -68.15642, -68.14583, -68.13126, -68.11301, -68.0915, -68.06696, 
        -68.03996, -68.00993, -67.97938, -67.94778, -67.9156, -67.88282, 
        -67.84889, -67.81332, -67.77578, -67.7364, -67.69554, -67.65327, 
        -67.61012, -67.56622, -67.52167, -67.47659, -67.43037, -67.38293, 
        -67.33385, -67.28305, -67.2311, -67.1775, -67.12221, -67.06551, 
        -67.00675, -66.94612, -66.88254, -66.81812, -66.7518, -66.68377, 
        -66.6141, -66.54278, -66.46992, -66.39549, -66.31953, -66.24266, 
        -66.16443, -66.08491, -66.00394, -65.9212, -65.83647, -65.74913, 
        -65.65959, -65.56759, -65.4727, -65.37511, -65.27394, -65.16917, 
        -65.06091, -64.94954, -64.83617, -64.72146, -64.60638, -64.4923, 
        -64.37912, -64.26697, -64.15845, -64.05238, -63.94867, -63.84701, 
        -63.74723, -63.64902, -63.55222, -63.45728, -63.36404, -63.27308, 
        -63.18422, -63.09741, -63.0127, -62.92967, -62.84795, -62.76637, 
        -62.68383, -62.59917, -62.5109, -62.41851, -62.32133, -62.21954, 
        -62.11338, -62.00385, -61.89196, -61.77907, -61.66616, -61.5544, 
        -61.44444, -61.33707, -61.23311, -61.13266, -61.03669, -60.94428, 
        -60.8576, -60.77603, -60.69979, -60.62869, -60.56284, -60.50209, 
        -60.44577, -60.39325, -60.34343, -60.29513, -60.24784, -60.20054, 
        -60.15221, -60.10201, -60.04968, -59.99553, -59.94057, -59.88597, 
        -59.83331, -59.78331, -59.73669, -59.6935, -59.65385, -59.61782, 
        -59.58524, -59.55576, -59.52902, -59.50456, -59.4822, -59.46178, 
        -59.44305, -59.42558, -59.40888, -59.39188, -59.37373, -59.35381, 
        -59.33238, -59.30958, -59.28656, -59.26409, -59.2437, -59.22627, 
        -59.21144, -59.20221, -59.19804, -59.19915, -59.20565, -59.21785, 
        -59.23513,
  -48.62983, -48.83522, -49.03693, -49.23841, -49.44106, -49.64748, 
        -49.85894, -50.07688, -50.30194, -50.53475, -50.77552, -51.02206, 
        -51.27619, -51.53661, -51.80309, -52.07515, -52.35298, -52.63771, 
        -52.92844, -53.22537, -53.52861, -53.83781, -54.15187, -54.46972, 
        -54.7896, -55.10949, -55.42646, -55.74059, -56.04839, -56.348, 
        -56.63699, -56.91376, -57.1765, -57.42458, -57.65806, -57.87696, 
        -58.08279, -58.27659, -58.46005, -58.63445, -58.80089, -58.95985, 
        -59.11102, -59.25683, -59.39638, -59.52995, -59.6573, -59.7783, 
        -59.89282, -60.00051, -60.10184, -60.19716, -60.28727, -60.37287, 
        -60.45451, -60.53304, -60.60883, -60.68288, -60.75479, -60.82724, 
        -60.90021, -60.97355, -61.04801, -61.12336, -61.20003, -61.27828, 
        -61.35846, -61.44036, -61.5237, -61.60817, -61.69331, -61.77912, 
        -61.86572, -61.9535, -62.04211, -62.13134, -62.22348, -62.31854, 
        -62.41655, -62.51791, -62.62374, -62.73455, -62.85117, -62.97378, 
        -63.1017, -63.23399, -63.36909, -63.5058, -63.6426, -63.7788, 
        -63.91359, -64.04559, -64.17437, -64.29821, -64.41764, -64.53125, 
        -64.63786, -64.73695, -64.82815, -64.9117, -64.98923, -65.062, 
        -65.13222, -65.20245, -65.27422, -65.34891, -65.42662, -65.50687, 
        -65.58757, -65.66725, -65.74358, -65.81573, -65.88189, -65.94376, 
        -66.00108, -66.05473, -66.10593, -66.15637, -66.20737, -66.25986, 
        -66.31422, -66.37042, -66.42857, -66.48818, -66.54882, -66.6106, 
        -66.67408, -66.73984, -66.8079, -66.87812, -66.95064, -67.0245, 
        -67.09967, -67.17451, -67.25011, -67.32439, -67.39638, -67.46575, 
        -67.53238, -67.59589, -67.65574, -67.71171, -67.76331, -67.81017, 
        -67.85204, -67.88892, -67.92058, -67.94734, -67.96941, -67.9873, 
        -68.00167, -68.01226, -68.01907, -68.02242, -68.02195, -68.01685, 
        -68.00892, -67.99704, -67.9813, -67.96185, -67.93937, -67.91402, 
        -67.88617, -67.85635, -67.82499, -67.79287, -67.76015, -67.72669, 
        -67.692, -67.6559, -67.61796, -67.57798, -67.53629, -67.49338, 
        -67.4496, -67.40585, -67.36193, -67.31771, -67.27262, -67.22527, 
        -67.17749, -67.12805, -67.07723, -67.02526, -66.97171, -66.91676, 
        -66.86018, -66.80185, -66.74169, -66.67973, -66.61591, -66.55009, 
        -66.48228, -66.41272, -66.34127, -66.2686, -66.1941, -66.11788, 
        -66.04019, -65.96072, -65.87957, -65.79662, -65.71142, -65.62347, 
        -65.53275, -65.43919, -65.34122, -65.24116, -65.13744, -65.03015, 
        -64.9198, -64.80575, -64.6897, -64.57143, -64.45245, -64.33354, 
        -64.21549, -64.09856, -63.98339, -63.87035, -63.75945, -63.65024, 
        -63.54259, -63.43664, -63.33233, -63.23003, -63.12983, -63.03204, 
        -62.93675, -62.84396, -62.75348, -62.66489, -62.57753, -62.49031, 
        -62.40236, -62.31249, -62.21966, -62.1229, -62.02071, -61.91526, 
        -61.80606, -61.694, -61.57994, -61.46502, -61.35052, -61.23735, 
        -61.12664, -61.01883, -60.91502, -60.81562, -60.72142, -60.63251, 
        -60.54911, -60.4716, -60.39968, -60.33375, -60.27321, -60.21762, 
        -60.16679, -60.11956, -60.07519, -60.03224, -59.99037, -59.94883, 
        -59.90629, -59.86225, -59.81612, -59.76836, -59.71952, -59.67107, 
        -59.62403, -59.57946, -59.53756, -59.49882, -59.46316, -59.4306, 
        -59.40095, -59.37298, -59.34835, -59.32572, -59.3048, -59.28522, 
        -59.26661, -59.24852, -59.23028, -59.21106, -59.19032, -59.16766, 
        -59.14352, -59.11813, -59.09328, -59.07008, -59.04956, -59.03242, 
        -59.01989, -59.01264, -59.0111, -59.01538, -59.02561, -59.04147, 
        -59.06282,
  -48.374, -48.58168, -48.78576, -48.98853, -49.19286, -49.40046, 
        -49.61197, -49.83088, -50.05697, -50.2913, -50.5339, -50.78391, 
        -51.04096, -51.30408, -51.57334, -51.8484, -52.12901, -52.41546, 
        -52.70816, -53.00672, -53.3115, -53.62091, -53.93609, -54.25525, 
        -54.57672, -54.89867, -55.21892, -55.53565, -55.84647, -56.14913, 
        -56.44138, -56.72168, -56.98869, -57.24127, -57.47929, -57.70306, 
        -57.91253, -58.11108, -58.29904, -58.47784, -58.64815, -58.81033, 
        -58.965, -59.11213, -59.25191, -59.38446, -59.50962, -59.62764, 
        -59.73827, -59.84177, -59.9385, -60.02886, -60.11266, -60.19299, 
        -60.26928, -60.34256, -60.41356, -60.48319, -60.55214, -60.62115, 
        -60.69104, -60.76207, -60.83418, -60.90732, -60.98174, -61.0576, 
        -61.13504, -61.21424, -61.29498, -61.37607, -61.45925, -61.54391, 
        -61.62962, -61.71674, -61.80518, -61.89544, -61.98795, -62.0832, 
        -62.18201, -62.28476, -62.39242, -62.50581, -62.62539, -62.75164, 
        -62.88376, -63.0209, -63.16135, -63.30292, -63.4464, -63.58964, 
        -63.73175, -63.87152, -64.00826, -64.14109, -64.26873, -64.38964, 
        -64.50253, -64.60645, -64.70113, -64.78689, -64.86517, -64.93763, 
        -65.00652, -65.07455, -65.14328, -65.2133, -65.28684, -65.36225, 
        -65.43832, -65.51299, -65.58469, -65.65226, -65.71492, -65.77303, 
        -65.82679, -65.87749, -65.92681, -65.97594, -66.02646, -66.07885, 
        -66.13387, -66.19118, -66.25056, -66.31149, -66.37331, -66.43528, 
        -66.50002, -66.56671, -66.63588, -66.70711, -66.7806, -66.8561, 
        -66.93288, -67.01038, -67.08734, -67.16278, -67.23597, -67.30616, 
        -67.37333, -67.43695, -67.49676, -67.55252, -67.60385, -67.65051, 
        -67.69196, -67.72829, -67.75937, -67.78444, -67.80594, -67.82327, 
        -67.83662, -67.84634, -67.85222, -67.85467, -67.85321, -67.8478, 
        -67.83846, -67.82522, -67.80827, -67.78783, -67.76431, -67.73804, 
        -67.70941, -67.67903, -67.64709, -67.61417, -67.58059, -67.5462, 
        -67.51093, -67.47395, -67.43403, -67.39323, -67.35102, -67.30795, 
        -67.26446, -67.22081, -67.17737, -67.13407, -67.09048, -67.04571, 
        -66.99934, -66.95143, -66.90213, -66.85178, -66.80021, -66.74715, 
        -66.69238, -66.63593, -66.57848, -66.51904, -66.45757, -66.39377, 
        -66.32803, -66.26055, -66.1913, -66.12005, -66.04609, -65.97119, 
        -65.89439, -65.81535, -65.73434, -65.65102, -65.56499, -65.4763, 
        -65.3844, -65.28901, -65.19008, -65.08759, -64.98173, -64.87218, 
        -64.75949, -64.64354, -64.52494, -64.40416, -64.28185, -64.15882, 
        -64.03548, -63.91272, -63.7913, -63.67123, -63.55283, -63.43611, 
        -63.32099, -63.20789, -63.09671, -62.9876, -62.88004, -62.77586, 
        -62.67445, -62.57544, -62.47874, -62.38411, -62.29082, -62.19793, 
        -62.10442, -62.00924, -61.91133, -61.80996, -61.7049, -61.596, 
        -61.48369, -61.36905, -61.25275, -61.13598, -61.01977, -60.90542, 
        -60.79387, -60.68599, -60.58265, -60.48456, -60.39225, -60.30615, 
        -60.22635, -60.15281, -60.08564, -60.02462, -59.96922, -59.91894, 
        -59.87302, -59.83094, -59.79164, -59.75443, -59.71716, -59.6814, 
        -59.64519, -59.60767, -59.56846, -59.52773, -59.48583, -59.44402, 
        -59.40337, -59.36451, -59.32803, -59.29396, -59.26247, -59.23343, 
        -59.2067, -59.18206, -59.15927, -59.13793, -59.11769, -59.09818, 
        -59.079, -59.05971, -59.03971, -59.01835, -58.99499, -58.96978, 
        -58.94317, -58.91612, -58.88994, -58.866, -58.84517, -58.82848, 
        -58.8168, -58.81079, -58.81113, -58.81794, -58.8311, -58.85038, 
        -58.87516,
  -48.11349, -48.32191, -48.52683, -48.73044, -48.93564, -49.14375, 
        -49.35697, -49.57645, -49.80338, -50.03823, -50.28189, -50.53352, 
        -50.79261, -51.05781, -51.32897, -51.60483, -51.88704, -52.17485, 
        -52.46856, -52.76787, -53.07351, -53.38457, -53.70096, -54.02099, 
        -54.34388, -54.66789, -54.99088, -55.31059, -55.62462, -55.93078, 
        -56.22595, -56.51054, -56.78244, -57.04035, -57.2841, -57.5135, 
        -57.72943, -57.93321, -58.12604, -58.30946, -58.48402, -58.65001, 
        -58.80754, -58.95632, -59.09631, -59.22765, -59.34937, -59.46374, 
        -59.5702, -59.66909, -59.76078, -59.84598, -59.92549, -60.00042, 
        -60.07159, -60.13994, -60.20667, -60.27229, -60.33791, -60.40408, 
        -60.47142, -60.54018, -60.61026, -60.68008, -60.75182, -60.82447, 
        -60.89834, -60.9735, -61.05017, -61.12868, -61.20884, -61.29131, 
        -61.3755, -61.46173, -61.5499, -61.63969, -61.73197, -61.82735, 
        -61.92663, -62.0304, -62.13874, -62.25442, -62.37669, -62.50572, 
        -62.64117, -62.78215, -62.92752, -63.07594, -63.22625, -63.37704, 
        -63.52724, -63.67564, -63.82145, -63.96355, -64.10014, -64.22944, 
        -64.34946, -64.45921, -64.55827, -64.64594, -64.72597, -64.79894, 
        -64.86703, -64.93281, -64.99811, -65.06458, -65.13297, -65.20259, 
        -65.27245, -65.3412, -65.40718, -65.46943, -65.52728, -65.58105, 
        -65.63165, -65.68, -65.72768, -65.77583, -65.82494, -65.87782, 
        -65.93374, -65.9925, -66.05346, -66.1158, -66.17937, -66.24394, 
        -66.31014, -66.37799, -66.44784, -66.5203, -66.59543, -66.67232, 
        -66.75059, -66.82936, -66.90734, -66.98357, -67.0575, -67.12824, 
        -67.19524, -67.25755, -67.3168, -67.37213, -67.42292, -67.46918, 
        -67.5104, -67.54617, -67.57687, -67.60233, -67.62303, -67.63945, 
        -67.65163, -67.66009, -67.66479, -67.66555, -67.66256, -67.65543, 
        -67.64441, -67.62956, -67.61112, -67.58945, -67.56484, -67.53778, 
        -67.50774, -67.47666, -67.44394, -67.41014, -67.37575, -67.34023, 
        -67.30356, -67.26539, -67.22533, -67.184, -67.14157, -67.09859, 
        -67.05544, -67.01254, -66.97014, -66.92792, -66.88559, -66.8425, 
        -66.79795, -66.7522, -66.70484, -66.65615, -66.60629, -66.55499, 
        -66.50236, -66.44748, -66.39175, -66.3344, -66.27494, -66.2138, 
        -66.15032, -66.08495, -66.01777, -65.9485, -65.87731, -65.80394, 
        -65.72813, -65.64996, -65.56905, -65.48542, -65.39878, -65.30877, 
        -65.21518, -65.11791, -65.01701, -64.9123, -64.80401, -64.69216, 
        -64.57711, -64.45931, -64.33854, -64.21545, -64.09012, -63.96222, 
        -63.8343, -63.70595, -63.57793, -63.45088, -63.32517, -63.20131, 
        -63.07946, -62.95994, -62.84266, -62.7277, -62.61539, -62.50573, 
        -62.3986, -62.29362, -62.19103, -62.09022, -61.99101, -61.89232, 
        -61.79326, -61.69286, -61.59003, -61.48429, -61.37551, -61.26318, 
        -61.148, -61.03068, -60.91222, -60.79372, -60.67598, -60.56048, 
        -60.4483, -60.34043, -60.23676, -60.13993, -60.04985, -59.96657, 
        -59.89011, -59.82041, -59.75775, -59.70152, -59.65079, -59.60543, 
        -59.56436, -59.52681, -59.49232, -59.46015, -59.42961, -59.3996, 
        -59.36961, -59.33887, -59.30684, -59.27359, -59.23933, -59.20489, 
        -59.17111, -59.13882, -59.10809, -59.07938, -59.05238, -59.02699, 
        -59.00314, -58.98057, -58.95905, -58.93829, -58.91795, -58.89777, 
        -58.87745, -58.85634, -58.83428, -58.81075, -58.78497, -58.75755, 
        -58.72902, -58.70076, -58.67392, -58.6488, -58.62814, -58.6117, 
        -58.60043, -58.5952, -58.59666, -58.60519, -58.62056, -58.64256, 
        -58.67053,
  -47.8465, -48.05705, -48.26222, -48.46601, -48.6712, -48.87985, 
        -49.09327, -49.31298, -49.54, -49.77481, -50.01778, -50.27031, 
        -50.52995, -50.79649, -51.06924, -51.347, -51.63022, -51.91855, 
        -52.21276, -52.5129, -52.81892, -53.13099, -53.44815, -53.76937, 
        -54.09405, -54.41902, -54.74414, -55.06675, -55.38406, -55.69379, 
        -55.99414, -56.28339, -56.5605, -56.82424, -57.074, -57.30959, 
        -57.5314, -57.74097, -57.9393, -58.12785, -58.30708, -58.47573, 
        -58.63585, -58.78577, -58.92567, -59.05529, -59.175, -59.28519, 
        -59.38696, -59.48046, -59.56686, -59.64692, -59.72141, -59.79135, 
        -59.85809, -59.92265, -59.98597, -60.04774, -60.11082, -60.17501, 
        -60.24047, -60.30714, -60.3749, -60.44319, -60.51178, -60.58061, 
        -60.65006, -60.72034, -60.79233, -60.86632, -60.94263, -61.02186, 
        -61.10371, -61.1885, -61.2745, -61.36358, -61.45529, -61.55054, 
        -61.64996, -61.75451, -61.86486, -61.98197, -62.10586, -62.23693, 
        -62.37493, -62.51946, -62.66925, -62.82343, -62.98058, -63.13927, 
        -63.29821, -63.45609, -63.61072, -63.76279, -63.90902, -64.04736, 
        -64.17565, -64.29226, -64.39689, -64.48977, -64.57247, -64.64647, 
        -64.71412, -64.7775, -64.83911, -64.90063, -64.96285, -65.02587, 
        -65.08865, -65.15067, -65.21007, -65.26513, -65.31789, -65.36753, 
        -65.41508, -65.46126, -65.50723, -65.55487, -65.60509, -65.65885, 
        -65.71583, -65.77593, -65.83853, -65.90281, -65.96873, -66.03526, 
        -66.10291, -66.17197, -66.24332, -66.3177, -66.39439, -66.47175, 
        -66.55106, -66.63057, -66.70937, -66.78616, -66.86006, -66.93047, 
        -66.99706, -67.05989, -67.1187, -67.17342, -67.22379, -67.2695, 
        -67.31026, -67.34576, -67.37583, -67.40079, -67.42058, -67.4359, 
        -67.44679, -67.45351, -67.45621, -67.45381, -67.44852, -67.43921, 
        -67.42589, -67.40878, -67.38846, -67.36545, -67.33987, -67.31209, 
        -67.28223, -67.25057, -67.21726, -67.18277, -67.14703, -67.11017, 
        -67.07196, -67.03241, -66.9914, -66.94934, -66.90664, -66.86388, 
        -66.82148, -66.77962, -66.73856, -66.69786, -66.65627, -66.61492, 
        -66.57285, -66.52917, -66.48376, -66.43701, -66.3894, -66.34006, 
        -66.2893, -66.23743, -66.18375, -66.12859, -66.07133, -66.01234, 
        -65.95108, -65.88789, -65.8227, -65.75552, -65.68607, -65.61404, 
        -65.53934, -65.46207, -65.38168, -65.29771, -65.21002, -65.11831, 
        -65.02301, -64.92251, -64.81916, -64.71198, -64.6012, -64.48727, 
        -64.37013, -64.25012, -64.12734, -64.00176, -63.87382, -63.74343, 
        -63.61103, -63.4772, -63.34266, -63.20912, -63.07645, -62.94584, 
        -62.81792, -62.69261, -62.57022, -62.45073, -62.33374, -62.21923, 
        -62.10699, -61.99697, -61.88887, -61.78256, -61.67754, -61.57309, 
        -61.4688, -61.36352, -61.25532, -61.14575, -61.03318, -60.91793, 
        -60.80012, -60.68049, -60.55989, -60.43942, -60.32038, -60.20417, 
        -60.09151, -59.98389, -59.88224, -59.78705, -59.69896, -59.61843, 
        -59.54529, -59.47955, -59.4208, -59.36843, -59.32163, -59.28007, 
        -59.24285, -59.20953, -59.17923, -59.15182, -59.12642, -59.10252, 
        -59.07894, -59.05498, -59.03048, -59.00504, -58.97876, -58.95208, 
        -58.92559, -58.90028, -58.87589, -58.85273, -58.82957, -58.808, 
        -58.78702, -58.76633, -58.74579, -58.72519, -58.70429, -58.68293, 
        -58.66091, -58.63792, -58.61392, -58.58825, -58.56068, -58.53175, 
        -58.5021, -58.47302, -58.44569, -58.42108, -58.40018, -58.38367, 
        -58.37243, -58.36728, -58.36907, -58.37831, -58.395, -58.41886, 
        -58.44944,
  -47.57531, -47.78606, -47.99117, -48.19459, -48.39919, -48.60638, 
        -48.81953, -49.03897, -49.26575, -49.50034, -49.74369, -49.99612, 
        -50.2567, -50.52415, -50.79726, -51.07549, -51.35884, -51.64759, 
        -51.94199, -52.24287, -52.54883, -52.8616, -53.1804, -53.5033, 
        -53.82937, -54.15689, -54.48437, -54.8091, -55.12914, -55.44224, 
        -55.74649, -56.04036, -56.32285, -56.59234, -56.84804, -57.08887, 
        -57.31697, -57.53254, -57.73644, -57.92997, -58.11329, -58.28633, 
        -58.44852, -58.59919, -58.73818, -58.86542, -58.98144, -59.08703, 
        -59.18354, -59.27147, -59.35238, -59.42633, -59.49618, -59.56236, 
        -59.62583, -59.68764, -59.74871, -59.80975, -59.87151, -59.93439, 
        -59.99837, -60.0632, -60.12877, -60.19427, -60.25937, -60.32375, 
        -60.38794, -60.45287, -60.51842, -60.58733, -60.65911, -60.73462, 
        -60.81369, -60.89611, -60.98132, -61.06919, -61.16021, -61.25491, 
        -61.3541, -61.45861, -61.5694, -61.68689, -61.81182, -61.94428, 
        -62.08428, -62.23063, -62.38459, -62.54444, -62.70836, -62.87514, 
        -63.04324, -63.21133, -63.37742, -63.53984, -63.69644, -63.84457, 
        -63.98191, -64.10657, -64.21783, -64.31599, -64.40185, -64.47739, 
        -64.54472, -64.60582, -64.66248, -64.7183, -64.77393, -64.82963, 
        -64.885, -64.93914, -64.9912, -65.04124, -65.08887, -65.13444, 
        -65.17884, -65.22301, -65.26818, -65.31568, -65.36646, -65.4211, 
        -65.47932, -65.54111, -65.60588, -65.6727, -65.73951, -65.80791, 
        -65.87717, -65.9483, -66.02183, -66.09796, -66.17596, -66.25544, 
        -66.33585, -66.41603, -66.49512, -66.57178, -66.64532, -66.71534, 
        -66.78139, -66.84362, -66.90173, -66.95591, -67.00598, -67.0513, 
        -67.09179, -67.12579, -67.15548, -67.17982, -67.19886, -67.21292, 
        -67.22203, -67.22657, -67.22677, -67.22264, -67.21446, -67.20197, 
        -67.18569, -67.16618, -67.14377, -67.11913, -67.09229, -67.06354, 
        -67.03303, -67.00064, -66.96657, -66.93081, -66.89368, -66.85538, 
        -66.81565, -66.77358, -66.73137, -66.68849, -66.64582, -66.60356, 
        -66.5621, -66.52141, -66.48159, -66.44279, -66.40414, -66.36507, 
        -66.3247, -66.28316, -66.24032, -66.19608, -66.15047, -66.10313, 
        -66.05446, -66.00463, -65.95293, -65.8997, -65.84447, -65.78731, 
        -65.72842, -65.66737, -65.60431, -65.53764, -65.46947, -65.39907, 
        -65.32558, -65.24895, -65.1684, -65.08414, -64.99576, -64.9026, 
        -64.80531, -64.70341, -64.59724, -64.48752, -64.37418, -64.25787, 
        -64.13814, -64.01583, -63.8909, -63.76303, -63.63229, -63.4982, 
        -63.36145, -63.22273, -63.08274, -62.9429, -62.80401, -62.66729, 
        -62.53374, -62.40387, -62.27642, -62.15318, -62.03262, -61.91436, 
        -61.79818, -61.68377, -61.57092, -61.45965, -61.3495, -61.24006, 
        -61.13071, -61.02094, -60.9098, -60.7966, -60.68112, -60.56311, 
        -60.44302, -60.32131, -60.19895, -60.07702, -59.95695, -59.83999, 
        -59.72742, -59.62037, -59.51978, -59.42659, -59.34084, -59.263, 
        -59.19292, -59.13031, -59.07477, -59.02551, -58.98187, -58.94318, 
        -58.90915, -58.87813, -58.85165, -58.82819, -58.80751, -58.78899, 
        -58.77187, -58.75488, -58.73772, -58.72006, -58.70168, -58.68299, 
        -58.66433, -58.64612, -58.62847, -58.61123, -58.59407, -58.57665, 
        -58.5586, -58.53967, -58.51991, -58.49923, -58.4775, -58.45475, 
        -58.43103, -58.40626, -58.38034, -58.35295, -58.32404, -58.29402, 
        -58.26364, -58.23409, -58.2064, -58.18142, -58.16011, -58.14301, 
        -58.13103, -58.1252, -58.12634, -58.13532, -58.15244, -58.17764, 
        -58.21,
  -47.29618, -47.50649, -47.71133, -47.91388, -48.11747, -48.32487, 
        -48.53755, -48.75603, -48.98221, -49.21618, -49.45894, -49.71062, 
        -49.97124, -50.2392, -50.51182, -50.79038, -51.07393, -51.36306, 
        -51.65798, -51.96012, -52.26872, -52.58353, -52.90411, -53.2287, 
        -53.55612, -53.88489, -54.21354, -54.53973, -54.86178, -55.17747, 
        -55.48402, -55.78194, -56.06904, -56.34385, -56.60534, -56.85317, 
        -57.0873, -57.3087, -57.51795, -57.71574, -57.90263, -58.07808, 
        -58.24131, -58.3917, -58.52892, -58.65196, -58.76347, -58.86389, 
        -58.95448, -59.03679, -59.11246, -59.18276, -59.24909, -59.31252, 
        -59.37409, -59.43459, -59.49511, -59.5558, -59.61735, -59.6795, 
        -59.74239, -59.80573, -59.86796, -59.93035, -59.99141, -60.05094, 
        -60.1098, -60.16893, -60.22948, -60.29292, -60.35969, -60.43109, 
        -60.50653, -60.5861, -60.66931, -60.75559, -60.84522, -60.93903, 
        -61.03772, -61.14066, -61.2509, -61.36827, -61.49353, -61.62674, 
        -61.76822, -61.91839, -62.07631, -62.24123, -62.41217, -62.58723, 
        -62.76492, -62.94307, -63.11989, -63.29311, -63.46064, -63.61956, 
        -63.76685, -63.89956, -64.01846, -64.12259, -64.21239, -64.28961, 
        -64.35643, -64.41524, -64.46845, -64.5187, -64.56734, -64.61514, 
        -64.66239, -64.70852, -64.75362, -64.79725, -64.83955, -64.88091, 
        -64.92261, -64.96541, -65.01, -65.05677, -65.10812, -65.16419, 
        -65.22427, -65.28826, -65.35512, -65.4239, -65.49382, -65.56442, 
        -65.636, -65.70944, -65.78499, -65.86272, -65.94228, -66.02286, 
        -66.1039, -66.18427, -66.2633, -66.33983, -66.4128, -66.4822, 
        -66.54646, -66.60816, -66.66608, -66.71964, -66.76928, -66.81431, 
        -66.85458, -66.88952, -66.91888, -66.94256, -66.96064, -66.97308, 
        -66.9801, -66.98196, -66.97916, -66.97159, -66.95988, -66.94402, 
        -66.92435, -66.90181, -66.87687, -66.85026, -66.82109, -66.79121, 
        -66.75968, -66.72621, -66.69111, -66.65424, -66.61559, -66.57538, 
        -66.53375, -66.49122, -66.44788, -66.4044, -66.36157, -66.31953, 
        -66.27909, -66.23993, -66.20182, -66.16454, -66.12775, -66.09085, 
        -66.05286, -66.01353, -65.97283, -65.93069, -65.88725, -65.84153, 
        -65.79527, -65.74734, -65.69743, -65.64594, -65.59293, -65.53769, 
        -65.48051, -65.42097, -65.35957, -65.29568, -65.22868, -65.15918, 
        -65.08639, -65.01035, -64.93013, -64.84524, -64.75597, -64.66151, 
        -64.56201, -64.45792, -64.34915, -64.23655, -64.12008, -64.00089, 
        -63.87891, -63.754, -63.62658, -63.49479, -63.36105, -63.22353, 
        -63.08249, -62.93908, -62.79406, -62.64904, -62.50489, -62.36335, 
        -62.22527, -62.09142, -61.96189, -61.83601, -61.71281, -61.59188, 
        -61.47275, -61.35511, -61.23872, -61.12326, -61.00871, -60.89495, 
        -60.78149, -60.66772, -60.55296, -60.43661, -60.31854, -60.19823, 
        -60.07607, -59.9528, -59.82919, -59.70631, -59.5856, -59.46847, 
        -59.35536, -59.24932, -59.15027, -59.05891, -58.9758, -58.90063, 
        -58.83321, -58.7733, -58.72017, -58.67318, -58.6318, -58.59552, 
        -58.56366, -58.53619, -58.51289, -58.49314, -58.47667, -58.46302, 
        -58.45148, -58.44123, -58.43108, -58.42079, -58.41032, -58.39953, 
        -58.38872, -58.37778, -58.36679, -58.35557, -58.34362, -58.33027, 
        -58.31517, -58.29824, -58.27937, -58.25865, -58.23632, -58.21242, 
        -58.18726, -58.16086, -58.13347, -58.10498, -58.07509, -58.0445, 
        -58.0126, -57.98277, -57.95457, -57.92889, -57.90657, -57.88821, 
        -57.87477, -57.86741, -57.8671, -57.87495, -57.89161, -57.91702, 
        -57.95072,
  -47.01013, -47.21933, -47.42332, -47.62506, -47.82748, -48.03363, 
        -48.2452, -48.46274, -48.68792, -48.92014, -49.16217, -49.41323, 
        -49.67392, -49.9421, -50.21619, -50.49544, -50.77983, -51.07004, 
        -51.3667, -51.67053, -51.98153, -52.29911, -52.62204, -52.94852, 
        -53.2761, -53.60526, -53.93404, -54.26053, -54.58327, -54.90041, 
        -55.21018, -55.51097, -55.8018, -56.08101, -56.34731, -56.6008, 
        -56.84079, -57.06751, -57.28153, -57.48296, -57.67115, -57.84756, 
        -58.01035, -58.15892, -58.29282, -58.41272, -58.51959, -58.61413, 
        -58.69886, -58.77571, -58.84643, -58.91312, -58.97684, -59.03887, 
        -59.10018, -59.16117, -59.22152, -59.28316, -59.34511, -59.4074, 
        -59.46965, -59.53163, -59.59244, -59.65145, -59.70824, -59.76291, 
        -59.81613, -59.86926, -59.9239, -59.9814, -60.04303, -60.1098, 
        -60.18154, -60.2567, -60.3373, -60.42126, -60.50935, -60.60245, 
        -60.70002, -60.80278, -60.91199, -61.02861, -61.15348, -61.28693, 
        -61.43005, -61.58264, -61.74454, -61.91472, -62.0924, -62.27562, 
        -62.46241, -62.65012, -62.83782, -63.02242, -63.20125, -63.37125, 
        -63.52953, -63.673, -63.80036, -63.91082, -64.00487, -64.08421, 
        -64.15045, -64.20681, -64.25562, -64.29998, -64.34175, -64.38162, 
        -64.42065, -64.45911, -64.49585, -64.53333, -64.57037, -64.60809, 
        -64.64713, -64.6884, -64.73278, -64.78122, -64.83405, -64.89159, 
        -64.95356, -65.01978, -65.08845, -65.15907, -65.23096, -65.30407, 
        -65.37867, -65.45442, -65.5318, -65.61091, -65.69068, -65.77245, 
        -65.85393, -65.93449, -66.01315, -66.08913, -66.16179, -66.2304, 
        -66.29523, -66.35619, -66.41364, -66.46732, -66.51662, -66.56152, 
        -66.60166, -66.6365, -66.66574, -66.68867, -66.70524, -66.7156, 
        -66.72026, -66.7193, -66.71188, -66.70056, -66.68462, -66.66476, 
        -66.64165, -66.6157, -66.58797, -66.55896, -66.52899, -66.49784, 
        -66.46495, -66.4304, -66.39377, -66.35532, -66.315, -66.27267, 
        -66.22914, -66.18471, -66.14022, -66.09633, -66.05321, -66.01168, 
        -65.97207, -65.93438, -65.89732, -65.86166, -65.82657, -65.79136, 
        -65.75562, -65.71905, -65.68027, -65.64001, -65.59887, -65.55662, 
        -65.51314, -65.46709, -65.41934, -65.36967, -65.31804, -65.26493, 
        -65.20884, -65.15062, -65.08993, -65.0269, -64.9614, -64.8923, 
        -64.81995, -64.74368, -64.66359, -64.57875, -64.48798, -64.39113, 
        -64.28982, -64.18317, -64.07209, -63.95639, -63.83698, -63.71443, 
        -63.58944, -63.46239, -63.33169, -63.19781, -63.06017, -62.91904, 
        -62.77438, -62.62645, -62.47723, -62.3278, -62.17987, -62.03473, 
        -61.89346, -61.7569, -61.62505, -61.49716, -61.37247, -61.24974, 
        -61.12879, -61.00884, -60.88974, -60.77143, -60.65362, -60.53625, 
        -60.41849, -60.30136, -60.18364, -60.06474, -59.94434, -59.82222, 
        -59.69868, -59.57399, -59.44947, -59.32629, -59.2056, -59.08906, 
        -58.97779, -58.87325, -58.7761, -58.68697, -58.60618, -58.53371, 
        -58.46893, -58.41136, -58.3602, -58.31511, -58.27531, -58.24054, 
        -58.21059, -58.18506, -58.16416, -58.14754, -58.13484, -58.12547, 
        -58.1189, -58.11444, -58.11083, -58.10765, -58.10441, -58.10125, 
        -58.09768, -58.0928, -58.08832, -58.08294, -58.07593, -58.0667, 
        -58.05479, -58.03995, -58.02244, -58.00229, -57.9798, -57.9553, 
        -57.92909, -57.90165, -57.87314, -57.84385, -57.81363, -57.78262, 
        -57.75167, -57.72116, -57.69228, -57.66554, -57.64163, -57.62136, 
        -57.60575, -57.59613, -57.59364, -57.59951, -57.61477, -57.63961, 
        -57.67401,
  -46.71384, -46.92197, -47.12467, -47.32553, -47.52581, -47.73048, 
        -47.94048, -48.15678, -48.3806, -48.61302, -48.85458, -49.10559, 
        -49.3662, -49.63493, -49.91021, -50.191, -50.47747, -50.77015, 
        -51.06978, -51.37556, -51.68989, -52.01075, -52.33623, -52.66455, 
        -52.99349, -53.32204, -53.64994, -53.97543, -54.29753, -54.61451, 
        -54.92484, -55.22719, -55.52043, -55.80315, -56.07235, -56.33061, 
        -56.57555, -56.80693, -57.02463, -57.2285, -57.41851, -57.59423, 
        -57.75491, -57.90004, -58.02974, -58.14451, -58.24529, -58.33435, 
        -58.41351, -58.48533, -58.55125, -58.6152, -58.6778, -58.74018, 
        -58.80261, -58.86571, -58.92916, -58.99257, -59.05572, -59.11859, 
        -59.18057, -59.24115, -59.29928, -59.35499, -59.40755, -59.45722, 
        -59.50472, -59.55073, -59.5994, -59.65129, -59.70778, -59.7698, 
        -59.83741, -59.91014, -59.9873, -60.06917, -60.15519, -60.24707, 
        -60.34291, -60.44386, -60.55164, -60.66682, -60.79088, -60.92493, 
        -61.06847, -61.22368, -61.38956, -61.5653, -61.74964, -61.94091, 
        -62.13695, -62.33577, -62.53468, -62.73095, -62.9216, -63.10325, 
        -63.27266, -63.42633, -63.56242, -63.67977, -63.77843, -63.85959, 
        -63.92555, -63.97847, -64.02325, -64.06179, -64.09642, -64.12874, 
        -64.15985, -64.19033, -64.22104, -64.25223, -64.28455, -64.3187, 
        -64.35543, -64.39558, -64.4401, -64.48936, -64.54382, -64.60313, 
        -64.66711, -64.73491, -64.80526, -64.87663, -64.9509, -65.02657, 
        -65.10358, -65.18159, -65.261, -65.34156, -65.42344, -65.50576, 
        -65.58754, -65.66815, -65.74646, -65.82201, -65.89398, -65.96211, 
        -66.02669, -66.08739, -66.14464, -66.19807, -66.24738, -66.29245, 
        -66.33154, -66.36625, -66.39495, -66.41674, -66.43173, -66.43993, 
        -66.44166, -66.43714, -66.42676, -66.41119, -66.39098, -66.36695, 
        -66.33986, -66.31049, -66.27982, -66.24825, -66.21614, -66.18313, 
        -66.14866, -66.11246, -66.07406, -66.03352, -65.99092, -65.94534, 
        -65.89957, -65.85332, -65.80753, -65.76271, -65.71962, -65.67881, 
        -65.64021, -65.60401, -65.56937, -65.5356, -65.50233, -65.46876, 
        -65.43496, -65.40014, -65.36362, -65.32588, -65.28687, -65.24694, 
        -65.20559, -65.16211, -65.11673, -65.06881, -65.01871, -64.96623, 
        -64.91103, -64.85262, -64.79247, -64.72995, -64.66441, -64.59567, 
        -64.52364, -64.44753, -64.36696, -64.28124, -64.18964, -64.09227, 
        -63.98894, -63.88024, -63.76623, -63.64761, -63.52526, -63.39972, 
        -63.27159, -63.14085, -63.00687, -62.86957, -62.72818, -62.5829, 
        -62.4341, -62.28244, -62.12957, -61.97714, -61.82673, -61.67948, 
        -61.53546, -61.39746, -61.26424, -61.13541, -61.00987, -60.88637, 
        -60.76427, -60.64296, -60.52235, -60.40216, -60.28208, -60.1624, 
        -60.04294, -59.92334, -59.8032, -59.68213, -59.55993, -59.43635, 
        -59.31157, -59.18625, -59.06144, -58.93848, -58.81874, -58.70338, 
        -58.59378, -58.49108, -58.39609, -58.30948, -58.2313, -58.16144, 
        -58.09924, -58.04386, -57.99457, -57.951, -57.91257, -57.87817, 
        -57.84958, -57.82568, -57.80674, -57.79262, -57.78313, -57.77755, 
        -57.77533, -57.77551, -57.77747, -57.78056, -57.78392, -57.78737, 
        -57.79038, -57.79314, -57.79472, -57.79481, -57.79271, -57.78746, 
        -57.77899, -57.76682, -57.75113, -57.73215, -57.71009, -57.68561, 
        -57.65905, -57.6311, -57.60211, -57.57261, -57.54224, -57.511, 
        -57.47969, -57.44886, -57.41891, -57.39059, -57.36469, -57.34206, 
        -57.32376, -57.31113, -57.30566, -57.30882, -57.32184, -57.34543, 
        -57.37984,
  -46.40575, -46.61203, -46.81324, -47.0125, -47.2126, -47.41543, 
        -47.62354, -47.83846, -48.06113, -48.29254, -48.5338, -48.78497, 
        -49.04597, -49.31636, -49.59268, -49.87635, -50.16647, -50.46331, 
        -50.76742, -51.07878, -51.39658, -51.72045, -52.0481, -52.3774, 
        -52.70589, -53.03327, -53.35935, -53.68282, -54.00275, -54.31749, 
        -54.62749, -54.93048, -55.22503, -55.51009, -55.78357, -56.04535, 
        -56.29387, -56.52811, -56.74768, -56.95205, -57.1411, -57.31418, 
        -57.47128, -57.61157, -57.73483, -57.8438, -57.93906, -58.02251, 
        -58.09681, -58.16492, -58.22933, -58.29234, -58.35526, -58.41919, 
        -58.48428, -58.55036, -58.6166, -58.68245, -58.74739, -58.81105, 
        -58.87285, -58.93092, -58.98703, -59.03932, -59.08784, -59.13277, 
        -59.1749, -59.21606, -59.25893, -59.30514, -59.35654, -59.41358, 
        -59.47602, -59.54454, -59.61874, -59.69759, -59.78192, -59.87075, 
        -59.96399, -60.06293, -60.16895, -60.28278, -60.40644, -60.54106, 
        -60.68744, -60.84563, -61.01589, -61.19734, -61.38853, -61.58781, 
        -61.79317, -62.00231, -62.21242, -62.42043, -62.62288, -62.81604, 
        -62.9955, -63.15934, -63.30423, -63.42842, -63.53177, -63.61517, 
        -63.68132, -63.73349, -63.77428, -63.80716, -63.83485, -63.85965, 
        -63.88291, -63.90578, -63.92972, -63.95506, -63.98272, -64.01362, 
        -64.04835, -64.08809, -64.13178, -64.18195, -64.23772, -64.29884, 
        -64.3644, -64.43346, -64.50523, -64.57973, -64.65622, -64.73418, 
        -64.81297, -64.89301, -64.97417, -65.05623, -65.13905, -65.22162, 
        -65.30357, -65.38413, -65.4622, -65.53738, -65.60789, -65.67573, 
        -65.74023, -65.80105, -65.85836, -65.9119, -65.96128, -66.00641, 
        -66.04653, -66.08079, -66.10851, -66.12899, -66.14216, -66.1478, 
        -66.14629, -66.13795, -66.12341, -66.10326, -66.07868, -66.0504, 
        -66.01911, -65.98602, -65.9522, -65.9168, -65.88217, -65.84665, 
        -65.80998, -65.77162, -65.73089, -65.68771, -65.64229, -65.59507, 
        -65.5471, -65.49901, -65.45177, -65.4062, -65.36308, -65.32294, 
        -65.28563, -65.25079, -65.21755, -65.1853, -65.15376, -65.12198, 
        -65.08968, -65.05631, -65.02172, -64.98553, -64.94901, -64.91151, 
        -64.87224, -64.83124, -64.78815, -64.74202, -64.69318, -64.64097, 
        -64.58614, -64.52875, -64.46858, -64.40599, -64.34022, -64.27145, 
        -64.19942, -64.12315, -64.04224, -63.95542, -63.86267, -63.76381, 
        -63.65843, -63.5473, -63.43061, -63.30905, -63.18372, -63.05519, 
        -62.92369, -62.78794, -62.6501, -62.50874, -62.36318, -62.21394, 
        -62.061, -61.90587, -61.7503, -61.59575, -61.44397, -61.29602, 
        -61.15273, -61.01466, -60.88161, -60.75273, -60.62701, -60.50347, 
        -60.38114, -60.25927, -60.13779, -60.01645, -59.89524, -59.77411, 
        -59.65295, -59.5317, -59.40992, -59.28736, -59.16373, -59.03915, 
        -58.91377, -58.78834, -58.66407, -58.54203, -58.42268, -58.30922, 
        -58.20185, -58.10176, -58.00962, -57.92586, -57.85059, -57.78333, 
        -57.72362, -57.67055, -57.62326, -57.58118, -57.54407, -57.51179, 
        -57.48449, -57.46207, -57.44478, -57.43263, -57.42545, -57.42267, 
        -57.42365, -57.42751, -57.43394, -57.44181, -57.45082, -57.45996, 
        -57.46914, -57.47747, -57.48474, -57.49017, -57.49278, -57.4919, 
        -57.48704, -57.47788, -57.46452, -57.44722, -57.4263, -57.40231, 
        -57.376, -57.34817, -57.31924, -57.28874, -57.2585, -57.22756, 
        -57.19608, -57.1645, -57.13338, -57.10332, -57.07516, -57.04985, 
        -57.02837, -57.01231, -57.0032, -57.00314, -57.01358, -57.0358, 
        -57.07011,
  -46.08604, -46.29021, -46.49014, -46.68768, -46.88622, -47.08731, 
        -47.29377, -47.5068, -47.72713, -47.9577, -48.19867, -48.45037, 
        -48.71279, -48.98513, -49.26616, -49.55453, -49.85008, -50.15266, 
        -50.46208, -50.77848, -51.10085, -51.42721, -51.75639, -52.08428, 
        -52.41174, -52.73702, -53.06037, -53.38065, -53.69784, -54.01147, 
        -54.32013, -54.62263, -54.91793, -55.20418, -55.47958, -55.74314, 
        -55.99359, -56.22906, -56.44858, -56.65067, -56.83682, -57.00609, 
        -57.15804, -57.2927, -57.41097, -57.51375, -57.6033, -57.68178, 
        -57.7523, -57.81796, -57.88125, -57.94441, -58.00908, -58.07584, 
        -58.14452, -58.21343, -58.28325, -58.3522, -58.41909, -58.48391, 
        -58.54574, -58.60368, -58.65764, -58.70701, -58.75179, -58.7922, 
        -58.82943, -58.86567, -58.90332, -58.94417, -58.98984, -59.0415, 
        -59.09797, -59.16206, -59.23212, -59.3084, -59.38913, -59.47549, 
        -59.56713, -59.66358, -59.76735, -59.88009, -60.00383, -60.13972, 
        -60.28819, -60.45029, -60.62551, -60.81265, -61.01102, -61.21849, 
        -61.43214, -61.65148, -61.87276, -62.09231, -62.30635, -62.51061, 
        -62.70168, -62.87529, -63.02844, -63.15946, -63.26764, -63.35387, 
        -63.42069, -63.47112, -63.50863, -63.53641, -63.55764, -63.57491, 
        -63.59071, -63.60546, -63.623, -63.64284, -63.66602, -63.69381, 
        -63.72688, -63.76624, -63.81102, -63.86166, -63.91868, -63.98125, 
        -64.04816, -64.1184, -64.19161, -64.26736, -64.34551, -64.42542, 
        -64.506, -64.58751, -64.67002, -64.75218, -64.83584, -64.91885, 
        -65.00095, -65.08119, -65.15917, -65.23415, -65.30562, -65.37357, 
        -65.43813, -65.49939, -65.55721, -65.61102, -65.66061, -65.70566, 
        -65.74542, -65.77906, -65.80551, -65.82424, -65.83489, -65.83749, 
        -65.83245, -65.81901, -65.79999, -65.7752, -65.7458, -65.71293, 
        -65.67732, -65.64046, -65.60302, -65.56551, -65.52794, -65.4895, 
        -65.45, -65.40871, -65.36506, -65.319, -65.27043, -65.22044, 
        -65.16978, -65.11973, -65.07143, -65.02512, -64.98204, -64.9425, 
        -64.90558, -64.87241, -64.8406, -64.81007, -64.77977, -64.74931, 
        -64.71889, -64.68693, -64.65457, -64.62141, -64.58722, -64.55255, 
        -64.51546, -64.47659, -64.43523, -64.39089, -64.34341, -64.29137, 
        -64.23645, -64.17821, -64.11761, -64.05473, -63.98839, -63.91929, 
        -63.84663, -63.76991, -63.68863, -63.59994, -63.50571, -63.40483, 
        -63.29758, -63.18418, -63.06469, -62.9407, -62.81217, -62.68023, 
        -62.54533, -62.40656, -62.26434, -62.11812, -61.96829, -61.81486, 
        -61.65814, -61.49995, -61.34213, -61.18657, -61.03454, -60.8871, 
        -60.7451, -60.60816, -60.4761, -60.34817, -60.22307, -60.10009, 
        -59.97832, -59.85665, -59.73497, -59.61249, -59.49094, -59.36932, 
        -59.24767, -59.12564, -59.00317, -58.87975, -58.75537, -58.63031, 
        -58.50489, -58.38006, -58.25689, -58.13657, -58.02013, -57.90919, 
        -57.8049, -57.7081, -57.6192, -57.53873, -57.46662, -57.40228, 
        -57.3451, -57.29427, -57.24906, -57.20873, -57.17312, -57.14201, 
        -57.11588, -57.09493, -57.07907, -57.06874, -57.06324, -57.0624, 
        -57.06589, -57.07255, -57.08184, -57.09335, -57.10659, -57.11946, 
        -57.13319, -57.14639, -57.1585, -57.16859, -57.17578, -57.17926, 
        -57.1782, -57.17237, -57.16188, -57.14679, -57.12768, -57.10515, 
        -57.07976, -57.05256, -57.02431, -56.99532, -56.96554, -56.93504, 
        -56.9035, -56.87135, -56.83913, -56.80728, -56.77679, -56.7487, 
        -56.72375, -56.70401, -56.69086, -56.6869, -56.69442, -56.71484, 
        -56.74889,
  -45.75558, -45.95703, -46.15438, -46.34908, -46.54558, -46.74547, 
        -46.95033, -47.1621, -47.38248, -47.61257, -47.85336, -48.10582, 
        -48.37058, -48.6456, -48.93092, -49.22475, -49.5264, -49.83548, 
        -50.15022, -50.47177, -50.79753, -51.12625, -51.45565, -51.78378, 
        -52.10956, -52.43234, -52.75213, -53.06895, -53.38305, -53.69384, 
        -54.00094, -54.30276, -54.59795, -54.88377, -55.16018, -55.4242, 
        -55.67408, -55.90825, -56.12567, -56.32544, -56.50731, -56.6711, 
        -56.81732, -56.94597, -57.05797, -57.15516, -57.23958, -57.31424, 
        -57.38198, -57.44522, -57.50868, -57.57342, -57.64102, -57.71154, 
        -57.78427, -57.85824, -57.93199, -58.00405, -58.07353, -58.13941, 
        -58.20136, -58.25878, -58.31094, -58.35799, -58.39953, -58.43641, 
        -58.46896, -58.50095, -58.53418, -58.56955, -58.60976, -58.65582, 
        -58.708, -58.76715, -58.83286, -58.9043, -58.98161, -59.06472, 
        -59.15277, -59.247, -59.34942, -59.46129, -59.58558, -59.72193, 
        -59.87428, -60.04074, -60.22142, -60.41492, -60.6208, -60.83669, 
        -61.06063, -61.29018, -61.52219, -61.75232, -61.97691, -62.1916, 
        -62.39215, -62.57464, -62.73553, -62.87288, -62.98593, -63.07502, 
        -63.14198, -63.19132, -63.22585, -63.24911, -63.26439, -63.2753, 
        -63.28437, -63.29333, -63.30462, -63.31921, -63.3385, -63.36337, 
        -63.39494, -63.43283, -63.47749, -63.52868, -63.58653, -63.64991, 
        -63.71774, -63.78794, -63.86241, -63.93953, -64.01832, -64.09915, 
        -64.18099, -64.2638, -64.3474, -64.4313, -64.51537, -64.59863, 
        -64.68077, -64.7612, -64.83913, -64.91418, -64.98585, -65.05437, 
        -65.1198, -65.1818, -65.24017, -65.29444, -65.34417, -65.38795, 
        -65.42696, -65.4596, -65.48428, -65.50076, -65.50856, -65.50782, 
        -65.4988, -65.48183, -65.45804, -65.42829, -65.39383, -65.35606, 
        -65.31608, -65.27511, -65.23389, -65.19273, -65.15149, -65.10947, 
        -65.06645, -65.02163, -64.97452, -64.92483, -64.87207, -64.81918, 
        -64.7661, -64.71415, -64.66457, -64.6178, -64.57504, -64.53654, 
        -64.50172, -64.46988, -64.4396, -64.41035, -64.38186, -64.35264, 
        -64.32328, -64.29314, -64.26268, -64.23206, -64.20078, -64.16837, 
        -64.13361, -64.09669, -64.05746, -64.01437, -63.96736, -63.91486, 
        -63.8594, -63.801, -63.73954, -63.67572, -63.60841, -63.53867, 
        -63.46582, -63.38849, -63.3061, -63.21721, -63.1218, -63.01951, 
        -62.91021, -62.79441, -62.67229, -62.54538, -62.41435, -62.27913, 
        -62.14012, -61.99686, -61.84997, -61.69912, -61.54459, -61.38691, 
        -61.22658, -61.06601, -60.90683, -60.7509, -60.59859, -60.45254, 
        -60.31246, -60.17786, -60.04779, -59.9215, -59.79794, -59.67635, 
        -59.55565, -59.43517, -59.31426, -59.19333, -59.07228, -58.95119, 
        -58.82973, -58.70795, -58.58551, -58.46227, -58.33789, -58.21276, 
        -58.08793, -57.96443, -57.84324, -57.72537, -57.61193, -57.50431, 
        -57.40356, -57.31057, -57.22547, -57.14858, -57.07966, -57.01827, 
        -56.96355, -56.91483, -56.8705, -56.83181, -56.79781, -56.76825, 
        -56.74358, -56.7238, -56.7097, -56.70066, -56.69663, -56.69699, 
        -56.7016, -56.70995, -56.72144, -56.73558, -56.75163, -56.76876, 
        -56.78627, -56.8035, -56.8197, -56.83394, -56.84523, -56.85279, 
        -56.85569, -56.85332, -56.84579, -56.83335, -56.81639, -56.79559, 
        -56.77211, -56.74642, -56.71937, -56.69144, -56.66262, -56.63292, 
        -56.60184, -56.56933, -56.53598, -56.50243, -56.46977, -56.43895, 
        -56.41057, -56.38697, -56.36984, -56.36222, -56.36666, -56.38398, 
        -56.41806,
  -45.41492, -45.61291, -45.80737, -46.0008, -46.19555, -46.39414, 
        -46.59835, -46.80949, -47.02943, -47.25943, -47.50115, -47.75464, 
        -48.02121, -48.29892, -48.58841, -48.88772, -49.19576, -49.51134, 
        -49.83282, -50.15887, -50.4874, -50.81647, -51.14486, -51.47129, 
        -51.79448, -52.11406, -52.43018, -52.74359, -53.05342, -53.36203, 
        -53.66743, -53.9684, -54.26327, -54.5501, -54.82598, -55.0885, 
        -55.33603, -55.56696, -55.78009, -55.97511, -56.15131, -56.30914, 
        -56.44924, -56.57099, -56.67757, -56.77003, -56.8508, -56.92271, 
        -56.989, -57.05285, -57.11742, -57.18463, -57.25566, -57.33022, 
        -57.40731, -57.48567, -57.56335, -57.63882, -57.71069, -57.77813, 
        -57.8395, -57.89659, -57.94779, -57.99302, -58.03242, -58.06709, 
        -58.09814, -58.12723, -58.15607, -58.18727, -58.22219, -58.26266, 
        -58.30948, -58.36346, -58.4242, -58.49104, -58.56409, -58.64197, 
        -58.72673, -58.81845, -58.91937, -59.03112, -59.15602, -59.29659, 
        -59.45261, -59.62434, -59.81075, -60.01156, -60.22529, -60.44965, 
        -60.68238, -60.92156, -61.1629, -61.40268, -61.63652, -61.85911, 
        -62.0679, -62.25798, -62.42563, -62.56865, -62.68625, -62.77843, 
        -62.84751, -62.89639, -62.92889, -62.94863, -62.95943, -62.96453, 
        -62.96746, -62.9705, -62.97619, -62.9861, -63.00172, -63.02382, 
        -63.05165, -63.08786, -63.13166, -63.18277, -63.24087, -63.30442, 
        -63.37289, -63.44487, -63.52002, -63.59743, -63.67671, -63.75793, 
        -63.84038, -63.92383, -64.00787, -64.0921, -64.17641, -64.25977, 
        -64.34191, -64.42233, -64.50052, -64.57526, -64.64776, -64.71728, 
        -64.78372, -64.84675, -64.90632, -64.96108, -65.01109, -65.05546, 
        -65.09355, -65.12453, -65.14688, -65.16065, -65.16518, -65.16051, 
        -65.14712, -65.12538, -65.09637, -65.06133, -65.0215, -64.97852, 
        -64.93359, -64.88699, -64.84129, -64.79595, -64.75051, -64.70441, 
        -64.65712, -64.60799, -64.5567, -64.50331, -64.44809, -64.39223, 
        -64.33672, -64.28319, -64.23278, -64.18589, -64.14364, -64.10582, 
        -64.07218, -64.04176, -64.01286, -63.98521, -63.9577, -63.9302, 
        -63.90261, -63.8746, -63.84556, -63.81732, -63.78865, -63.75891, 
        -63.72653, -63.69154, -63.6533, -63.61123, -63.56517, -63.51373, 
        -63.4584, -63.39921, -63.33684, -63.27243, -63.20456, -63.13406, 
        -63.06033, -62.9823, -62.8991, -62.80907, -62.7124, -62.60845, 
        -62.49726, -62.37949, -62.25511, -62.12536, -61.99099, -61.85162, 
        -61.70856, -61.56098, -61.40923, -61.25341, -61.09416, -60.93241, 
        -60.76934, -60.60673, -60.44669, -60.29114, -60.14119, -59.99725, 
        -59.85962, -59.7277, -59.60062, -59.47702, -59.35574, -59.23608, 
        -59.11717, -58.99829, -58.87917, -58.75963, -58.63987, -58.52018, 
        -58.40015, -58.27935, -58.15769, -58.03505, -57.91162, -57.78766, 
        -57.66443, -57.54185, -57.42339, -57.30882, -57.19926, -57.09572, 
        -56.99911, -56.91012, -56.8289, -56.75558, -56.68961, -56.63069, 
        -56.57814, -56.53122, -56.48959, -56.45262, -56.42032, -56.39251, 
        -56.3693, -56.35107, -56.33809, -56.33032, -56.32722, -56.32834, 
        -56.33359, -56.34292, -56.35587, -56.37166, -56.38956, -56.40903, 
        -56.42947, -56.4501, -56.46976, -56.48761, -56.50262, -56.51384, 
        -56.52027, -56.5211, -56.51645, -56.50638, -56.49201, -56.47386, 
        -56.45174, -56.42799, -56.40279, -56.37665, -56.34951, -56.32103, 
        -56.29065, -56.25836, -56.22429, -56.18948, -56.15485, -56.12139, 
        -56.09014, -56.06307, -56.04245, -56.03149, -56.03341, -56.05021, 
        -56.08374,
  -45.069, -45.26339, -45.45475, -45.64578, -45.83921, -46.03684, 
        -46.24105, -46.45139, -46.6723, -46.90332, -47.14595, -47.40117, 
        -47.66996, -47.95042, -48.24408, -48.54789, -48.86074, -49.18127, 
        -49.50719, -49.83609, -50.16518, -50.49319, -50.8186, -51.14236, 
        -51.46229, -51.77792, -52.09076, -52.40105, -52.70928, -53.01561, 
        -53.3197, -53.62008, -53.91402, -54.1996, -54.47413, -54.73367, 
        -54.9772, -55.20319, -55.40971, -55.59873, -55.76905, -55.92057, 
        -56.05484, -56.17262, -56.27507, -56.36427, -56.44279, -56.51339, 
        -56.5793, -56.64399, -56.71041, -56.78054, -56.85508, -56.93384, 
        -57.01425, -57.09673, -57.17833, -57.25698, -57.33131, -57.4005, 
        -57.46394, -57.52131, -57.57219, -57.61684, -57.65536, -57.68895, 
        -57.71877, -57.74589, -57.7722, -57.79964, -57.83043, -57.8652, 
        -57.90754, -57.95652, -58.01181, -58.07396, -58.14265, -58.21727, 
        -58.29818, -58.38748, -58.48664, -58.5987, -58.72539, -58.86883, 
        -59.02918, -59.20638, -59.39967, -59.60694, -59.82863, -60.05981, 
        -60.30124, -60.54832, -60.79781, -61.04543, -61.28678, -61.51748, 
        -61.73309, -61.92919, -62.10244, -62.25017, -62.37164, -62.46675, 
        -62.53724, -62.58619, -62.61747, -62.63464, -62.64168, -62.64161, 
        -62.63982, -62.6381, -62.63913, -62.64483, -62.65654, -62.67503, 
        -62.70097, -62.73501, -62.77707, -62.82729, -62.8846, -62.94798, 
        -63.01635, -63.08853, -63.16361, -63.2409, -63.32014, -63.40105, 
        -63.48329, -63.56572, -63.64973, -63.73383, -63.81765, -63.90069, 
        -63.98288, -64.06374, -64.14262, -64.21938, -64.29319, -64.36427, 
        -64.43237, -64.49693, -64.55744, -64.61292, -64.66315, -64.70718, 
        -64.74419, -64.77316, -64.79288, -64.80328, -64.80389, -64.79374, 
        -64.77549, -64.74834, -64.71371, -64.67282, -64.62719, -64.57841, 
        -64.52802, -64.47719, -64.42666, -64.37627, -64.32591, -64.27492, 
        -64.22273, -64.16901, -64.11326, -64.05582, -63.99712, -63.93837, 
        -63.88092, -63.82604, -63.77481, -63.7277, -63.68581, -63.64812, 
        -63.61561, -63.58645, -63.55887, -63.53263, -63.50678, -63.48109, 
        -63.45563, -63.42995, -63.40483, -63.37972, -63.35391, -63.32668, 
        -63.29636, -63.26321, -63.2263, -63.18507, -63.13925, -63.08792, 
        -63.03248, -62.97347, -62.91093, -62.84569, -62.77715, -62.70602, 
        -62.63174, -62.55198, -62.46771, -62.37663, -62.27867, -62.17355, 
        -62.06096, -61.94109, -61.81445, -61.68225, -61.545, -61.40306, 
        -61.25626, -61.1041, -60.94759, -60.78722, -60.62363, -60.45801, 
        -60.29225, -60.12833, -59.96837, -59.81361, -59.66528, -59.52398, 
        -59.38946, -59.26066, -59.13681, -59.01641, -58.89808, -58.78096, 
        -58.66437, -58.54668, -58.43003, -58.31308, -58.19561, -58.07791, 
        -57.95996, -57.84108, -57.7211, -57.60016, -57.47837, -57.35644, 
        -57.23565, -57.11703, -57.00209, -56.89175, -56.78671, -56.68777, 
        -56.59578, -56.51085, -56.43329, -56.36297, -56.29967, -56.24269, 
        -56.19186, -56.1462, -56.10592, -56.07048, -56.03991, -56.01378, 
        -55.99239, -55.9756, -55.96382, -55.95681, -55.95417, -55.95575, 
        -55.96124, -55.97081, -55.98354, -56.00048, -56.01991, -56.04124, 
        -56.06407, -56.08747, -56.11021, -56.13129, -56.14948, -56.16372, 
        -56.17304, -56.17667, -56.17482, -56.16754, -56.15571, -56.14005, 
        -56.12144, -56.10034, -56.0775, -56.05363, -56.0285, -56.00198, 
        -55.97281, -55.94114, -55.90693, -55.87141, -55.83556, -55.80013, 
        -55.76682, -55.73729, -55.7142, -55.70092, -55.70082, -55.71658, 
        -55.74993,
  -44.72046, -44.91133, -45.09846, -45.28723, -45.47966, -45.67727, 
        -45.88198, -46.0949, -46.31754, -46.55042, -46.79498, -47.05212, 
        -47.32238, -47.60482, -47.90004, -48.20612, -48.52179, -48.84352, 
        -49.17094, -49.5003, -49.82824, -50.15309, -50.47558, -50.79578, 
        -51.11188, -51.42403, -51.73351, -52.04089, -52.3467, -52.65123, 
        -52.95417, -53.25342, -53.54567, -53.82921, -54.10057, -54.35647, 
        -54.59497, -54.8153, -55.01697, -55.19978, -55.36418, -55.51038, 
        -55.63975, -55.75344, -55.85341, -55.94103, -56.01879, -56.08933, 
        -56.1551, -56.22129, -56.28993, -56.36295, -56.44093, -56.5237, 
        -56.60926, -56.69577, -56.78076, -56.86235, -56.93921, -57.01041, 
        -57.07553, -57.13404, -57.18594, -57.231, -57.27028, -57.30339, 
        -57.33324, -57.35978, -57.38477, -57.4104, -57.43885, -57.47166, 
        -57.51003, -57.55485, -57.60621, -57.66404, -57.72793, -57.79839, 
        -57.87586, -57.9623, -58.06032, -58.17253, -58.29962, -58.44551, 
        -58.60986, -58.79224, -58.99151, -59.20613, -59.43495, -59.67454, 
        -59.92291, -60.17626, -60.4319, -60.68559, -60.93237, -61.16811, 
        -61.3882, -61.58871, -61.76611, -61.91751, -62.0421, -62.13859, 
        -62.2104, -62.25993, -62.29072, -62.30663, -62.31166, -62.30981, 
        -62.30473, -62.29965, -62.29701, -62.299, -62.30671, -62.32121, 
        -62.34369, -62.37469, -62.41435, -62.46239, -62.51803, -62.58036, 
        -62.64699, -62.71864, -62.79313, -62.8697, -62.94801, -63.02794, 
        -63.10942, -63.19195, -63.2751, -63.3584, -63.44139, -63.52436, 
        -63.60654, -63.6879, -63.76778, -63.84583, -63.92161, -63.99473, 
        -64.06489, -64.13127, -64.19297, -64.24863, -64.29903, -64.34266, 
        -64.37833, -64.40482, -64.4217, -64.42821, -64.42419, -64.40993, 
        -64.38581, -64.35275, -64.3119, -64.26456, -64.21262, -64.1575, 
        -64.10132, -64.04452, -63.98816, -63.93217, -63.87624, -63.81993, 
        -63.76251, -63.70373, -63.64233, -63.58053, -63.51848, -63.45706, 
        -63.39753, -63.3413, -63.28934, -63.24246, -63.20097, -63.16495, 
        -63.13351, -63.10534, -63.07942, -63.05482, -63.03085, -63.00747, 
        -62.98457, -62.9624, -62.94061, -62.91893, -62.89635, -62.87158, 
        -62.84383, -62.81212, -62.77619, -62.73559, -62.68865, -62.63801, 
        -62.58279, -62.52396, -62.4616, -62.39594, -62.32734, -62.25574, 
        -62.1808, -62.10122, -62.01591, -61.92421, -61.82517, -61.71878, 
        -61.60501, -61.48369, -61.3554, -61.22106, -61.08125, -60.93599, 
        -60.7854, -60.62967, -60.46887, -60.30415, -60.13669, -59.9679, 
        -59.80006, -59.63528, -59.47465, -59.32145, -59.17543, -59.03671, 
        -58.90527, -58.77993, -58.65941, -58.54228, -58.42733, -58.3133, 
        -58.19972, -58.08587, -57.97226, -57.85857, -57.74444, -57.62968, 
        -57.51422, -57.398, -57.28045, -57.1618, -57.04263, -56.92363, 
        -56.80654, -56.69208, -56.5815, -56.47583, -56.3756, -56.28174, 
        -56.19419, -56.1132, -56.03882, -55.97092, -55.9095, -55.85387, 
        -55.80293, -55.75858, -55.71929, -55.68502, -55.65574, -55.63129, 
        -55.61137, -55.59595, -55.58513, -55.57858, -55.57638, -55.57805, 
        -55.58356, -55.59329, -55.60709, -55.62497, -55.64594, -55.66898, 
        -55.69386, -55.71979, -55.74526, -55.76901, -55.78985, -55.8066, 
        -55.81837, -55.82436, -55.82483, -55.82012, -55.81096, -55.79814, 
        -55.7821, -55.76372, -55.74352, -55.72213, -55.69949, -55.67506, 
        -55.64774, -55.61731, -55.58394, -55.54862, -55.51263, -55.4768, 
        -55.44261, -55.41199, -55.38673, -55.37219, -55.37082, -55.38573, 
        -55.41879,
  -44.37283, -44.56007, -44.74551, -44.93244, -45.12391, -45.32203, 
        -45.52833, -45.74345, -45.96834, -46.20377, -46.45044, -46.70944, 
        -46.97939, -47.2622, -47.55686, -47.86261, -48.17745, -48.49949, 
        -48.82544, -49.15238, -49.47685, -49.79762, -50.11473, -50.42958, 
        -50.74167, -51.05041, -51.3564, -51.65978, -51.96332, -52.26618, 
        -52.5677, -52.8655, -53.15666, -53.43761, -53.70527, -53.95667, 
        -54.18996, -54.40474, -54.60048, -54.77787, -54.93713, -55.07912, 
        -55.20452, -55.31646, -55.41516, -55.50259, -55.58091, -55.65276, 
        -55.7212, -55.78947, -55.86038, -55.93602, -56.01723, -56.10358, 
        -56.19302, -56.28284, -56.37106, -56.4556, -56.53489, -56.60762, 
        -56.67506, -56.7356, -56.7895, -56.83692, -56.87846, -56.91475, 
        -56.94611, -56.97417, -56.99994, -57.02555, -57.05322, -57.08489, 
        -57.12107, -57.16383, -57.21185, -57.26694, -57.32611, -57.39359, 
        -57.46833, -57.55223, -57.64872, -57.76025, -57.88906, -58.03668, 
        -58.20378, -58.39079, -58.59539, -58.81624, -59.05075, -59.29619, 
        -59.54963, -59.80765, -60.06733, -60.32418, -60.57319, -60.81176, 
        -61.03448, -61.23726, -61.41705, -61.57082, -61.69737, -61.79645, 
        -61.86961, -61.92001, -61.95097, -61.96689, -61.97144, -61.96859, 
        -61.96218, -61.95506, -61.94973, -61.94837, -61.95218, -61.96188, 
        -61.98038, -62.00763, -62.04373, -62.08848, -62.14149, -62.20184, 
        -62.26786, -62.33817, -62.41124, -62.48653, -62.56316, -62.64169, 
        -62.72157, -62.80249, -62.88411, -62.96591, -63.04813, -63.13074, 
        -63.21323, -63.29543, -63.3755, -63.4554, -63.53347, -63.60911, 
        -63.68151, -63.7498, -63.81314, -63.87075, -63.92145, -63.96431, 
        -63.99831, -64.02234, -64.03562, -64.03786, -64.0287, -64.00852, 
        -63.97807, -63.93828, -63.89043, -63.83609, -63.77711, -63.71528, 
        -63.65132, -63.58804, -63.52538, -63.46309, -63.4013, -63.33917, 
        -63.27629, -63.21219, -63.147, -63.08115, -63.01552, -62.95146, 
        -62.89012, -62.8326, -62.77989, -62.73288, -62.69172, -62.6562, 
        -62.62556, -62.59848, -62.57409, -62.55138, -62.52977, -62.50897, 
        -62.48851, -62.47022, -62.45277, -62.43513, -62.41589, -62.39428, 
        -62.36884, -62.33892, -62.30382, -62.26337, -62.2177, -62.16735, 
        -62.11272, -62.05432, -61.99218, -61.92679, -61.85858, -61.78685, 
        -61.71148, -61.63104, -61.54494, -61.45253, -61.35281, -61.24556, 
        -61.13065, -61.00852, -60.87952, -60.74373, -60.6011, -60.45337, 
        -60.29961, -60.14071, -59.97668, -59.80849, -59.63787, -59.46694, 
        -59.29781, -59.13269, -58.97367, -58.82209, -58.67866, -58.54273, 
        -58.41417, -58.29205, -58.17485, -58.06121, -57.94962, -57.83916, 
        -57.72903, -57.61893, -57.50875, -57.39851, -57.28812, -57.17672, 
        -57.0646, -56.95134, -56.837, -56.72163, -56.60589, -56.49006, 
        -56.37737, -56.26787, -56.16244, -56.062, -55.9668, -55.87749, 
        -55.79432, -55.71704, -55.64518, -55.57922, -55.51873, -55.46379, 
        -55.41446, -55.37059, -55.33221, -55.29894, -55.27071, -55.24733, 
        -55.22852, -55.21412, -55.20385, -55.19763, -55.19518, -55.19672, 
        -55.20223, -55.21201, -55.22613, -55.24463, -55.26705, -55.29224, 
        -55.31929, -55.34739, -55.37529, -55.40146, -55.42451, -55.44333, 
        -55.45689, -55.46487, -55.4675, -55.46423, -55.45761, -55.44732, 
        -55.43409, -55.41832, -55.40084, -55.38209, -55.3623, -55.34054, 
        -55.31576, -55.28732, -55.25562, -55.22176, -55.18696, -55.15194, 
        -55.11848, -55.08817, -55.06401, -55.04937, -55.04763, -55.0621, 
        -55.09476,
  -44.0312, -44.21527, -44.39844, -44.58372, -44.7747, -44.9739, 
        -45.18188, -45.39869, -45.62644, -45.86436, -46.11312, -46.37263, 
        -46.64303, -46.92434, -47.21619, -47.51826, -47.8292, -48.14704, 
        -48.4687, -48.79066, -49.10971, -49.42373, -49.73524, -50.0443, 
        -50.35073, -50.65502, -50.95773, -51.25904, -51.56025, -51.861, 
        -52.16034, -52.45567, -52.74374, -53.02103, -53.28474, -53.53144, 
        -53.75986, -53.96863, -54.15945, -54.33245, -54.48809, -54.62753, 
        -54.7527, -54.86457, -54.96427, -55.05307, -55.13328, -55.20724, 
        -55.27815, -55.34882, -55.42216, -55.50057, -55.58453, -55.67284, 
        -55.76518, -55.85804, -55.94915, -56.03647, -56.11876, -56.19529, 
        -56.26553, -56.32932, -56.3864, -56.43777, -56.48316, -56.523, 
        -56.55831, -56.58963, -56.61866, -56.64667, -56.67531, -56.70734, 
        -56.74471, -56.78738, -56.83501, -56.88815, -56.94666, -57.01232, 
        -57.0849, -57.16798, -57.26318, -57.37314, -57.50056, -57.64841, 
        -57.81748, -58.00658, -58.21497, -58.43936, -58.67748, -58.9267, 
        -59.18321, -59.44367, -59.70476, -59.96321, -60.21377, -60.45271, 
        -60.67574, -60.87877, -61.05886, -61.21314, -61.34016, -61.44001, 
        -61.51415, -61.5655, -61.59747, -61.6144, -61.61889, -61.61694, 
        -61.61073, -61.60323, -61.5963, -61.59211, -61.59265, -61.59949, 
        -61.61399, -61.63684, -61.66841, -61.70903, -61.75844, -61.81562, 
        -61.87904, -61.94693, -62.01801, -62.09115, -62.16576, -62.24203, 
        -62.31858, -62.39715, -62.47665, -62.55717, -62.63868, -62.72114, 
        -62.80425, -62.88752, -62.97035, -63.05238, -63.133, -63.2111, 
        -63.2859, -63.35622, -63.42103, -63.47931, -63.52996, -63.57175, 
        -63.60368, -63.6246, -63.63395, -63.63124, -63.61535, -63.58885, 
        -63.55152, -63.50447, -63.44912, -63.38715, -63.32051, -63.25111, 
        -63.18068, -63.11052, -63.04095, -62.97221, -62.90387, -62.83591, 
        -62.76749, -62.69808, -62.62827, -62.55845, -62.48954, -62.42293, 
        -62.3598, -62.30106, -62.24776, -62.19941, -62.15818, -62.12291, 
        -62.09264, -62.06668, -62.04366, -62.02294, -62.004, -61.98674, 
        -61.9711, -61.95742, -61.94438, -61.9314, -61.91629, -61.89785, 
        -61.87514, -61.8467, -61.81249, -61.77235, -61.72696, -61.67687, 
        -61.62259, -61.56479, -61.50326, -61.43852, -61.37084, -61.29946, 
        -61.22279, -61.1419, -61.05531, -60.96227, -60.86199, -60.75435, 
        -60.63902, -60.51665, -60.38739, -60.25147, -60.10877, -59.95977, 
        -59.80442, -59.64346, -59.47731, -59.30718, -59.13503, -58.96286, 
        -58.79328, -58.62846, -58.47044, -58.32045, -58.17925, -58.046, 
        -57.9201, -57.80073, -57.6867, -57.57642, -57.46827, -57.36157, 
        -57.25424, -57.14798, -57.04154, -56.93503, -56.8281, -56.7204, 
        -56.61171, -56.50195, -56.39131, -56.2802, -56.16902, -56.0591, 
        -55.9516, -55.84764, -55.74799, -55.653, -55.56293, -55.47811, 
        -55.39841, -55.32388, -55.25422, -55.18937, -55.12944, -55.07473, 
        -55.02549, -54.98196, -54.94427, -54.9118, -54.88429, -54.86171, 
        -54.84336, -54.82935, -54.81915, -54.81265, -54.80977, -54.81099, 
        -54.81527, -54.8252, -54.83989, -54.85938, -54.88327, -54.91068, 
        -54.94018, -54.97054, -55.00061, -55.02889, -55.05384, -55.07412, 
        -55.08913, -55.09887, -55.10345, -55.10333, -55.09919, -55.0916, 
        -55.08077, -55.06779, -55.05297, -55.03711, -55.02029, -55.00148, 
        -54.97963, -54.95415, -54.92553, -54.89453, -54.8621, -54.8295, 
        -54.79782, -54.76938, -54.74673, -54.73304, -54.73169, -54.74594, 
        -54.77803,
  -43.69745, -43.87862, -44.05894, -44.24323, -44.43402, -44.63391, 
        -44.84351, -45.06361, -45.29386, -45.53363, -45.78314, -46.04164, 
        -46.30989, -46.58727, -46.87373, -47.16938, -47.47301, -47.78396, 
        -48.09901, -48.41417, -48.72615, -49.03473, -49.33948, -49.64252, 
        -49.94321, -50.24267, -50.54065, -50.83847, -51.13636, -51.43437, 
        -51.73042, -52.02118, -52.30507, -52.57813, -52.83685, -53.07926, 
        -53.30339, -53.50893, -53.69636, -53.86629, -54.01983, -54.1586, 
        -54.28431, -54.39767, -54.49971, -54.59133, -54.67461, -54.75084, 
        -54.82489, -54.89848, -54.97469, -55.0556, -55.14207, -55.23362, 
        -55.32826, -55.42361, -55.51728, -55.60718, -55.69262, -55.77243, 
        -55.84638, -55.91403, -55.97612, -56.03235, -56.08203, -56.12777, 
        -56.16879, -56.20607, -56.24033, -56.27341, -56.30684, -56.34348, 
        -56.38377, -56.42891, -56.47856, -56.53274, -56.59214, -56.65766, 
        -56.73084, -56.81319, -56.90743, -57.01554, -57.14209, -57.28891, 
        -57.45681, -57.64662, -57.85516, -58.08108, -58.32056, -58.57064, 
        -58.828, -59.08821, -59.34904, -59.60613, -59.8553, -60.09249, 
        -60.31343, -60.51458, -60.69259, -60.84529, -60.97018, -61.06939, 
        -61.14358, -61.19584, -61.22921, -61.24796, -61.2558, -61.25591, 
        -61.25149, -61.24471, -61.23745, -61.2318, -61.22966, -61.23322, 
        -61.24364, -61.26182, -61.28849, -61.32409, -61.36883, -61.42085, 
        -61.4804, -61.545, -61.61288, -61.68334, -61.75557, -61.82894, 
        -61.90345, -61.9794, -62.05687, -62.13608, -62.21711, -62.30002, 
        -62.38416, -62.46908, -62.55415, -62.63857, -62.72161, -62.80206, 
        -62.87904, -62.95116, -63.01593, -63.07431, -63.12403, -63.16422, 
        -63.19336, -63.2107, -63.21546, -63.20734, -63.18646, -63.15328, 
        -63.10871, -63.0538, -62.99022, -62.91998, -62.8452, -62.76791, 
        -62.6897, -62.61193, -62.53518, -62.45944, -62.38505, -62.31108, 
        -62.23709, -62.16199, -62.08773, -62.01429, -61.94249, -61.87357, 
        -61.80869, -61.74905, -61.69503, -61.64721, -61.60558, -61.57016, 
        -61.54008, -61.51471, -61.49302, -61.47421, -61.45807, -61.44471, 
        -61.43398, -61.42515, -61.41726, -61.409, -61.39841, -61.38348, 
        -61.36304, -61.33628, -61.30217, -61.26271, -61.21745, -61.16755, 
        -61.11337, -61.05593, -60.99546, -60.9317, -60.8646, -60.7936, 
        -60.71803, -60.63713, -60.55014, -60.45683, -60.35634, -60.24873, 
        -60.13383, -60.01181, -59.88324, -59.74788, -59.60587, -59.4569, 
        -59.30161, -59.1403, -58.97381, -58.80342, -58.63131, -58.45949, 
        -58.28932, -58.12547, -57.96883, -57.82058, -57.681, -57.55, 
        -57.42653, -57.30952, -57.19813, -57.09076, -56.9859, -56.88269, 
        -56.78003, -56.67743, -56.57468, -56.47179, -56.36818, -56.26404, 
        -56.15905, -56.05313, -55.94658, -55.84005, -55.73415, -55.62984, 
        -55.5282, -55.43029, -55.33664, -55.2473, -55.16223, -55.08154, 
        -55.0048, -54.93231, -54.86397, -54.79984, -54.73926, -54.68462, 
        -54.63554, -54.59217, -54.55474, -54.52285, -54.49598, -54.47359, 
        -54.45533, -54.44083, -54.43007, -54.42301, -54.41953, -54.42013, 
        -54.42513, -54.43527, -54.45092, -54.47183, -54.4976, -54.52734, 
        -54.55946, -54.59219, -54.62419, -54.65426, -54.68084, -54.70233, 
        -54.71854, -54.72955, -54.73581, -54.73782, -54.73595, -54.7309, 
        -54.72281, -54.71237, -54.70049, -54.68779, -54.67404, -54.65838, 
        -54.64014, -54.61849, -54.59386, -54.56672, -54.53807, -54.50791, 
        -54.47966, -54.45406, -54.43394, -54.42204, -54.42181, -54.43629, 
        -54.46755,
  -43.37181, -43.55024, -43.72998, -43.91366, -44.10405, -44.30415, 
        -44.51493, -44.73625, -44.9676, -45.20803, -45.45644, -45.7113, 
        -45.97501, -46.24601, -46.52466, -46.81211, -47.10803, -47.41039, 
        -47.71677, -48.02408, -48.3287, -48.62965, -48.92758, -49.2241, 
        -49.51863, -49.81271, -50.10494, -50.39832, -50.69213, -50.98593, 
        -51.27773, -51.56473, -51.8436, -52.11104, -52.36501, -52.60303, 
        -52.82314, -53.02549, -53.21036, -53.37871, -53.53189, -53.67155, 
        -53.79809, -53.91421, -54.01952, -54.11508, -54.20246, -54.28384, 
        -54.36158, -54.43864, -54.51792, -54.60164, -54.69033, -54.78373, 
        -54.88025, -54.9776, -55.07346, -55.16635, -55.25397, -55.33749, 
        -55.41579, -55.4887, -55.55616, -55.61868, -55.67622, -55.72945, 
        -55.77832, -55.8233, -55.86515, -55.90514, -55.94546, -55.98816, 
        -56.0346, -56.08495, -56.13921, -56.19655, -56.25939, -56.32819, 
        -56.40385, -56.4879, -56.58305, -56.69135, -56.81673, -56.96133, 
        -57.12724, -57.31387, -57.52042, -57.74453, -57.98199, -58.23012, 
        -58.48503, -58.74311, -59.0008, -59.25382, -59.49938, -59.73244, 
        -59.94939, -60.14616, -60.31983, -60.46861, -60.59119, -60.68837, 
        -60.76169, -60.81382, -60.84842, -60.86946, -60.88031, -60.8836, 
        -60.88181, -60.8768, -60.87036, -60.86439, -60.85984, -60.86084, 
        -60.86742, -60.8809, -60.90254, -60.93299, -60.97227, -61.01996, 
        -61.07464, -61.1349, -61.19913, -61.26603, -61.33471, -61.40483, 
        -61.47647, -61.5499, -61.62571, -61.7039, -61.78516, -61.86915, 
        -61.95411, -62.04129, -62.12871, -62.21545, -62.3007, -62.38326, 
        -62.4617, -62.53458, -62.60048, -62.65826, -62.7065, -62.74393, 
        -62.76961, -62.78253, -62.78231, -62.76842, -62.74111, -62.70082, 
        -62.64847, -62.58551, -62.51361, -62.4349, -62.35169, -62.26517, 
        -62.17887, -62.0932, -62.00897, -61.92659, -61.84573, -61.76603, 
        -61.68701, -61.60842, -61.53046, -61.45401, -61.37982, -61.30918, 
        -61.2429, -61.1822, -61.12758, -61.07925, -61.03712, -61.00114, 
        -60.97082, -60.9457, -60.92493, -60.90804, -60.8952, -60.88486, 
        -60.87883, -60.87533, -60.87286, -60.86958, -60.86322, -60.85197, 
        -60.83427, -60.80938, -60.77732, -60.73825, -60.69329, -60.64352, 
        -60.5896, -60.53255, -60.47256, -60.40955, -60.34345, -60.27296, 
        -60.19776, -60.11684, -60.02989, -59.93659, -59.83656, -59.72958, 
        -59.61549, -59.49492, -59.36688, -59.23347, -59.09335, -58.94641, 
        -58.79282, -58.6331, -58.46822, -58.29956, -58.12901, -57.95889, 
        -57.79145, -57.62952, -57.47466, -57.32798, -57.18998, -57.06042, 
        -56.93889, -56.82378, -56.71447, -56.60936, -56.50733, -56.40705, 
        -56.30747, -56.20831, -56.10891, -56.0091, -55.90873, -55.80774, 
        -55.70627, -55.60405, -55.50171, -55.39894, -55.29839, -55.20023, 
        -55.10491, -55.01318, -54.92509, -54.8411, -54.76106, -54.68439, 
        -54.61053, -54.53971, -54.47236, -54.40892, -54.34968, -54.29527, 
        -54.24638, -54.20322, -54.16616, -54.13461, -54.10797, -54.08549, 
        -54.0667, -54.05134, -54.03952, -54.03122, -54.02675, -54.02658, 
        -54.03139, -54.04192, -54.0587, -54.08131, -54.10915, -54.14132, 
        -54.17607, -54.21139, -54.24553, -54.27708, -54.3047, -54.32741, 
        -54.34373, -54.35592, -54.36372, -54.36751, -54.36792, -54.36532, 
        -54.36005, -54.35271, -54.34415, -54.33471, -54.32439, -54.31247, 
        -54.298, -54.28082, -54.26059, -54.23796, -54.21384, -54.18918, 
        -54.16527, -54.14365, -54.12675, -54.11737, -54.11877, -54.1335, 
        -54.16409,
  -43.05563, -43.23196, -43.41012, -43.59299, -43.78286, -43.98259, 
        -44.1921, -44.41343, -44.6442, -44.88284, -45.12798, -45.37913, 
        -45.63605, -45.89885, -46.16831, -46.44579, -46.73143, -47.02414, 
        -47.32088, -47.61982, -47.91683, -48.20945, -48.50035, -48.78949, 
        -49.07854, -49.36666, -49.6547, -49.9429, -50.23167, -50.51996, 
        -50.80584, -51.08683, -51.3595, -51.62134, -51.86984, -52.1032, 
        -52.31885, -52.51869, -52.70211, -52.87009, -53.02421, -53.16565, 
        -53.29573, -53.41523, -53.52458, -53.6246, -53.71673, -53.8027, 
        -53.88498, -53.96595, -54.04894, -54.13541, -54.22515, -54.32032, 
        -54.41843, -54.51762, -54.61575, -54.71129, -54.80328, -54.89109, 
        -54.97454, -55.05314, -55.1268, -55.19644, -55.26215, -55.32423, 
        -55.38246, -55.4366, -55.48732, -55.53536, -55.58433, -55.63591, 
        -55.69065, -55.7489, -55.81034, -55.87556, -55.94529, -56.02002, 
        -56.10061, -56.18966, -56.2874, -56.39668, -56.52211, -56.66449, 
        -56.82692, -57.00923, -57.21021, -57.4283, -57.66096, -57.90432, 
        -58.15501, -58.40866, -58.66161, -58.91037, -59.15031, -59.37741, 
        -59.58804, -59.77838, -59.94541, -60.08787, -60.2054, -60.29827, 
        -60.36896, -60.41988, -60.45518, -60.47735, -60.49118, -60.49779, 
        -60.499, -60.49673, -60.49226, -60.48695, -60.48327, -60.48227, 
        -60.48563, -60.49516, -60.51202, -60.53714, -60.57056, -60.6124, 
        -60.66174, -60.71684, -60.77659, -60.83924, -60.90405, -60.96983, 
        -61.03858, -61.10975, -61.18393, -61.26195, -61.34409, -61.4298, 
        -61.518, -61.60766, -61.6979, -61.78712, -61.87435, -61.95823, 
        -62.03711, -62.10994, -62.17506, -62.23103, -62.27657, -62.31033, 
        -62.33149, -62.33921, -62.33305, -62.31187, -62.27775, -62.23023, 
        -62.1702, -62.09909, -62.01888, -61.93192, -61.84036, -61.74641, 
        -61.65196, -61.55844, -61.46695, -61.3777, -61.29079, -61.20572, 
        -61.12204, -61.03981, -60.95885, -60.87996, -60.8041, -60.73215, 
        -60.66522, -60.60398, -60.54787, -60.49895, -60.45618, -60.41976, 
        -60.38907, -60.36385, -60.34367, -60.32855, -60.31859, -60.31323, 
        -60.31212, -60.31384, -60.31673, -60.31812, -60.31592, -60.30806, 
        -60.29315, -60.27018, -60.23899, -60.20058, -60.15594, -60.10622, 
        -60.05239, -59.99529, -59.93579, -59.87363, -59.80705, -59.73731, 
        -59.66232, -59.58187, -59.49549, -59.40281, -59.30353, -59.1978, 
        -59.0857, -58.96734, -58.84293, -58.71239, -58.57572, -58.43219, 
        -58.28204, -58.12591, -57.96454, -57.79953, -57.63259, -57.46558, 
        -57.30118, -57.1417, -56.98912, -56.84428, -56.70764, -56.57917, 
        -56.45844, -56.34478, -56.23687, -56.13344, -56.03236, -55.93438, 
        -55.83752, -55.74088, -55.64421, -55.54708, -55.44914, -55.35114, 
        -55.25275, -55.15387, -55.05536, -54.95806, -54.86297, -54.77056, 
        -54.68133, -54.59554, -54.51327, -54.43469, -54.35927, -54.2863, 
        -54.21529, -54.14627, -54.08023, -54.01748, -53.95883, -53.90517, 
        -53.85688, -53.81437, -53.77754, -53.74613, -53.71943, -53.69654, 
        -53.67696, -53.66032, -53.64687, -53.63599, -53.63021, -53.62929, 
        -53.63379, -53.64481, -53.66281, -53.68731, -53.71748, -53.75208, 
        -53.78944, -53.82722, -53.86335, -53.8962, -53.92474, -53.94835, 
        -53.96679, -53.98022, -53.9894, -53.99511, -53.99785, -53.99802, 
        -53.9959, -53.99212, -53.9871, -53.98142, -53.97475, -53.96675, 
        -53.95655, -53.94382, -53.92831, -53.91056, -53.89119, -53.87136, 
        -53.8522, -53.83522, -53.82232, -53.8161, -53.81946, -53.83485, 
        -53.86436,
  -42.74518, -42.91895, -43.09566, -43.27763, -43.46671, -43.66518, 
        -43.87445, -44.09378, -44.32214, -44.55684, -44.79692, -45.04112, 
        -45.2896, -45.54305, -45.80238, -46.06788, -46.34228, -46.62386, 
        -46.91046, -47.19966, -47.4881, -47.77456, -48.05883, -48.34238, 
        -48.6263, -48.90908, -49.19144, -49.47425, -49.75699, -50.03888, 
        -50.31801, -50.59076, -50.85647, -51.11151, -51.35415, -51.58266, 
        -51.79564, -51.99333, -52.17585, -52.34401, -52.49916, -52.6428, 
        -52.77603, -52.89907, -53.01247, -53.11711, -53.21305, -53.30396, 
        -53.39106, -53.47669, -53.56337, -53.65257, -53.74579, -53.84317, 
        -53.94314, -54.04436, -54.145, -54.24363, -54.33928, -54.43181, 
        -54.52047, -54.605, -54.68561, -54.76202, -54.83626, -54.90754, 
        -54.97542, -55.03923, -55.10025, -55.15939, -55.21905, -55.2811, 
        -55.34594, -55.41381, -55.48524, -55.55999, -55.63884, -55.722, 
        -55.81096, -55.90696, -56.00978, -56.12265, -56.24863, -56.39068, 
        -56.55072, -56.72804, -56.9239, -57.1364, -57.36232, -57.59848, 
        -57.84173, -58.089, -58.33559, -58.57713, -58.80986, -59.02931, 
        -59.23164, -59.41324, -59.57059, -59.70485, -59.81472, -59.90131, 
        -59.96727, -60.01566, -60.05029, -60.07438, -60.09032, -60.09981, 
        -60.10445, -60.10517, -60.10328, -60.09978, -60.09634, -60.09446, 
        -60.09575, -60.10202, -60.11475, -60.13487, -60.16196, -60.19795, 
        -60.24159, -60.29136, -60.34602, -60.40379, -60.46421, -60.5273, 
        -60.59327, -60.66255, -60.73589, -60.81416, -60.89774, -60.98554, 
        -61.07636, -61.16882, -61.26192, -61.35334, -61.44209, -61.52644, 
        -61.60498, -61.67543, -61.73826, -61.79113, -61.83272, -61.86184, 
        -61.87762, -61.8795, -61.86718, -61.84026, -61.79909, -61.74437, 
        -61.67694, -61.59782, -61.50969, -61.41445, -61.31468, -61.21272, 
        -61.11035, -61.00939, -60.91074, -60.81514, -60.72239, -60.6314, 
        -60.54391, -60.4588, -60.37582, -60.29551, -60.21862, -60.14613, 
        -60.07909, -60.01764, -59.96217, -59.91265, -59.86941, -59.83241, 
        -59.80109, -59.77556, -59.75613, -59.74277, -59.73542, -59.7336, 
        -59.73653, -59.74308, -59.75071, -59.75673, -59.75835, -59.75381, 
        -59.74039, -59.71897, -59.68874, -59.65078, -59.60627, -59.55641, 
        -59.50254, -59.44567, -59.38642, -59.32469, -59.25936, -59.18993, 
        -59.11566, -59.03609, -58.95068, -58.85917, -58.76146, -58.65798, 
        -58.54862, -58.43364, -58.313, -58.18657, -58.05421, -57.91533, 
        -57.77014, -57.6189, -57.46252, -57.30234, -57.1402, -56.97709, 
        -56.81648, -56.66061, -56.51112, -56.36845, -56.23323, -56.10576, 
        -55.98579, -55.87292, -55.76594, -55.66369, -55.56476, -55.46833, 
        -55.37324, -55.27866, -55.18377, -55.08859, -54.99308, -54.89729, 
        -54.80124, -54.7051, -54.60948, -54.51612, -54.42538, -54.33783, 
        -54.25371, -54.17332, -54.09646, -54.0229, -53.95197, -53.88268, 
        -53.81502, -53.74884, -53.68356, -53.62231, -53.56498, -53.5126, 
        -53.46576, -53.4243, -53.38815, -53.35696, -53.32986, -53.30637, 
        -53.28563, -53.26738, -53.25201, -53.24018, -53.23282, -53.23085, 
        -53.23518, -53.24652, -53.2656, -53.2919, -53.32465, -53.36166, 
        -53.40126, -53.44121, -53.47924, -53.51339, -53.54285, -53.56716, 
        -53.58663, -53.60123, -53.61179, -53.61963, -53.62511, -53.62855, 
        -53.6302, -53.63032, -53.62948, -53.62778, -53.6252, -53.62137, 
        -53.6154, -53.60696, -53.59516, -53.5822, -53.56792, -53.55313, 
        -53.53885, -53.52666, -53.51809, -53.51515, -53.52043, -53.53633, 
        -53.56485,
  -42.43694, -42.61165, -42.78713, -42.96712, -43.15492, -43.35185, 
        -43.55844, -43.77444, -43.99823, -44.22731, -44.4596, -44.69584, 
        -44.93478, -45.1779, -45.42641, -45.68164, -45.94414, -46.21413, 
        -46.48983, -46.76926, -47.04957, -47.32882, -47.60729, -47.8854, 
        -48.1635, -48.44027, -48.71735, -48.99406, -49.27042, -49.54508, 
        -49.81623, -50.08215, -50.34003, -50.5879, -50.82413, -51.04756, 
        -51.25728, -51.4524, -51.63392, -51.80222, -51.95872, -52.10313, 
        -52.23873, -52.3648, -52.48209, -52.59095, -52.69251, -52.78852, 
        -52.88058, -52.97097, -53.06142, -53.15428, -53.2504, -53.35014, 
        -53.45245, -53.55608, -53.65947, -53.76038, -53.86003, -53.95718, 
        -54.05107, -54.14199, -54.22978, -54.31509, -54.3982, -54.47855, 
        -54.55572, -54.62968, -54.70115, -54.77135, -54.84261, -54.91554, 
        -54.99172, -55.07119, -55.15277, -55.23911, -55.32938, -55.42408, 
        -55.5235, -55.62862, -55.73982, -55.8595, -55.98999, -56.13363, 
        -56.29163, -56.4651, -56.65588, -56.86148, -57.0799, -57.30841, 
        -57.54404, -57.78294, -58.02037, -58.25399, -58.47827, -58.68839, 
        -58.88085, -59.05223, -59.20008, -59.32396, -59.42414, -59.50242, 
        -59.56182, -59.60577, -59.63804, -59.66116, -59.67809, -59.6897, 
        -59.69693, -59.70068, -59.70145, -59.6992, -59.69705, -59.69511, 
        -59.69522, -59.6992, -59.70853, -59.72437, -59.74752, -59.77835, 
        -59.81642, -59.86071, -59.90981, -59.96261, -60.0188, -60.07834, 
        -60.1417, -60.20949, -60.28232, -60.3612, -60.44605, -60.53505, 
        -60.62867, -60.7241, -60.81975, -60.91306, -61.00258, -61.08662, 
        -61.16366, -61.23246, -61.2917, -61.34011, -61.37664, -61.40012, 
        -61.40986, -61.40533, -61.38627, -61.35264, -61.30461, -61.24265, 
        -61.16775, -61.08131, -60.98578, -60.88212, -60.77512, -60.66563, 
        -60.556, -60.44786, -60.34278, -60.2412, -60.14334, -60.04906, 
        -59.95827, -59.871, -59.78681, -59.706, -59.62913, -59.5569, 
        -59.49018, -59.42907, -59.37363, -59.32402, -59.28035, -59.24287, 
        -59.21129, -59.18579, -59.16671, -59.15364, -59.14812, -59.14922, 
        -59.1558, -59.16606, -59.17773, -59.18756, -59.19277, -59.19071, 
        -59.18019, -59.16011, -59.13069, -59.09303, -59.04829, -58.9982, 
        -58.94421, -58.88734, -58.82816, -58.76654, -58.70171, -58.63287, 
        -58.55944, -58.48104, -58.3973, -58.30756, -58.21245, -58.11211, 
        -58.00568, -57.89494, -57.77887, -57.65741, -57.53039, -57.39719, 
        -57.25779, -57.11241, -56.96219, -56.80814, -56.6517, -56.49503, 
        -56.33994, -56.18813, -56.04191, -55.90187, -55.76838, -55.64184, 
        -55.52256, -55.41031, -55.30399, -55.20225, -55.10413, -55.00869, 
        -54.91466, -54.82124, -54.72791, -54.63401, -54.53997, -54.44571, 
        -54.35107, -54.25587, -54.1628, -54.07209, -53.98494, -53.90109, 
        -53.82112, -53.74494, -53.67285, -53.60386, -53.53699, -53.47168, 
        -53.40741, -53.34442, -53.28319, -53.2244, -53.16928, -53.11864, 
        -53.07376, -53.03408, -52.99899, -52.96809, -52.94072, -52.91628, 
        -52.89425, -52.87437, -52.85697, -52.84319, -52.83412, -52.83106, 
        -52.83496, -52.84678, -52.86697, -52.89503, -52.9297, -52.9691, 
        -53.01073, -53.05239, -53.09201, -53.1274, -53.15665, -53.18166, 
        -53.20169, -53.2175, -53.22992, -53.24002, -53.24857, -53.256, 
        -53.26195, -53.2668, -53.27043, -53.27322, -53.27509, -53.27524, 
        -53.27337, -53.26912, -53.26268, -53.25437, -53.24489, -53.23502, 
        -53.22593, -53.21851, -53.21416, -53.21477, -53.22231, -53.23875, 
        -53.26598,
  -42.13205, -42.30612, -42.48067, -42.65928, -42.84487, -43.03805, 
        -43.2411, -43.45256, -43.67043, -43.89242, -44.1178, -44.34539, 
        -44.57459, -44.80717, -45.04496, -45.28858, -45.53933, -45.79785, 
        -46.06225, -46.33142, -46.60233, -46.87529, -47.148, -47.42098, 
        -47.69381, -47.96613, -48.23751, -48.50817, -48.77727, -49.04404, 
        -49.30694, -49.56476, -49.8146, -50.05433, -50.28458, -50.50128, 
        -50.70694, -50.90023, -51.08013, -51.24765, -51.40458, -51.55116, 
        -51.68856, -51.81692, -51.93701, -52.04927, -52.15496, -52.25549, 
        -52.35249, -52.44746, -52.54237, -52.63811, -52.73767, -52.84039, 
        -52.94532, -53.0518, -53.15805, -53.26336, -53.3671, -53.46892, 
        -53.56848, -53.66567, -53.76085, -53.85396, -53.94537, -54.03439, 
        -54.12067, -54.20454, -54.28528, -54.36634, -54.44895, -54.53346, 
        -54.62165, -54.71294, -54.8079, -54.90713, -55.01068, -55.11815, 
        -55.22988, -55.34605, -55.46779, -55.59646, -55.73347, -55.88034, 
        -56.03863, -56.20961, -56.3967, -56.59724, -56.80827, -57.02945, 
        -57.25712, -57.48771, -57.71771, -57.94242, -58.15722, -58.35726, 
        -58.53885, -58.69865, -58.83461, -58.94658, -59.03558, -59.10391, 
        -59.15483, -59.1924, -59.2191, -59.23958, -59.25584, -59.26818, 
        -59.27702, -59.28306, -59.28632, -59.28737, -59.28654, -59.28542, 
        -59.28525, -59.28771, -59.29458, -59.30694, -59.32601, -59.3522, 
        -59.38535, -59.42412, -59.46788, -59.51585, -59.56666, -59.62276, 
        -59.68369, -59.75014, -59.82288, -59.90272, -59.98915, -60.08133, 
        -60.17738, -60.27512, -60.37261, -60.46714, -60.55678, -60.63936, 
        -60.71382, -60.77876, -60.83322, -60.87615, -60.9065, -60.92358, 
        -60.92665, -60.9143, -60.88839, -60.84806, -60.79334, -60.7247, 
        -60.64324, -60.55036, -60.44846, -60.33945, -60.22582, -60.10987, 
        -59.99382, -59.87966, -59.76875, -59.66179, -59.55931, -59.46125, 
        -59.36792, -59.27919, -59.19465, -59.11418, -59.03792, -58.96682, 
        -58.901, -58.83966, -58.78486, -58.73557, -58.69216, -58.65472, 
        -58.62283, -58.59745, -58.57877, -58.56766, -58.56388, -58.56685, 
        -58.57583, -58.58883, -58.60323, -58.61581, -58.62363, -58.62376, 
        -58.61477, -58.59516, -58.56621, -58.52827, -58.4832, -58.43262, 
        -58.37829, -58.32127, -58.26109, -58.19953, -58.13502, -58.06703, 
        -57.99506, -57.91838, -57.83712, -57.7504, -57.65892, -57.56242, 
        -57.46143, -57.35595, -57.24531, -57.1296, -57.00832, -56.88121, 
        -56.74817, -56.60936, -56.46556, -56.31823, -56.16836, -56.01779, 
        -55.868, -55.72139, -55.57907, -55.44184, -55.31058, -55.1855, 
        -55.06722, -54.95551, -54.84848, -54.74699, -54.64922, -54.55442, 
        -54.46125, -54.36865, -54.2762, -54.18319, -54.08989, -53.99636, 
        -53.90242, -53.80931, -53.71768, -53.62896, -53.54404, -53.4628, 
        -53.3858, -53.3129, -53.24427, -53.17932, -53.11638, -53.0546, 
        -52.994, -52.93468, -52.87704, -52.8218, -52.76994, -52.72213, 
        -52.67926, -52.64148, -52.60769, -52.57706, -52.54945, -52.5241, 
        -52.5006, -52.47829, -52.45923, -52.44365, -52.43317, -52.42918, 
        -52.43272, -52.44498, -52.46617, -52.4957, -52.53204, -52.57314, 
        -52.61663, -52.65974, -52.70048, -52.73691, -52.76786, -52.79337, 
        -52.81404, -52.83094, -52.84532, -52.85805, -52.8702, -52.88205, 
        -52.89304, -52.90315, -52.91194, -52.91964, -52.92588, -52.93003, 
        -52.932, -52.93159, -52.92926, -52.92528, -52.92048, -52.91569, 
        -52.91154, -52.9089, -52.90874, -52.91276, -52.92253, -52.93966, 
        -52.96607,
  -41.82761, -42.00277, -42.17503, -42.34802, -42.53237, -42.72325, 
        -42.92308, -43.12927, -43.34064, -43.55451, -43.77147, -43.99015, 
        -44.20996, -44.43279, -44.6601, -44.89194, -45.13131, -45.37816, 
        -45.63107, -45.89093, -46.15435, -46.42038, -46.68707, -46.95495, 
        -47.22233, -47.48898, -47.75413, -48.0176, -48.2794, -48.53805, 
        -48.79137, -49.04045, -49.28161, -49.51431, -49.73765, -49.95039, 
        -50.15168, -50.34173, -50.51933, -50.68587, -50.84232, -50.98917, 
        -51.12747, -51.2575, -51.37954, -51.49343, -51.60231, -51.70676, 
        -51.80799, -51.90755, -52.00707, -52.10815, -52.21175, -52.31752, 
        -52.42575, -52.53508, -52.64429, -52.75323, -52.8609, -52.96725, 
        -53.07205, -53.17564, -53.27682, -53.37757, -53.4768, -53.57396, 
        -53.66895, -53.76191, -53.85362, -53.94557, -54.03872, -54.13475, 
        -54.23445, -54.3382, -54.44604, -54.55847, -54.67564, -54.79625, 
        -54.9209, -55.04837, -55.18148, -55.32003, -55.46511, -55.6179, 
        -55.78049, -55.95402, -56.13938, -56.33627, -56.54338, -56.75819, 
        -56.97906, -57.2025, -57.42439, -57.64019, -57.84517, -58.03461, 
        -58.20448, -58.35067, -58.47358, -58.57262, -58.64923, -58.7066, 
        -58.74789, -58.77727, -58.79849, -58.81477, -58.82858, -58.83984, 
        -58.849, -58.85612, -58.86139, -58.86415, -58.86472, -58.86443, 
        -58.86443, -58.86615, -58.87115, -58.88004, -58.89589, -58.91809, 
        -58.94664, -58.98045, -59.01916, -59.06249, -59.11062, -59.16339, 
        -59.22216, -59.2876, -59.36044, -59.44107, -59.5289, -59.62279, 
        -59.72058, -59.82, -59.91863, -60.01329, -60.10168, -60.18184, 
        -60.2516, -60.31181, -60.36055, -60.3972, -60.42084, -60.43121, 
        -60.42738, -60.40926, -60.37674, -60.32997, -60.2692, -60.19486, 
        -60.1079, -60.00972, -59.90233, -59.78804, -59.66903, -59.54771, 
        -59.42631, -59.30701, -59.19118, -59.07978, -58.97242, -58.87136, 
        -58.77613, -58.68655, -58.60212, -58.52246, -58.44761, -58.37789, 
        -58.31371, -58.25479, -58.20108, -58.1526, -58.10985, -58.07281, 
        -58.04129, -58.01625, -57.99805, -57.98751, -57.98474, -57.98895, 
        -57.99908, -58.01313, -58.02888, -58.04292, -58.05196, -58.05222, 
        -58.04388, -58.02477, -57.9956, -57.95713, -57.91146, -57.86036, 
        -57.80556, -57.74826, -57.68901, -57.62762, -57.56379, -57.4969, 
        -57.42667, -57.35267, -57.27468, -57.19214, -57.10527, -57.01416, 
        -56.9185, -56.81841, -56.71379, -56.60408, -56.48899, -56.36806, 
        -56.24119, -56.10876, -55.97172, -55.83007, -55.68669, -55.54224, 
        -55.39839, -55.25709, -55.11914, -54.98571, -54.85725, -54.73444, 
        -54.61766, -54.50694, -54.40119, -54.29992, -54.20228, -54.10792, 
        -54.01535, -53.92334, -53.83126, -53.73877, -53.64584, -53.55265, 
        -53.45925, -53.36657, -53.27572, -53.18776, -53.10357, -53.02384, 
        -52.94859, -52.87776, -52.81131, -52.74914, -52.68959, -52.63124, 
        -52.5732, -52.51782, -52.46444, -52.41331, -52.36539, -52.32084, 
        -52.28049, -52.24431, -52.21174, -52.18173, -52.15368, -52.12722, 
        -52.10255, -52.0796, -52.05924, -52.04248, -52.03114, -52.02649, 
        -52.03016, -52.04298, -52.06506, -52.0958, -52.13376, -52.17641, 
        -52.22121, -52.26548, -52.30692, -52.34397, -52.37545, -52.40118, 
        -52.42228, -52.44027, -52.45656, -52.47229, -52.48825, -52.5047, 
        -52.52124, -52.53691, -52.55159, -52.56475, -52.57549, -52.58284, 
        -52.58852, -52.5918, -52.59323, -52.59344, -52.59339, -52.59343, 
        -52.5941, -52.59626, -52.60041, -52.60783, -52.61965, -52.63772, 
        -52.66324,
  -41.52785, -41.70296, -41.87238, -42.04084, -42.21759, -42.39802, 
        -42.60176, -42.80507, -43.00959, -43.21506, -43.42364, -43.63274, 
        -43.84351, -44.05763, -44.27586, -44.4992, -44.72783, -44.96307, 
        -45.20512, -45.45517, -45.70866, -45.9683, -46.22859, -46.49032, 
        -46.75047, -47.01057, -47.26891, -47.52512, -47.77905, -48.02969, 
        -48.27573, -48.5156, -48.74848, -48.97406, -49.19048, -49.39766, 
        -49.59441, -49.78046, -49.95593, -50.12024, -50.27459, -50.42102, 
        -50.55941, -50.68995, -50.8132, -50.9297, -51.04113, -51.14874, 
        -51.25372, -51.35767, -51.4618, -51.56734, -51.67501, -51.78443, 
        -51.89569, -52.00799, -52.11914, -52.23106, -52.34239, -52.45335, 
        -52.56352, -52.67313, -52.78196, -52.88977, -52.99622, -53.10096, 
        -53.20411, -53.30576, -53.4067, -53.5085, -53.6122, -53.71917, 
        -53.83017, -53.94482, -54.06509, -54.19051, -54.32045, -54.45419, 
        -54.59145, -54.73258, -54.87742, -55.02683, -55.18173, -55.34274, 
        -55.51141, -55.68894, -55.87582, -56.07206, -56.2768, -56.48816, 
        -56.70471, -56.92085, -57.13587, -57.34334, -57.53875, -57.7173, 
        -57.87505, -58.00935, -58.1188, -58.20432, -58.26807, -58.31365, 
        -58.34444, -58.36451, -58.37814, -58.38847, -58.39798, -58.40673, 
        -58.41463, -58.42175, -58.4264, -58.43017, -58.43189, -58.43215, 
        -58.43245, -58.43365, -58.43756, -58.4456, -58.45877, -58.47768, 
        -58.50202, -58.53169, -58.56602, -58.60511, -58.6497, -58.69983, 
        -58.75647, -58.82111, -58.89383, -58.97521, -59.06297, -59.15795, 
        -59.25677, -59.35674, -59.45512, -59.54871, -59.63478, -59.71157, 
        -59.77769, -59.83242, -59.87503, -59.905, -59.92181, -59.92525, 
        -59.91457, -59.88994, -59.85136, -59.79891, -59.73305, -59.65407, 
        -59.56285, -59.46072, -59.34848, -59.23029, -59.10725, -58.98176, 
        -58.85614, -58.7327, -58.61298, -58.49809, -58.38866, -58.28513, 
        -58.1884, -58.09843, -58.01445, -57.93603, -57.86286, -57.7951, 
        -57.73275, -57.67566, -57.62367, -57.57661, -57.53504, -57.49881, 
        -57.46809, -57.44363, -57.425, -57.4148, -57.41228, -57.41666, 
        -57.42659, -57.44044, -57.45586, -57.46968, -57.47871, -57.48021, 
        -57.47132, -57.45166, -57.42189, -57.38299, -57.33661, -57.28487, 
        -57.22965, -57.17193, -57.1127, -57.0518, -56.98918, -56.92397, 
        -56.85647, -56.78597, -56.71228, -56.6349, -56.55344, -56.46705, 
        -56.37744, -56.28337, -56.18457, -56.081, -55.97198, -55.85711, 
        -55.73645, -55.61018, -55.47932, -55.34495, -55.20797, -55.06958, 
        -54.93161, -54.7957, -54.66285, -54.53358, -54.40894, -54.28917, 
        -54.17456, -54.06535, -53.96052, -53.85971, -53.76225, -53.66807, 
        -53.57594, -53.48441, -53.3926, -53.30023, -53.20731, -53.11332, 
        -53.02027, -52.92787, -52.83723, -52.7497, -52.6658, -52.5863, 
        -52.5114, -52.44119, -52.37595, -52.31533, -52.25787, -52.2026, 
        -52.14899, -52.09742, -52.04832, -52.00154, -51.95745, -51.91654, 
        -51.87844, -51.84367, -51.81172, -51.78199, -51.75335, -51.7258, 
        -51.69962, -51.6755, -51.6541, -51.63713, -51.6256, -51.62132, 
        -51.62546, -51.63908, -51.6623, -51.6941, -51.7331, -51.77705, 
        -51.82285, -51.86716, -51.90918, -51.94653, -51.97828, -52.00433, 
        -52.0257, -52.04477, -52.06274, -52.08147, -52.10131, -52.12251, 
        -52.14455, -52.16643, -52.18731, -52.20603, -52.22178, -52.23434, 
        -52.24377, -52.25061, -52.25583, -52.26042, -52.26496, -52.2699, 
        -52.27544, -52.28229, -52.2906, -52.30142, -52.31579, -52.33489, 
        -52.36006,
  -41.22919, -41.40266, -41.57093, -41.73972, -41.91363, -42.09597, 
        -42.2855, -42.4807, -42.67805, -42.8772, -43.07766, -43.27906, 
        -43.48244, -43.68988, -43.90018, -44.11493, -44.33457, -44.55927, 
        -44.79147, -45.02891, -45.27441, -45.52366, -45.77688, -46.03059, 
        -46.28443, -46.53674, -46.78725, -47.0357, -47.28126, -47.52335, 
        -47.76077, -47.99264, -48.21741, -48.43524, -48.6442, -48.84606, 
        -49.03789, -49.2199, -49.39173, -49.55376, -49.70752, -49.85332, 
        -49.99149, -50.12222, -50.24588, -50.36348, -50.4765, -50.58639, 
        -50.69481, -50.80281, -50.91004, -51.01984, -51.13116, -51.24416, 
        -51.35872, -51.47371, -51.58858, -51.70333, -51.81838, -51.93316, 
        -52.04817, -52.16354, -52.27841, -52.39269, -52.50581, -52.61792, 
        -52.72853, -52.83708, -52.94683, -53.05788, -53.17161, -53.28902, 
        -53.41071, -53.53753, -53.66939, -53.80676, -53.94857, -54.09398, 
        -54.24292, -54.39566, -54.55196, -54.71296, -54.8779, -55.04812, 
        -55.22371, -55.40704, -55.59793, -55.79643, -56.00178, -56.21276, 
        -56.42684, -56.64055, -56.84964, -57.0499, -57.23618, -57.40395, 
        -57.54975, -57.67113, -57.76722, -57.83939, -57.89019, -57.92363, 
        -57.94307, -57.95235, -57.95766, -57.96129, -57.96519, -57.96999, 
        -57.97525, -57.98087, -57.98567, -57.98935, -57.99117, -57.99174, 
        -57.99191, -57.99261, -57.9957, -58.00228, -58.01333, -58.02935, 
        -58.05026, -58.07588, -58.10637, -58.14065, -58.18181, -58.22954, 
        -58.28491, -58.34862, -58.42127, -58.50306, -58.59223, -58.68769, 
        -58.78643, -58.88573, -58.98251, -59.07374, -59.15654, -59.22915, 
        -59.29021, -59.33915, -59.37548, -59.3988, -59.40891, -59.40567, 
        -59.38765, -59.35709, -59.31306, -59.25586, -59.18593, -59.10345, 
        -59.00939, -58.90472, -58.79114, -58.67073, -58.54538, -58.41706, 
        -58.28844, -58.16176, -58.0393, -57.92189, -57.81028, -57.70518, 
        -57.60748, -57.51728, -57.43391, -57.35682, -57.28537, -57.21872, 
        -57.15871, -57.10361, -57.0535, -57.0083, -56.9682, -56.93335, 
        -56.90368, -56.8803, -56.86296, -56.85291, -56.85012, -56.85346, 
        -56.86185, -56.87365, -56.88684, -56.89893, -56.90643, -56.9064, 
        -56.89646, -56.87597, -56.84531, -56.80563, -56.75873, -56.70668, 
        -56.65109, -56.59261, -56.53358, -56.47392, -56.41238, -56.34953, 
        -56.28564, -56.21931, -56.15049, -56.07869, -56.0034, -55.9244, 
        -55.84092, -55.75313, -55.66032, -55.56258, -55.45956, -55.35036, 
        -55.23532, -55.11474, -54.98978, -54.86143, -54.73049, -54.59843, 
        -54.46621, -54.33587, -54.20856, -54.08439, -53.96386, -53.84789, 
        -53.7355, -53.62815, -53.52471, -53.42476, -53.32792, -53.23391, 
        -53.1418, -53.0506, -52.95892, -52.86658, -52.77403, -52.68118, 
        -52.58845, -52.49657, -52.40634, -52.31882, -52.23487, -52.15477, 
        -52.07949, -52.00892, -51.94357, -51.88315, -51.82709, -51.77389, 
        -51.72349, -51.67496, -51.62953, -51.58649, -51.54603, -51.50796, 
        -51.47203, -51.43803, -51.40594, -51.37535, -51.34583, -51.31606, 
        -51.28843, -51.26321, -51.24152, -51.2247, -51.21406, -51.21094, 
        -51.21642, -51.23142, -51.25596, -51.28914, -51.32914, -51.37391, 
        -51.4207, -51.46642, -51.50883, -51.54636, -51.57808, -51.6045, 
        -51.62614, -51.64595, -51.66605, -51.68758, -51.71115, -51.73699, 
        -51.76458, -51.7927, -51.81966, -51.84433, -51.86556, -51.88276, 
        -51.89634, -51.90712, -51.91616, -51.925, -51.93417, -51.94395, 
        -51.95433, -51.96557, -51.97822, -51.9927, -52.0099, -52.03065, 
        -52.05635,
  -40.93605, -41.1096, -41.2782, -41.44447, -41.61689, -41.78893, 
        -41.97347, -42.16219, -42.34856, -42.54162, -42.73748, -42.93359, 
        -43.13281, -43.3332, -43.53507, -43.74352, -43.95515, -44.17138, 
        -44.39274, -44.62134, -44.85604, -45.09652, -45.33969, -45.58389, 
        -45.82846, -46.07135, -46.31303, -46.55237, -46.78904, -47.0216, 
        -47.25036, -47.47355, -47.69048, -47.90115, -48.10484, -48.30076, 
        -48.48771, -48.66548, -48.8338, -48.99349, -49.14534, -49.29023, 
        -49.42802, -49.55866, -49.68278, -49.8002, -49.91418, -50.02584, 
        -50.13687, -50.2481, -50.36009, -50.47347, -50.58821, -50.70446, 
        -50.82173, -50.93924, -51.05632, -51.1738, -51.29173, -51.41043, 
        -51.52985, -51.64914, -51.76977, -51.89009, -52.00968, -52.12841, 
        -52.24575, -52.36283, -52.48059, -52.60039, -52.72344, -52.85043, 
        -52.98252, -53.11968, -53.26171, -53.40928, -53.56131, -53.71731, 
        -53.87595, -54.03908, -54.20606, -54.37692, -54.55252, -54.73232, 
        -54.91727, -55.10828, -55.30515, -55.5084, -55.71719, -55.93009, 
        -56.14427, -56.35604, -56.56131, -56.7551, -56.93324, -57.09077, 
        -57.22406, -57.33269, -57.41564, -57.47472, -57.51306, -57.53447, 
        -57.54292, -57.54328, -57.53994, -57.53597, -57.53351, -57.53338, 
        -57.53505, -57.53784, -57.54052, -57.54285, -57.54383, -57.54359, 
        -57.543, -57.54316, -57.54421, -57.54935, -57.55836, -57.5717, 
        -57.58948, -57.6118, -57.63879, -57.67102, -57.70937, -57.75481, 
        -57.80869, -57.87178, -57.94445, -58.02599, -58.11496, -58.2099, 
        -58.30737, -58.40475, -58.4991, -58.58727, -58.66468, -58.73246, 
        -58.78812, -58.83133, -58.86156, -58.87861, -58.88249, -58.87307, 
        -58.8504, -58.81482, -58.76621, -58.70528, -58.6323, -58.54773, 
        -58.45207, -58.34662, -58.23235, -58.11137, -57.98517, -57.8556, 
        -57.72504, -57.59658, -57.47226, -57.35209, -57.23903, -57.13293, 
        -57.0347, -56.94471, -56.86201, -56.78627, -56.7165, -56.65278, 
        -56.59492, -56.54199, -56.49401, -56.45073, -56.41239, -56.37922, 
        -56.351, -56.32821, -56.31139, -56.3012, -56.29727, -56.29854, 
        -56.30409, -56.31247, -56.32181, -56.33026, -56.33376, -56.33112, 
        -56.31912, -56.29723, -56.26568, -56.22546, -56.17837, -56.12629, 
        -56.07118, -56.01415, -55.95597, -55.89762, -55.8384, -55.77865, 
        -55.71842, -55.65655, -55.5929, -55.5268, -55.45761, -55.38506, 
        -55.30795, -55.22613, -55.13924, -55.04729, -54.94975, -54.8461, 
        -54.73636, -54.62029, -54.50093, -54.37828, -54.25344, -54.12741, 
        -54.0015, -53.87704, -53.75529, -53.63683, -53.52154, -53.40977, 
        -53.30206, -53.19773, -53.09633, -52.99784, -52.90165, -52.80797, 
        -52.71592, -52.6244, -52.53284, -52.44062, -52.34813, -52.25584, 
        -52.16383, -52.07257, -51.9827, -51.89532, -51.81126, -51.73053, 
        -51.65431, -51.583, -51.51671, -51.45559, -51.39849, -51.34652, 
        -51.29784, -51.25248, -51.20932, -51.16928, -51.13089, -51.09451, 
        -51.05939, -51.02545, -50.99222, -50.95978, -50.92828, -50.89788, 
        -50.86901, -50.84304, -50.82162, -50.80563, -50.79658, -50.79559, 
        -50.80329, -50.82038, -50.84674, -50.88134, -50.92301, -50.96878, 
        -51.01611, -51.06215, -51.10474, -51.14201, -51.17362, -51.20014, 
        -51.22293, -51.24393, -51.26535, -51.28915, -51.31647, -51.34707, 
        -51.38023, -51.41437, -51.44776, -51.47764, -51.50463, -51.52696, 
        -51.54516, -51.56017, -51.57354, -51.58643, -51.59983, -51.61407, 
        -51.62941, -51.64547, -51.66251, -51.68109, -51.70165, -51.72499, 
        -51.75234,
  -40.65808, -40.82957, -40.9946, -41.16643, -41.32897, -41.49513, 
        -41.67762, -41.85186, -42.02171, -42.21324, -42.40602, -42.59981, 
        -42.79244, -42.98743, -43.18011, -43.38575, -43.59295, -43.80224, 
        -44.01519, -44.23343, -44.45784, -44.6871, -44.91903, -45.15205, 
        -45.38457, -45.61705, -45.84853, -46.07811, -46.30605, -46.53081, 
        -46.75081, -46.9656, -47.1748, -47.37802, -47.57516, -47.76571, 
        -47.94789, -48.12111, -48.28613, -48.44222, -48.59301, -48.73647, 
        -48.87355, -49.00421, -49.12873, -49.24789, -49.36295, -49.4762, 
        -49.58922, -49.70322, -49.81791, -49.93403, -50.05161, -50.17018, 
        -50.2894, -50.40744, -50.52676, -50.64664, -50.76718, -50.88905, 
        -51.01249, -51.1372, -51.26272, -51.3885, -51.51416, -51.63907, 
        -51.76297, -51.88685, -52.01212, -52.14014, -52.27157, -52.40769, 
        -52.54779, -52.69403, -52.84503, -53.00105, -53.16166, -53.32625, 
        -53.49473, -53.66698, -53.84333, -54.02369, -54.20913, -54.3989, 
        -54.59295, -54.79247, -54.9969, -55.20694, -55.4214, -55.6379, 
        -55.85284, -56.06412, -56.26649, -56.45508, -56.6255, -56.77361, 
        -56.8968, -56.99342, -57.06376, -57.11034, -57.13643, -57.14618, 
        -57.14406, -57.13471, -57.12283, -57.11118, -57.10215, -57.09628, 
        -57.09351, -57.09168, -57.09149, -57.09132, -57.09004, -57.0884, 
        -57.08656, -57.08552, -57.08624, -57.08955, -57.09656, -57.10738, 
        -57.12233, -57.14166, -57.16563, -57.19518, -57.23116, -57.27471, 
        -57.32733, -57.38941, -57.46133, -57.54118, -57.62938, -57.72275, 
        -57.81809, -57.91269, -58.00359, -58.0873, -58.16135, -58.22382, 
        -58.27424, -58.31178, -58.33649, -58.34799, -58.3463, -58.3316, 
        -58.30426, -58.26414, -58.21194, -58.14818, -58.07323, -57.98764, 
        -57.89185, -57.78569, -57.6728, -57.55259, -57.42683, -57.29741, 
        -57.16645, -57.03754, -56.91217, -56.79223, -56.67872, -56.57214, 
        -56.47421, -56.38432, -56.30249, -56.22779, -56.15953, -56.0979, 
        -56.04171, -55.99084, -55.9449, -55.90355, -55.86718, -55.83524, 
        -55.80833, -55.78514, -55.76817, -55.75751, -55.75169, -55.75034, 
        -55.75222, -55.75594, -55.76044, -55.76392, -55.76364, -55.75712, 
        -55.74289, -55.7195, -55.68704, -55.64661, -55.59973, -55.54807, 
        -55.49395, -55.43801, -55.38152, -55.32501, -55.26839, -55.21217, 
        -55.15556, -55.09831, -55.03953, -54.97769, -54.91457, -54.84792, 
        -54.77689, -54.70103, -54.61987, -54.53339, -54.44092, -54.34252, 
        -54.23806, -54.12838, -54.01464, -53.89768, -53.779, -53.65933, 
        -53.53997, -53.4221, -53.30662, -53.1942, -53.08456, -52.97773, 
        -52.87426, -52.77341, -52.6747, -52.57807, -52.48304, -52.38976, 
        -52.29758, -52.20569, -52.11378, -52.02161, -51.9286, -51.83684, 
        -51.74554, -51.65511, -51.56614, -51.47935, -51.39492, -51.31402, 
        -51.23674, -51.16416, -51.09677, -51.03441, -50.97734, -50.92512, 
        -50.87744, -50.83364, -50.79197, -50.75323, -50.71569, -50.67934, 
        -50.64341, -50.60759, -50.57195, -50.53646, -50.5021, -50.46942, 
        -50.43913, -50.41301, -50.39209, -50.37763, -50.37117, -50.373, 
        -50.38376, -50.40374, -50.43275, -50.46983, -50.51295, -50.55903, 
        -50.60694, -50.65323, -50.69575, -50.7331, -50.76458, -50.79132, 
        -50.81465, -50.8367, -50.85966, -50.88609, -50.91692, -50.95222, 
        -50.99072, -51.03084, -51.0706, -51.1078, -51.14091, -51.16903, 
        -51.19235, -51.21208, -51.22989, -51.24695, -51.2647, -51.28339, 
        -51.30332, -51.32421, -51.34615, -51.36938, -51.39397, -51.42118, 
        -51.45184,
  -40.39262, -40.55963, -40.73072, -40.89483, -41.0507, -41.21711, 
        -41.3853, -41.5449, -41.69901, -41.88657, -42.08836, -42.27844, 
        -42.46263, -42.65429, -42.84564, -43.04105, -43.24726, -43.45108, 
        -43.65639, -43.8649, -44.07917, -44.29652, -44.51643, -44.73732, 
        -44.95859, -45.17978, -45.40054, -45.62042, -45.83908, -46.0549, 
        -46.26644, -46.47293, -46.67429, -46.8702, -47.06004, -47.24447, 
        -47.42168, -47.59114, -47.75295, -47.90741, -48.05619, -48.19881, 
        -48.3352, -48.46605, -48.59117, -48.71117, -48.8277, -48.94255, 
        -49.05751, -49.17224, -49.28893, -49.40718, -49.52644, -49.64647, 
        -49.7666, -49.88665, -50.00703, -50.1286, -50.25138, -50.37601, 
        -50.50262, -50.63102, -50.76101, -50.89193, -51.02276, -51.15371, 
        -51.28275, -51.41282, -51.54507, -51.68024, -51.81976, -51.96384, 
        -52.11274, -52.2665, -52.42469, -52.58767, -52.75519, -52.92709, 
        -53.10289, -53.28278, -53.46723, -53.65644, -53.85048, -54.04963, 
        -54.25229, -54.46095, -54.67502, -54.89307, -55.11398, -55.33563, 
        -55.55418, -55.76584, -55.96604, -56.14986, -56.31308, -56.45201, 
        -56.56443, -56.6496, -56.70796, -56.74263, -56.75673, -56.75534, 
        -56.74208, -56.72376, -56.70393, -56.68489, -56.66928, -56.65778, 
        -56.65011, -56.64483, -56.64083, -56.63738, -56.6335, -56.6295, 
        -56.62569, -56.62263, -56.62134, -56.6228, -56.62761, -56.63605, 
        -56.64827, -56.66495, -56.68546, -56.71251, -56.74661, -56.78859, 
        -56.8399, -56.90088, -56.97175, -57.05111, -57.13744, -57.22831, 
        -57.32074, -57.41179, -57.49787, -57.57679, -57.64562, -57.70293, 
        -57.74821, -57.78064, -57.80052, -57.80726, -57.80098, -57.78103, 
        -57.74966, -57.70603, -57.65116, -57.58538, -57.50932, -57.42358, 
        -57.32884, -57.22545, -57.11438, -56.99651, -56.87251, -56.7447, 
        -56.61508, -56.48671, -56.36175, -56.24174, -56.12853, -56.0226, 
        -55.92522, -55.8361, -55.7549, -55.68134, -55.61349, -55.55313, 
        -55.4986, -55.44922, -55.4051, -55.36554, -55.33046, -55.2998, 
        -55.27337, -55.2516, -55.23447, -55.22249, -55.21463, -55.20972, 
        -55.20737, -55.20609, -55.20505, -55.20286, -55.19735, -55.18695, 
        -55.16953, -55.14442, -55.11127, -55.07103, -55.02503, -54.97352, 
        -54.92068, -54.86658, -54.81208, -54.75795, -54.70441, -54.65123, 
        -54.59828, -54.54477, -54.4905, -54.43463, -54.37662, -54.31537, 
        -54.24981, -54.17938, -54.10358, -54.02221, -53.93478, -53.84118, 
        -53.74206, -53.63797, -53.53004, -53.41911, -53.30673, -53.19392, 
        -53.08183, -52.97094, -52.86217, -52.7561, -52.65188, -52.55069, 
        -52.45185, -52.35497, -52.25937, -52.16489, -52.07142, -51.97837, 
        -51.88581, -51.79347, -51.70129, -51.60917, -51.51749, -51.42654, 
        -51.33609, -51.24678, -51.15882, -51.07259, -50.98855, -50.90714, 
        -50.82931, -50.75556, -50.68658, -50.62284, -50.56446, -50.51183, 
        -50.46394, -50.41995, -50.3787, -50.33914, -50.30063, -50.26215, 
        -50.2231, -50.18366, -50.14397, -50.10336, -50.06512, -50.0295, 
        -49.99775, -49.97142, -49.9515, -49.93937, -49.93603, -49.9417, 
        -49.95649, -49.98051, -50.013, -50.05301, -50.09835, -50.14679, 
        -50.19545, -50.24191, -50.28437, -50.32142, -50.35288, -50.3798, 
        -50.40387, -50.4272, -50.45215, -50.48083, -50.51531, -50.55481, 
        -50.59856, -50.64452, -50.69041, -50.73407, -50.77364, -50.80799, 
        -50.83702, -50.86173, -50.88427, -50.90575, -50.928, -50.95133, 
        -50.97595, -51.00177, -51.02866, -51.05698, -51.08698, -51.11953, 
        -51.15483,
  -40.14854, -40.30534, -40.46827, -40.63153, -40.79377, -40.94515, 
        -41.09573, -41.25726, -41.41185, -41.58513, -41.78286, -41.97047, 
        -42.15508, -42.34196, -42.5308, -42.71955, -42.91642, -43.11642, 
        -43.31532, -43.51719, -43.72066, -43.92711, -44.13422, -44.34294, 
        -44.55203, -44.76199, -44.97197, -45.18192, -45.39037, -45.59744, 
        -45.80043, -45.99893, -46.1924, -46.38107, -46.56551, -46.74457, 
        -46.91683, -47.08251, -47.24081, -47.3932, -47.53961, -47.68072, 
        -47.81681, -47.94788, -48.07264, -48.19398, -48.31208, -48.42883, 
        -48.54543, -48.66265, -48.78068, -48.90009, -49.02008, -49.14061, 
        -49.26054, -49.38073, -49.50152, -49.62383, -49.74824, -49.87475, 
        -50.00293, -50.13449, -50.26783, -50.40305, -50.53913, -50.67485, 
        -50.81045, -50.94678, -51.08493, -51.22672, -51.37272, -51.52378, 
        -51.67902, -51.83913, -52.00306, -52.17164, -52.34451, -52.52112, 
        -52.70297, -52.88924, -53.08076, -53.2776, -53.48035, -53.68816, 
        -53.9017, -54.12085, -54.34449, -54.57159, -54.80002, -55.02686, 
        -55.24839, -55.46045, -55.65854, -55.83743, -55.99363, -56.12257, 
        -56.22463, -56.29829, -56.34491, -56.36753, -56.37033, -56.35849, 
        -56.33686, -56.31008, -56.28268, -56.25705, -56.23519, -56.21865, 
        -56.20588, -56.19596, -56.18781, -56.18064, -56.17351, -56.16637, 
        -56.15977, -56.15333, -56.14966, -56.14885, -56.1514, -56.15746, 
        -56.16748, -56.18188, -56.20132, -56.22659, -56.25882, -56.29952, 
        -56.34951, -56.40932, -56.47832, -56.55575, -56.63939, -56.72686, 
        -56.81525, -56.90145, -56.98269, -57.05489, -57.11821, -57.17024, 
        -57.21038, -57.23825, -57.25395, -57.25708, -57.24738, -57.22468, 
        -57.19002, -57.14413, -57.08704, -57.02, -56.94363, -56.8588, 
        -56.76575, -56.66483, -56.55648, -56.44153, -56.32055, -56.19565, 
        -56.06852, -55.9421, -55.81735, -55.69902, -55.5873, -55.48274, 
        -55.38644, -55.29842, -55.21842, -55.14605, -55.08021, -55.02066, 
        -54.96723, -54.91902, -54.87625, -54.83759, -54.80329, -54.77345, 
        -54.74743, -54.72569, -54.70805, -54.69406, -54.68368, -54.67542, 
        -54.66873, -54.66235, -54.65467, -54.64687, -54.63647, -54.62177, 
        -54.60144, -54.57454, -54.54112, -54.50156, -54.45685, -54.40811, 
        -54.35705, -54.30505, -54.25318, -54.20155, -54.15054, -54.10001, 
        -54.05008, -53.99995, -53.94915, -53.89698, -53.84296, -53.78621, 
        -53.72548, -53.66006, -53.58901, -53.51223, -53.42976, -53.34132, 
        -53.24674, -53.14832, -53.04638, -52.94223, -52.83686, -52.73153, 
        -52.62695, -52.52366, -52.4223, -52.32318, -52.22665, -52.13167, 
        -52.0377, -51.94496, -51.85275, -51.76078, -51.66843, -51.57564, 
        -51.48277, -51.38999, -51.29746, -51.2053, -51.11415, -51.0238, 
        -50.93453, -50.84644, -50.75949, -50.6739, -50.59026, -50.50897, 
        -50.43073, -50.35577, -50.28445, -50.21923, -50.15948, -50.10549, 
        -50.05632, -50.01119, -49.96872, -49.92695, -49.8852, -49.84281, 
        -49.7988, -49.75355, -49.70814, -49.66323, -49.62037, -49.58113, 
        -49.54779, -49.52137, -49.50309, -49.49394, -49.49454, -49.50485, 
        -49.52463, -49.55354, -49.59026, -49.6336, -49.68208, -49.73172, 
        -49.78157, -49.82819, -49.87029, -49.90703, -49.9385, -49.96559, 
        -49.99046, -50.01517, -50.04201, -50.0734, -50.11105, -50.15488, 
        -50.20248, -50.25358, -50.30555, -50.35555, -50.40179, -50.44257, 
        -50.47783, -50.50838, -50.53602, -50.56244, -50.58919, -50.61696, 
        -50.6462, -50.67707, -50.70961, -50.74418, -50.78097, -50.82084, 
        -50.86459,
  -39.91027, -40.06721, -40.2302, -40.3947, -40.56833, -40.7236, 
        -40.87006, -41.00624, -41.14801, -41.31484, -41.49144, -41.68075, 
        -41.86366, -42.04787, -42.23414, -42.41948, -42.60495, -42.79636, 
        -42.99013, -43.18545, -43.37998, -43.57487, -43.77101, -43.96727, 
        -44.16536, -44.36444, -44.56456, -44.76484, -44.96463, -45.16306, 
        -45.35796, -45.54845, -45.73453, -45.91643, -46.09465, -46.26779, 
        -46.43521, -46.59703, -46.75113, -46.90098, -47.04575, -47.18546, 
        -47.32098, -47.45242, -47.57909, -47.7019, -47.8219, -47.94035, 
        -48.05845, -48.1768, -48.29579, -48.41575, -48.53593, -48.65554, 
        -48.77375, -48.89329, -49.01369, -49.13599, -49.26104, -49.38877, 
        -49.51941, -49.65331, -49.78952, -49.92799, -50.06804, -50.20824, 
        -50.34883, -50.49016, -50.63368, -50.78033, -50.93209, -51.08765, 
        -51.24804, -51.41261, -51.58118, -51.75447, -51.93171, -52.1133, 
        -52.29999, -52.4917, -52.689, -52.89269, -53.10318, -53.32039, 
        -53.54408, -53.77367, -54.00795, -54.24462, -54.48075, -54.71178, 
        -54.93615, -55.14828, -55.34353, -55.51729, -55.66618, -55.78687, 
        -55.87815, -55.94025, -55.97511, -55.98591, -55.97749, -55.95552, 
        -55.92493, -55.89044, -55.85606, -55.82461, -55.79755, -55.77575, 
        -55.75734, -55.74286, -55.73058, -55.71955, -55.70869, -55.69817, 
        -55.68834, -55.68, -55.67383, -55.67066, -55.67083, -55.67488, 
        -55.68306, -55.6957, -55.71337, -55.73717, -55.76812, -55.80756, 
        -55.85632, -55.91453, -55.98078, -56.05546, -56.13559, -56.21864, 
        -56.30193, -56.38237, -56.45763, -56.52496, -56.58242, -56.6289, 
        -56.66415, -56.6882, -56.70063, -56.70071, -56.68818, -56.66306, 
        -56.626, -56.57768, -56.51935, -56.45184, -56.37552, -56.29214, 
        -56.20046, -56.10266, -55.99769, -55.88587, -55.76888, -55.64782, 
        -55.52489, -55.4015, -55.28059, -55.16489, -55.05568, -54.95372, 
        -54.85918, -54.77227, -54.69389, -54.62246, -54.55771, -54.49891, 
        -54.4457, -54.39843, -54.35601, -54.31814, -54.28423, -54.25311, 
        -54.2274, -54.20507, -54.18639, -54.17065, -54.15709, -54.14563, 
        -54.13483, -54.12391, -54.11227, -54.09925, -54.08434, -54.06605, 
        -54.0436, -54.01554, -53.98188, -53.94324, -53.90018, -53.85372, 
        -53.80507, -53.75522, -53.70594, -53.65673, -53.60837, -53.55963, 
        -53.51162, -53.46364, -53.4144, -53.3652, -53.31414, -53.26039, 
        -53.20363, -53.14223, -53.0756, -53.00333, -52.9255, -52.84267, 
        -52.75496, -52.66314, -52.56782, -52.47058, -52.37316, -52.2756, 
        -52.17918, -52.08423, -51.99047, -51.89889, -51.80887, -51.72014, 
        -51.63155, -51.54271, -51.45391, -51.36407, -51.27299, -51.18068, 
        -51.08715, -50.99382, -50.90027, -50.80817, -50.71741, -50.62791, 
        -50.53969, -50.45274, -50.36683, -50.28215, -50.19879, -50.11774, 
        -50.03905, -49.96381, -49.89227, -49.82548, -49.76428, -49.70837, 
        -49.65744, -49.61007, -49.56461, -49.51914, -49.4721, -49.4235, 
        -49.37315, -49.32113, -49.26887, -49.21783, -49.16988, -49.12699, 
        -49.09156, -49.06524, -49.04915, -49.04343, -49.04876, -49.06421, 
        -49.08971, -49.124, -49.16557, -49.21206, -49.26299, -49.31485, 
        -49.36511, -49.41207, -49.45361, -49.48988, -49.52103, -49.54861, 
        -49.57429, -49.60062, -49.63002, -49.66428, -49.70494, -49.75263, 
        -49.80557, -49.86181, -49.91929, -49.97535, -50.02787, -50.07515, 
        -50.11688, -50.15359, -50.18702, -50.2187, -50.25023, -50.28265, 
        -50.31696, -50.35345, -50.39243, -50.43423, -50.47907, -50.52768, 
        -50.58156,
  -39.72095, -39.8871, -40.04176, -40.1939, -40.35868, -40.51157, 
        -40.64714, -40.78918, -40.93609, -41.08935, -41.23466, -41.39913, 
        -41.58303, -41.76903, -41.95151, -42.13108, -42.31145, -42.4907, 
        -42.67618, -42.86528, -43.05341, -43.23942, -43.42541, -43.61251, 
        -43.80058, -43.99005, -44.18092, -44.37185, -44.56264, -44.75237, 
        -44.93933, -45.1222, -45.30124, -45.47583, -45.64797, -45.81618, 
        -45.97941, -46.13703, -46.28932, -46.43668, -46.5793, -46.71793, 
        -46.85294, -46.98444, -47.11203, -47.23645, -47.35817, -47.47837, 
        -47.59766, -47.71573, -47.83511, -47.95494, -48.07448, -48.19299, 
        -48.31101, -48.42916, -48.54856, -48.67024, -48.79504, -48.92325, 
        -49.05466, -49.18946, -49.32811, -49.46901, -49.61169, -49.75438, 
        -49.89865, -50.04399, -50.1919, -50.34327, -50.49875, -50.65851, 
        -50.82291, -50.99141, -51.16339, -51.33978, -51.52028, -51.70547, 
        -51.89576, -52.09149, -52.29385, -52.50364, -52.72166, -52.94681, 
        -53.18105, -53.42199, -53.66726, -53.91343, -54.15677, -54.39407, 
        -54.62102, -54.83244, -55.02411, -55.19194, -55.33275, -55.44357, 
        -55.52381, -55.57406, -55.59673, -55.59561, -55.57581, -55.54271, 
        -55.50348, -55.46182, -55.42136, -55.38435, -55.35307, -55.32692, 
        -55.30508, -55.28646, -55.27021, -55.25528, -55.24069, -55.22667, 
        -55.21357, -55.20223, -55.19341, -55.18789, -55.18612, -55.1884, 
        -55.19516, -55.20558, -55.22219, -55.24501, -55.27499, -55.31345, 
        -55.36092, -55.41728, -55.48211, -55.55349, -55.62932, -55.70716, 
        -55.78438, -55.85834, -55.92691, -55.98804, -56.03958, -56.08078, 
        -56.11107, -56.13125, -56.14069, -56.13842, -56.12259, -56.09587, 
        -56.05718, -56.00772, -55.94821, -55.88062, -55.8055, -55.72373, 
        -55.63557, -55.54075, -55.43956, -55.33189, -55.21935, -55.10326, 
        -54.98463, -54.86595, -54.7494, -54.63773, -54.53189, -54.43275, 
        -54.34109, -54.25682, -54.17981, -54.10847, -54.04418, -53.98606, 
        -53.93331, -53.8862, -53.84401, -53.80577, -53.77186, -53.74174, 
        -53.71524, -53.69187, -53.67143, -53.65357, -53.63761, -53.62297, 
        -53.60857, -53.5936, -53.57785, -53.56091, -53.54228, -53.52131, 
        -53.49688, -53.46868, -53.4356, -53.39844, -53.35671, -53.31276, 
        -53.26677, -53.21962, -53.17223, -53.12495, -53.07802, -53.03098, 
        -52.98402, -52.93718, -52.89014, -52.84233, -52.79329, -52.74213, 
        -52.68802, -52.62988, -52.56697, -52.49932, -52.42672, -52.34958, 
        -52.26822, -52.18306, -52.09538, -52.00594, -51.9164, -51.82711, 
        -51.73886, -51.65218, -51.56646, -51.4813, -51.39797, -51.31497, 
        -51.23174, -51.14713, -51.06118, -50.97331, -50.88332, -50.79146, 
        -50.69817, -50.60448, -50.51163, -50.41982, -50.32942, -50.24095, 
        -50.1539, -50.06792, -49.98276, -49.89894, -49.81641, -49.73557, 
        -49.65705, -49.58099, -49.50866, -49.44066, -49.3776, -49.31961, 
        -49.266, -49.21496, -49.16517, -49.11474, -49.06179, -49.00556, 
        -48.94733, -48.88674, -48.82713, -48.7697, -48.71689, -48.67076, 
        -48.63382, -48.60781, -48.5942, -48.59216, -48.60232, -48.62325, 
        -48.65434, -48.6941, -48.74076, -48.79226, -48.8459, -48.89949, 
        -48.9503, -48.99682, -49.03806, -49.07389, -49.10512, -49.13271, 
        -49.15946, -49.18709, -49.21881, -49.25596, -49.2997, -49.35094, 
        -49.40808, -49.46923, -49.5319, -49.59354, -49.65178, -49.70545, 
        -49.75351, -49.79671, -49.83613, -49.87346, -49.91032, -49.94818, 
        -49.98816, -50.03114, -50.07737, -50.12637, -50.18041, -50.23951, 
        -50.30503,
  -39.56799, -39.72282, -39.87447, -40.01954, -40.17156, -40.30766, 
        -40.44985, -40.58891, -40.73164, -40.86941, -41.00115, -41.1364, 
        -41.31062, -41.49582, -41.67725, -41.849, -42.02582, -42.20185, 
        -42.37689, -42.56068, -42.74172, -42.92184, -43.09879, -43.27741, 
        -43.45694, -43.63805, -43.82002, -44.00147, -44.18377, -44.36516, 
        -44.54448, -44.7207, -44.89352, -45.06331, -45.23008, -45.39341, 
        -45.55233, -45.70642, -45.85585, -46.00064, -46.14171, -46.27911, 
        -46.41365, -46.5441, -46.67245, -46.79799, -46.92127, -47.04255, 
        -47.16263, -47.28201, -47.40123, -47.52044, -47.63885, -47.75594, 
        -47.87247, -47.98909, -48.10714, -48.22795, -48.35189, -48.47864, 
        -48.61024, -48.74561, -48.88473, -49.02699, -49.17164, -49.31742, 
        -49.46414, -49.61259, -49.76332, -49.91737, -50.07569, -50.23845, 
        -50.40535, -50.57593, -50.7502, -50.92881, -51.11065, -51.29819, 
        -51.49127, -51.69048, -51.89722, -52.11284, -52.33803, -52.5731, 
        -52.81769, -53.06963, -53.32533, -53.58083, -53.83168, -54.07371, 
        -54.30237, -54.51252, -54.70008, -54.86157, -54.99257, -55.09292, 
        -55.16127, -55.19905, -55.20906, -55.19554, -55.16441, -55.12208, 
        -55.07403, -55.02527, -54.97935, -54.93773, -54.90234, -54.87242, 
        -54.84707, -54.82488, -54.80498, -54.78648, -54.7684, -54.75111, 
        -54.73392, -54.71984, -54.70852, -54.70081, -54.69741, -54.69857, 
        -54.7042, -54.71489, -54.73104, -54.75325, -54.78252, -54.8201, 
        -54.86606, -54.92047, -54.98216, -55.04966, -55.12058, -55.19258, 
        -55.26316, -55.33019, -55.39095, -55.44509, -55.4905, -55.5265, 
        -55.55283, -55.56944, -55.57602, -55.57146, -55.55524, -55.52697, 
        -55.48718, -55.43686, -55.37719, -55.30981, -55.23584, -55.15594, 
        -55.07061, -54.97941, -54.88242, -54.77951, -54.67185, -54.56094, 
        -54.44706, -54.33403, -54.22278, -54.11545, -54.01391, -53.9188, 
        -53.83052, -53.74876, -53.67341, -53.60431, -53.5409, -53.48329, 
        -53.43064, -53.38323, -53.34061, -53.30222, -53.26802, -53.23716, 
        -53.20956, -53.18488, -53.16284, -53.14301, -53.12453, -53.10689, 
        -53.08932, -53.07014, -53.05123, -53.03126, -53.00994, -52.98725, 
        -52.96215, -52.93421, -52.90261, -52.86754, -52.82927, -52.78825, 
        -52.74531, -52.70075, -52.65548, -52.60986, -52.56376, -52.5175, 
        -52.47092, -52.42405, -52.37729, -52.3302, -52.28244, -52.23264, 
        -52.18024, -52.12484, -52.06573, -52.00267, -51.93441, -51.86307, 
        -51.78813, -51.71022, -51.63039, -51.54917, -51.46762, -51.38659, 
        -51.3065, -51.22762, -51.1496, -51.07232, -50.9953, -50.91781, 
        -50.83928, -50.75846, -50.67505, -50.58919, -50.50042, -50.40934, 
        -50.31633, -50.22276, -50.12983, -50.03865, -49.9492, -49.86156, 
        -49.77552, -49.69064, -49.60656, -49.52348, -49.44182, -49.36145, 
        -49.28202, -49.20586, -49.13279, -49.06331, -48.99819, -48.93752, 
        -48.88056, -48.82518, -48.77023, -48.71289, -48.65288, -48.58888, 
        -48.5225, -48.4552, -48.38906, -48.32613, -48.26937, -48.22131, 
        -48.18391, -48.15896, -48.14771, -48.14975, -48.16431, -48.19005, 
        -48.2262, -48.27066, -48.32146, -48.37635, -48.4324, -48.48703, 
        -48.53813, -48.58423, -48.6249, -48.66003, -48.69099, -48.71881, 
        -48.74623, -48.77557, -48.80915, -48.84885, -48.89468, -48.94931, 
        -49.01046, -49.07616, -49.14341, -49.21006, -49.27383, -49.33334, 
        -49.38764, -49.43729, -49.48299, -49.52636, -49.56923, -49.61327, 
        -49.65982, -49.71019, -49.76484, -49.82402, -49.88862, -49.95936, 
        -50.03819,
  -39.42449, -39.56975, -39.71602, -39.85746, -39.99775, -40.12155, 
        -40.26485, -40.39588, -40.53308, -40.66032, -40.78326, -40.90926, 
        -41.0672, -41.23558, -41.4158, -41.57233, -41.74792, -41.92532, 
        -42.09827, -42.27235, -42.44748, -42.62193, -42.79098, -42.96066, 
        -43.13277, -43.30613, -43.48058, -43.65521, -43.82972, -44.00339, 
        -44.17597, -44.34568, -44.51291, -44.67765, -44.83989, -44.99871, 
        -45.15385, -45.30372, -45.45065, -45.59335, -45.73259, -45.86934, 
        -46.00298, -46.13438, -46.26297, -46.38903, -46.51294, -46.63456, 
        -46.7547, -46.87398, -46.99261, -47.11075, -47.22764, -47.34336, 
        -47.45729, -47.5724, -47.68919, -47.80876, -47.9317, -48.05852, 
        -48.18942, -48.32443, -48.46356, -48.60587, -48.75089, -48.8976, 
        -49.04585, -49.19589, -49.34824, -49.50375, -49.66251, -49.82654, 
        -49.99445, -50.16628, -50.34198, -50.52171, -50.70634, -50.89564, 
        -51.0909, -51.29299, -51.50362, -51.72458, -51.95668, -52.20058, 
        -52.45496, -52.71705, -52.98272, -53.24702, -53.50372, -53.7499, 
        -53.97956, -54.18803, -54.37115, -54.52563, -54.6483, -54.73748, 
        -54.7935, -54.81811, -54.81475, -54.78828, -54.74526, -54.69246, 
        -54.63589, -54.57993, -54.52845, -54.48312, -54.44442, -54.41039, 
        -54.38202, -54.35691, -54.33414, -54.31247, -54.29136, -54.27126, 
        -54.25248, -54.23603, -54.22254, -54.21317, -54.20854, -54.20868, 
        -54.21398, -54.22446, -54.24025, -54.26213, -54.29095, -54.32735, 
        -54.37172, -54.42253, -54.4808, -54.54382, -54.60936, -54.67511, 
        -54.73887, -54.79861, -54.8531, -54.90039, -54.93968, -54.97063, 
        -54.99285, -55.00618, -55.01013, -55.00357, -54.98571, -54.95636, 
        -54.91597, -54.86538, -54.80592, -54.73922, -54.66567, -54.58829, 
        -54.50605, -54.41874, -54.32595, -54.22817, -54.12622, -54.0213, 
        -53.91472, -53.80769, -53.70241, -53.60067, -53.50394, -53.41319, 
        -53.32808, -53.24907, -53.17599, -53.10816, -53.04567, -52.98814, 
        -52.93568, -52.88814, -52.84505, -52.80621, -52.77003, -52.73833, 
        -52.70964, -52.68358, -52.65988, -52.63777, -52.61695, -52.59689, 
        -52.57688, -52.55629, -52.5349, -52.51278, -52.49014, -52.46672, 
        -52.44186, -52.41484, -52.38536, -52.35305, -52.31775, -52.27999, 
        -52.23988, -52.19802, -52.15488, -52.11073, -52.06561, -52.01945, 
        -51.97158, -51.92456, -51.87762, -51.83066, -51.78305, -51.73421, 
        -51.68365, -51.63071, -51.57502, -51.51605, -51.45385, -51.38858, 
        -51.32046, -51.24978, -51.17731, -51.1041, -51.03046, -50.95738, 
        -50.88485, -50.81296, -50.74179, -50.67082, -50.5994, -50.52655, 
        -50.45182, -50.37428, -50.29339, -50.20924, -50.1219, -50.03168, 
        -49.93859, -49.84578, -49.7537, -49.66357, -49.57533, -49.48888, 
        -49.40411, -49.32041, -49.23749, -49.15541, -49.07436, -48.99485, 
        -48.91682, -48.84053, -48.76649, -48.69577, -48.62849, -48.56463, 
        -48.5031, -48.44248, -48.38099, -48.31689, -48.24905, -48.17774, 
        -48.10376, -48.02975, -47.95824, -47.89156, -47.83258, -47.78399, 
        -47.74764, -47.72493, -47.71648, -47.72226, -47.74088, -47.7709, 
        -47.80961, -47.85757, -47.91133, -47.96811, -48.02539, -48.08053, 
        -48.13115, -48.17634, -48.21578, -48.25023, -48.28072, -48.30852, 
        -48.33638, -48.36675, -48.40198, -48.44382, -48.49339, -48.55113, 
        -48.61592, -48.68562, -48.75745, -48.82888, -48.89795, -48.96295, 
        -49.02308, -49.07884, -49.13098, -49.18077, -49.23037, -49.28117, 
        -49.33529, -49.39423, -49.45833, -49.52813, -49.60421, -49.68782, 
        -49.78097,
  -39.29163, -39.43023, -39.5675, -39.70393, -39.8268, -39.95369, 
        -40.0898, -40.21325, -40.34229, -40.46042, -40.58466, -40.70225, 
        -40.84492, -41.00734, -41.16883, -41.31024, -41.47823, -41.6572, 
        -41.83249, -42.00368, -42.17163, -42.33768, -42.50135, -42.66396, 
        -42.82872, -42.99571, -43.1633, -43.33112, -43.49897, -43.666, 
        -43.83236, -43.99712, -44.15853, -44.31856, -44.47651, -44.63155, 
        -44.78296, -44.93077, -45.075, -45.21618, -45.35414, -45.48951, 
        -45.62257, -45.75333, -45.88175, -46.00774, -46.13136, -46.25254, 
        -46.3712, -46.48975, -46.60738, -46.72409, -46.83953, -46.95384, 
        -47.06737, -47.18117, -47.29666, -47.41486, -47.5365, -47.66206, 
        -47.79189, -47.92603, -48.06388, -48.20535, -48.34846, -48.49524, 
        -48.64323, -48.79371, -48.94624, -49.10234, -49.26247, -49.42655, 
        -49.59472, -49.76691, -49.94297, -50.12342, -50.30863, -50.49915, 
        -50.69621, -50.90086, -51.11512, -51.3409, -51.57847, -51.83006, 
        -52.09324, -52.3644, -52.63881, -52.9108, -53.17447, -53.42436, 
        -53.65501, -53.86148, -54.03992, -54.18702, -54.29997, -54.37761, 
        -54.42049, -54.43121, -54.4137, -54.37366, -54.31712, -54.25368, 
        -54.1882, -54.1255, -54.06886, -54.02008, -53.97834, -53.94319, 
        -53.91262, -53.88519, -53.85991, -53.83572, -53.81216, -53.78981, 
        -53.76926, -53.75104, -53.7362, -53.72564, -53.72018, -53.71986, 
        -53.72403, -53.73449, -53.75028, -53.77207, -53.8002, -53.83529, 
        -53.87754, -53.92646, -53.9808, -54.03893, -54.09871, -54.15793, 
        -54.21463, -54.26731, -54.31451, -54.35509, -54.38871, -54.41473, 
        -54.43301, -54.4432, -54.44445, -54.43468, -54.4154, -54.38514, 
        -54.34457, -54.29416, -54.23545, -54.16993, -54.09926, -54.0247, 
        -53.94576, -53.86215, -53.77433, -53.68222, -53.5864, -53.48798, 
        -53.38793, -53.28782, -53.18916, -53.09303, -53.00128, -52.9142, 
        -52.83271, -52.75534, -52.68416, -52.61779, -52.55611, -52.49907, 
        -52.44683, -52.39934, -52.35585, -52.31619, -52.28047, -52.24762, 
        -52.21778, -52.19032, -52.16474, -52.14079, -52.11791, -52.09565, 
        -52.07362, -52.0511, -52.0282, -52.00486, -51.98171, -51.95831, 
        -51.93442, -51.90976, -51.88279, -51.85244, -51.82038, -51.78578, 
        -51.74873, -51.70974, -51.66903, -51.6264, -51.58211, -51.53645, 
        -51.48964, -51.44245, -51.39539, -51.34836, -51.30126, -51.25333, 
        -51.20425, -51.15347, -51.10063, -51.04576, -50.98846, -50.92893, 
        -50.86709, -50.80299, -50.73767, -50.67174, -50.60538, -50.53922, 
        -50.47321, -50.40651, -50.34086, -50.27506, -50.20807, -50.13909, 
        -50.06744, -49.9926, -49.914, -49.83154, -49.74555, -49.65694, 
        -49.56641, -49.47548, -49.38493, -49.29631, -49.20996, -49.12527, 
        -49.04216, -48.95995, -48.87822, -48.79721, -48.71724, -48.6385, 
        -48.5609, -48.48443, -48.40948, -48.33703, -48.26713, -48.19971, 
        -48.13322, -48.06672, -47.9982, -47.92676, -47.85155, -47.77203, 
        -47.69207, -47.61324, -47.53839, -47.47036, -47.41159, -47.36455, 
        -47.33099, -47.3116, -47.30683, -47.31594, -47.33781, -47.37085, 
        -47.41306, -47.46259, -47.51746, -47.57444, -47.6314, -47.68551, 
        -47.73468, -47.77859, -47.81666, -47.84991, -47.8795, -47.90691, 
        -47.93492, -47.96562, -48.00167, -48.04501, -48.09694, -48.15736, 
        -48.22547, -48.29912, -48.37546, -48.4517, -48.52557, -48.59552, 
        -48.66127, -48.72285, -48.78124, -48.83757, -48.89423, -48.95287, 
        -49.01458, -49.08297, -49.15765, -49.23909, -49.3278, -49.42527, 
        -49.5333,
  -39.15631, -39.29534, -39.428, -39.55516, -39.68092, -39.8078, 
        -39.92752, -40.03995, -40.16328, -40.27744, -40.38161, -40.49319, 
        -40.61905, -40.78126, -40.93473, -41.0613, -41.22609, -41.40231, 
        -41.5747, -41.74181, -41.90658, -42.06748, -42.2262, -42.38398, 
        -42.54337, -42.70372, -42.86525, -43.02665, -43.18912, -43.35079, 
        -43.51219, -43.67186, -43.8301, -43.98652, -44.1408, -44.29276, 
        -44.44101, -44.58613, -44.72829, -44.86736, -45.00375, -45.13825, 
        -45.26944, -45.39905, -45.52663, -45.65163, -45.77419, -45.89417, 
        -46.01247, -46.13002, -46.24649, -46.36162, -46.47569, -46.58865, 
        -46.70107, -46.81387, -46.92806, -47.04468, -47.1638, -47.28757, 
        -47.41565, -47.54834, -47.6847, -47.82373, -47.9663, -48.11138, 
        -48.25814, -48.40805, -48.5601, -48.7164, -48.87585, -49.03881, 
        -49.20691, -49.37895, -49.55478, -49.73531, -49.91979, -50.11103, 
        -50.30938, -50.51611, -50.7336, -50.9639, -51.20788, -51.46606, 
        -51.73634, -52.01479, -52.29624, -52.57458, -52.84335, -53.09624, 
        -53.32729, -53.5316, -53.70546, -53.84484, -53.94695, -54.01246, 
        -54.04165, -54.03786, -54.0056, -53.95156, -53.8833, -53.80874, 
        -53.73405, -53.66487, -53.60362, -53.5514, -53.50744, -53.47049, 
        -53.43838, -53.40933, -53.38224, -53.35611, -53.33083, -53.30605, 
        -53.28421, -53.26511, -53.24963, -53.2387, -53.23285, -53.23289, 
        -53.23795, -53.24856, -53.26438, -53.28601, -53.31329, -53.34684, 
        -53.38652, -53.43189, -53.48176, -53.53471, -53.58851, -53.64116, 
        -53.69102, -53.7357, -53.77605, -53.81044, -53.83846, -53.86015, 
        -53.87434, -53.88136, -53.88019, -53.86913, -53.84866, -53.81757, 
        -53.77694, -53.72739, -53.66983, -53.60647, -53.53821, -53.46627, 
        -53.39088, -53.31152, -53.22893, -53.14227, -53.05305, -52.96025, 
        -52.86742, -52.77467, -52.68254, -52.59149, -52.50441, -52.42119, 
        -52.34277, -52.26876, -52.19892, -52.1338, -52.07314, -52.01702, 
        -51.96506, -51.91727, -51.87344, -51.83352, -51.79707, -51.76304, 
        -51.7318, -51.7031, -51.67612, -51.65059, -51.62595, -51.6019, 
        -51.57702, -51.55325, -51.52939, -51.50569, -51.4827, -51.46022, 
        -51.43845, -51.41595, -51.39152, -51.36525, -51.33659, -51.30555, 
        -51.27197, -51.23573, -51.19727, -51.15672, -51.11403, -51.06945, 
        -51.0234, -50.97653, -50.92999, -50.8836, -50.83741, -50.79066, 
        -50.74305, -50.69444, -50.64454, -50.59237, -50.53942, -50.48468, 
        -50.4284, -50.37043, -50.31138, -50.25145, -50.19138, -50.13085, 
        -50.0704, -50.00967, -49.94834, -49.8864, -49.8229, -49.75681, 
        -49.68769, -49.61472, -49.53808, -49.45743, -49.37335, -49.28701, 
        -49.19912, -49.11065, -49.02276, -48.93652, -48.85274, -48.77046, 
        -48.68908, -48.60869, -48.52872, -48.44911, -48.36908, -48.29074, 
        -48.21359, -48.13686, -48.06122, -47.98711, -47.91449, -47.84254, 
        -47.77079, -47.69801, -47.62238, -47.54339, -47.46121, -47.377, 
        -47.29305, -47.21143, -47.136, -47.06926, -47.01329, -46.97019, 
        -46.94114, -46.92642, -46.92549, -46.93802, -46.96229, -46.99689, 
        -47.03995, -47.08942, -47.14331, -47.19865, -47.25331, -47.30526, 
        -47.35199, -47.39349, -47.42991, -47.46154, -47.48982, -47.5166, 
        -47.54396, -47.57373, -47.60993, -47.65417, -47.70765, -47.77031, 
        -47.84149, -47.91874, -47.99933, -48.08011, -48.15864, -48.23352, 
        -48.30437, -48.37157, -48.43599, -48.49913, -48.56321, -48.63026, 
        -48.70249, -48.78117, -48.86733, -48.96117, -49.0635, -49.17567, 
        -49.29923,
  -39.04449, -39.15288, -39.28187, -39.41392, -39.54282, -39.66291, 
        -39.77444, -39.88819, -39.99413, -40.09409, -40.19621, -40.3049, 
        -40.42929, -40.57549, -40.71402, -40.83659, -41.00264, -41.16549, 
        -41.32945, -41.49088, -41.64896, -41.80515, -41.96041, -42.11766, 
        -42.27396, -42.42958, -42.58463, -42.74197, -42.90007, -43.05791, 
        -43.21532, -43.37137, -43.52601, -43.67913, -43.83082, -43.97972, 
        -44.12561, -44.26767, -44.40783, -44.54499, -44.67996, -44.81292, 
        -44.94351, -45.07186, -45.19796, -45.32146, -45.4421, -45.56058, 
        -45.6773, -45.7934, -45.90818, -46.02208, -46.13495, -46.2459, 
        -46.35721, -46.4689, -46.58165, -46.69642, -46.81434, -46.93578, 
        -47.06145, -47.19151, -47.32521, -47.46258, -47.60218, -47.74414, 
        -47.88945, -48.03802, -48.18888, -48.34391, -48.5014, -48.6642, 
        -48.83166, -49.00264, -49.17837, -49.35859, -49.54413, -49.73582, 
        -49.93512, -50.14373, -50.3635, -50.5973, -50.84564, -51.10897, 
        -51.38435, -51.668, -51.95484, -52.23693, -52.50932, -52.76432, 
        -52.99538, -53.19726, -53.36614, -53.49786, -53.59082, -53.64383, 
        -53.65904, -53.64033, -53.59287, -53.52428, -53.44307, -53.3573, 
        -53.27388, -53.19787, -53.13229, -53.07707, -53.03015, -52.99212, 
        -52.959, -52.92892, -52.90056, -52.8732, -52.84682, -52.82222, 
        -52.79998, -52.78091, -52.76553, -52.75493, -52.74974, -52.75018, 
        -52.75565, -52.76678, -52.78275, -52.80371, -52.82966, -52.86099, 
        -52.8967, -52.93815, -52.98312, -53.03049, -53.0783, -53.12461, 
        -53.16792, -53.20708, -53.24125, -53.26991, -53.29279, -53.30998, 
        -53.3209, -53.32429, -53.32037, -53.30769, -53.28569, -53.25481, 
        -53.21462, -53.16614, -53.11092, -53.04939, -52.98412, -52.91497, 
        -52.84263, -52.76778, -52.69003, -52.60975, -52.52656, -52.44197, 
        -52.35605, -52.26977, -52.1837, -52.09898, -52.01593, -51.93589, 
        -51.85983, -51.78757, -51.71919, -51.65498, -51.59531, -51.53985, 
        -51.48854, -51.44087, -51.39688, -51.35563, -51.31826, -51.28375, 
        -51.25149, -51.22159, -51.19354, -51.16661, -51.14046, -51.11487, 
        -51.08952, -51.06492, -51.04083, -51.01724, -50.99494, -50.97383, 
        -50.9539, -50.93358, -50.91228, -50.88955, -50.86436, -50.83654, 
        -50.80618, -50.7731, -50.73718, -50.6988, -50.65842, -50.61475, 
        -50.57074, -50.52568, -50.48048, -50.43576, -50.39106, -50.34622, 
        -50.30061, -50.25421, -50.2071, -50.15903, -50.10996, -50.05945, 
        -50.00764, -49.95464, -49.90033, -49.84534, -49.78997, -49.73383, 
        -49.6775, -49.62026, -49.56242, -49.5033, -49.44217, -49.37831, 
        -49.3112, -49.24011, -49.16528, -49.08691, -49.00536, -48.92094, 
        -48.83623, -48.75137, -48.66689, -48.58393, -48.50306, -48.42383, 
        -48.34496, -48.26647, -48.18842, -48.11031, -48.03242, -47.95469, 
        -47.87762, -47.80076, -47.72415, -47.64819, -47.57237, -47.49608, 
        -47.41879, -47.33927, -47.25667, -47.1708, -47.08292, -46.99493, 
        -46.90866, -46.82686, -46.75372, -46.69054, -46.63976, -46.60262, 
        -46.57959, -46.57031, -46.57362, -46.58917, -46.61429, -46.64942, 
        -46.69177, -46.73949, -46.79081, -46.84298, -46.89431, -46.94214, 
        -46.98592, -47.02438, -47.05809, -47.08768, -47.1144, -47.13985, 
        -47.16641, -47.19647, -47.23279, -47.27767, -47.33231, -47.39685, 
        -47.47029, -47.55061, -47.63477, -47.71928, -47.80211, -47.8816, 
        -47.95769, -48.03012, -48.10093, -48.17101, -48.24307, -48.31909, 
        -48.40151, -48.49124, -48.58956, -48.69675, -48.81375, -48.94114, 
        -49.08028,
  -38.92872, -39.03909, -39.14799, -39.27561, -39.40818, -39.52414, 
        -39.63467, -39.73834, -39.83266, -39.92363, -40.03235, -40.14717, 
        -40.26124, -40.388, -40.50651, -40.6343, -40.77571, -40.93321, 
        -41.09091, -41.24586, -41.39681, -41.55464, -41.70825, -41.86583, 
        -42.02105, -42.17263, -42.32457, -42.47687, -42.63022, -42.78487, 
        -42.93939, -43.09147, -43.24295, -43.39358, -43.54294, -43.69024, 
        -43.83407, -43.97514, -44.11345, -44.2494, -44.38278, -44.514, 
        -44.64292, -44.76949, -44.89364, -45.01484, -45.13319, -45.24851, 
        -45.36362, -45.47774, -45.59098, -45.70369, -45.81547, -45.92646, 
        -46.037, -46.14715, -46.25789, -46.3704, -46.48563, -46.60417, 
        -46.72683, -46.85358, -46.9841, -47.11763, -47.25313, -47.39297, 
        -47.53595, -47.68221, -47.83202, -47.98567, -48.14302, -48.30529, 
        -48.47187, -48.64272, -48.81747, -48.99761, -49.18301, -49.37402, 
        -49.57382, -49.78383, -50.00577, -50.24077, -50.49222, -50.75844, 
        -51.03695, -51.32378, -51.61372, -51.89976, -52.17433, -52.43027, 
        -52.66064, -52.85958, -53.02279, -53.14649, -53.22909, -53.26984, 
        -53.27103, -53.23717, -53.17443, -53.09036, -52.99591, -52.89915, 
        -52.8071, -52.72481, -52.65497, -52.597, -52.54961, -52.5106, 
        -52.47681, -52.44619, -52.41735, -52.3895, -52.36268, -52.33779, 
        -52.31571, -52.29733, -52.28293, -52.27352, -52.26955, -52.26995, 
        -52.27668, -52.28839, -52.30421, -52.32425, -52.34868, -52.37741, 
        -52.41054, -52.44764, -52.48776, -52.52953, -52.57138, -52.61164, 
        -52.64867, -52.68179, -52.7103, -52.73375, -52.75217, -52.76506, 
        -52.7724, -52.77293, -52.76551, -52.75121, -52.72852, -52.69752, 
        -52.65837, -52.61211, -52.5595, -52.50158, -52.43959, -52.37429, 
        -52.30615, -52.23533, -52.16214, -52.08714, -52.01038, -51.93223, 
        -51.85302, -51.773, -51.69266, -51.61276, -51.53412, -51.45714, 
        -51.38168, -51.31068, -51.24344, -51.18062, -51.12168, -51.06668, 
        -51.01585, -50.96841, -50.92492, -50.88429, -50.8464, -50.81128, 
        -50.77842, -50.7478, -50.71882, -50.69073, -50.66338, -50.63666, 
        -50.61068, -50.58553, -50.56126, -50.53806, -50.51672, -50.49704, 
        -50.47877, -50.45992, -50.44151, -50.42169, -50.4, -50.37553, 
        -50.34803, -50.31774, -50.28486, -50.24949, -50.21194, -50.1721, 
        -50.13097, -50.08891, -50.04689, -50.00496, -49.96268, -49.92031, 
        -49.87714, -49.83368, -49.78934, -49.74415, -49.69822, -49.65101, 
        -49.60277, -49.55327, -49.50253, -49.45099, -49.3987, -49.34595, 
        -49.2913, -49.23693, -49.18128, -49.12424, -49.06533, -49.00328, 
        -48.93778, -48.86876, -48.79602, -48.7203, -48.64196, -48.56198, 
        -48.48129, -48.40071, -48.32071, -48.24162, -48.16399, -48.08797, 
        -48.01202, -47.93604, -47.85999, -47.7834, -47.70657, -47.6296, 
        -47.55275, -47.47573, -47.39814, -47.32008, -47.24123, -47.16069, 
        -47.07778, -46.99157, -46.90268, -46.81013, -46.71793, -46.62741, 
        -46.54114, -46.46172, -46.39267, -46.33546, -46.29169, -46.26186, 
        -46.24557, -46.24173, -46.24976, -46.26797, -46.2949, -46.32942, 
        -46.37005, -46.41513, -46.46272, -46.51082, -46.55751, -46.60114, 
        -46.64091, -46.67593, -46.70662, -46.73373, -46.75879, -46.78282, 
        -46.80845, -46.83813, -46.87445, -46.91972, -46.97519, -47.04112, 
        -47.11612, -47.1982, -47.28466, -47.37235, -47.45872, -47.54257, 
        -47.62308, -47.70089, -47.77783, -47.85445, -47.93544, -48.0209, 
        -48.11382, -48.21552, -48.32674, -48.44806, -48.57984, -48.72256, 
        -48.87762,
  -38.8133, -38.92376, -39.03049, -39.16049, -39.28353, -39.39667, 
        -39.49973, -39.59168, -39.67924, -39.78307, -39.88914, -39.99089, 
        -40.09372, -40.21249, -40.32018, -40.42899, -40.56097, -40.70543, 
        -40.85894, -41.00354, -41.15708, -41.31532, -41.47084, -41.62601, 
        -41.78148, -41.93208, -42.07903, -42.22835, -42.37751, -42.52813, 
        -42.68055, -42.8308, -42.98058, -43.12931, -43.27714, -43.42324, 
        -43.56596, -43.70607, -43.84315, -43.97753, -44.10961, -44.23829, 
        -44.36523, -44.48952, -44.61109, -44.72956, -44.84507, -44.95871, 
        -45.07157, -45.18365, -45.29548, -45.40689, -45.51805, -45.62818, 
        -45.73754, -45.84621, -45.95473, -46.06439, -46.17534, -46.2906, 
        -46.40934, -46.53249, -46.65923, -46.7891, -46.92243, -47.0593, 
        -47.1997, -47.344, -47.49253, -47.64487, -47.80148, -47.96279, 
        -48.12867, -48.29914, -48.47388, -48.65212, -48.83669, -49.02775, 
        -49.22789, -49.43822, -49.66105, -49.89785, -50.15038, -50.41737, 
        -50.69668, -50.98467, -51.2755, -51.56225, -51.83752, -52.09288, 
        -52.32137, -52.5166, -52.67398, -52.78848, -52.86057, -52.88877, 
        -52.87572, -52.82674, -52.74868, -52.65113, -52.54385, -52.43645, 
        -52.33605, -52.2481, -52.17436, -52.11383, -52.06527, -52.02544, 
        -51.99173, -51.96085, -51.93191, -51.90393, -51.87621, -51.85133, 
        -51.82987, -51.81264, -51.79977, -51.79217, -51.79031, -51.79371, 
        -51.80203, -51.81435, -51.83018, -51.84931, -51.87177, -51.89776, 
        -51.9273, -51.95999, -51.99508, -52.03145, -52.06768, -52.10214, 
        -52.13253, -52.16017, -52.18368, -52.20249, -52.21657, -52.22577, 
        -52.22989, -52.228, -52.21963, -52.20406, -52.18119, -52.15072, 
        -52.11332, -52.06966, -52.02014, -51.96514, -51.90683, -51.84512, 
        -51.78057, -51.71394, -51.64522, -51.57528, -51.50297, -51.43069, 
        -51.35744, -51.28293, -51.20787, -51.13229, -51.05719, -50.98282, 
        -50.91009, -50.84024, -50.77389, -50.71183, -50.65367, -50.5995, 
        -50.54921, -50.50221, -50.45873, -50.41814, -50.3801, -50.34451, 
        -50.31117, -50.28022, -50.25084, -50.22223, -50.19322, -50.16582, 
        -50.13941, -50.11411, -50.09001, -50.0675, -50.04683, -50.0282, 
        -50.01138, -49.99542, -49.97936, -49.96226, -49.94335, -49.92179, 
        -49.89728, -49.87003, -49.84011, -49.80804, -49.77375, -49.73767, 
        -49.70041, -49.66257, -49.62472, -49.58679, -49.5483, -49.5093, 
        -49.46943, -49.42795, -49.38662, -49.34395, -49.30043, -49.25584, 
        -49.21003, -49.16297, -49.11472, -49.06548, -49.01529, -48.96476, 
        -48.91318, -48.86074, -48.80705, -48.75164, -48.69412, -48.63392, 
        -48.57042, -48.50367, -48.43341, -48.36095, -48.28646, -48.2108, 
        -48.13478, -48.05907, -47.98396, -47.90931, -47.83541, -47.76263, 
        -47.68977, -47.61644, -47.54258, -47.46675, -47.39125, -47.31506, 
        -47.23843, -47.16135, -47.08302, -47.0032, -46.92144, -46.83677, 
        -46.74848, -46.65658, -46.56173, -46.46548, -46.3704, -46.27913, 
        -46.1948, -46.11984, -46.05634, -46.00645, -45.97079, -45.94881, 
        -45.93933, -45.94114, -45.95312, -45.97335, -46.00049, -46.0338, 
        -46.0718, -46.11331, -46.15677, -46.20035, -46.24263, -46.28186, 
        -46.31727, -46.3486, -46.37649, -46.40127, -46.42455, -46.44675, 
        -46.47217, -46.50205, -46.5389, -46.58468, -46.64052, -46.70678, 
        -46.78236, -46.86509, -46.95258, -47.0421, -47.131, -47.21799, 
        -47.3026, -47.38649, -47.4701, -47.55519, -47.64476, -47.7407, 
        -47.84495, -47.95903, -48.08356, -48.21924, -48.36614, -48.52422, 
        -48.69362,
  -38.71203, -38.81794, -38.92833, -39.04499, -39.16694, -39.27493, 
        -39.3638, -39.4641, -39.55927, -39.65489, -39.75311, -39.84611, 
        -39.94981, -40.05188, -40.15287, -40.25285, -40.3745, -40.51509, 
        -40.64781, -40.77402, -40.93658, -41.0942, -41.24836, -41.40341, 
        -41.55627, -41.7033, -41.84921, -41.99547, -42.14301, -42.29071, 
        -42.4391, -42.58768, -42.73489, -42.88272, -43.0295, -43.17462, 
        -43.31575, -43.45503, -43.59122, -43.72441, -43.85572, -43.98412, 
        -44.10929, -44.23161, -44.35062, -44.46629, -44.579, -44.68998, 
        -44.80044, -44.9104, -45.02032, -45.13054, -45.23952, -45.34864, 
        -45.45632, -45.56304, -45.66912, -45.77582, -45.88415, -45.99543, 
        -46.11014, -46.22861, -46.35099, -46.47711, -46.60722, -46.74145, 
        -46.87991, -47.02291, -47.17016, -47.32043, -47.47597, -47.63635, 
        -47.80135, -47.97125, -48.14542, -48.32384, -48.50797, -48.69907, 
        -48.89884, -49.10863, -49.33111, -49.56767, -49.81908, -50.08474, 
        -50.36287, -50.64966, -50.93853, -51.22401, -51.49759, -51.75071, 
        -51.97579, -52.16602, -52.31654, -52.42331, -52.48469, -52.50072, 
        -52.47387, -52.40984, -52.31714, -52.20577, -52.08632, -51.96885, 
        -51.86089, -51.76726, -51.68967, -51.62616, -51.57629, -51.5363, 
        -51.50238, -51.47145, -51.44225, -51.41482, -51.38832, -51.36411, 
        -51.34337, -51.32747, -51.31692, -51.31202, -51.31293, -51.31891, 
        -51.32927, -51.34294, -51.3592, -51.37767, -51.39842, -51.42039, 
        -51.44613, -51.47456, -51.50483, -51.5361, -51.56692, -51.59608, 
        -51.6225, -51.6453, -51.66396, -51.67846, -51.68876, -51.69485, 
        -51.69608, -51.69201, -51.68202, -51.66594, -51.64333, -51.61419, 
        -51.57858, -51.53724, -51.49002, -51.43905, -51.38433, -51.32591, 
        -51.2649, -51.20198, -51.13771, -51.07243, -51.00584, -50.93833, 
        -50.87, -50.80045, -50.72974, -50.65794, -50.58569, -50.51368, 
        -50.44286, -50.37427, -50.30883, -50.24706, -50.18968, -50.13621, 
        -50.08649, -50.04005, -49.99577, -49.95531, -49.91739, -49.88187, 
        -49.84849, -49.8173, -49.78796, -49.7593, -49.73158, -49.70384, 
        -49.67749, -49.65254, -49.62883, -49.60693, -49.58706, -49.56937, 
        -49.55354, -49.53895, -49.52463, -49.50938, -49.49277, -49.47369, 
        -49.45185, -49.42757, -49.40073, -49.37086, -49.34022, -49.30825, 
        -49.27562, -49.24258, -49.20952, -49.17648, -49.14272, -49.10799, 
        -49.07191, -49.03471, -48.99621, -48.95608, -48.91459, -48.87175, 
        -48.82756, -48.78223, -48.73563, -48.68797, -48.6393, -48.59025, 
        -48.54054, -48.48971, -48.4379, -48.38407, -48.32841, -48.27018, 
        -48.20921, -48.14518, -48.0784, -48.00863, -47.93856, -47.86762, 
        -47.79663, -47.72611, -47.6562, -47.58643, -47.51677, -47.44753, 
        -47.37769, -47.30676, -47.23494, -47.16197, -47.08787, -47.01252, 
        -46.93628, -46.85921, -46.78053, -46.69935, -46.61488, -46.52675, 
        -46.43427, -46.33799, -46.23891, -46.13966, -46.04288, -45.95243, 
        -45.87094, -45.80076, -45.7443, -45.70208, -45.67429, -45.65968, 
        -45.65646, -45.66323, -45.67713, -45.69875, -45.72564, -45.75708, 
        -45.79223, -45.83028, -45.86968, -45.90905, -45.94695, -45.98194, 
        -46.01334, -46.04117, -46.06629, -46.08928, -46.11191, -46.13514, 
        -46.16076, -46.1921, -46.23037, -46.27694, -46.33259, -46.39846, 
        -46.47381, -46.5559, -46.64265, -46.73198, -46.82178, -46.911, 
        -46.99936, -47.08843, -47.17851, -47.27257, -47.37143, -47.4784, 
        -47.59451, -47.72144, -47.86, -48.01053, -48.17255, -48.34538, 
        -48.52783,
  -38.61626, -38.71495, -38.82953, -38.93879, -39.05788, -39.15897, 
        -39.23862, -39.34171, -39.4421, -39.53725, -39.63046, -39.71556, 
        -39.81263, -39.90564, -39.99638, -40.09785, -40.21571, -40.33036, 
        -40.46976, -40.60082, -40.73904, -40.89817, -41.05042, -41.20055, 
        -41.34574, -41.48894, -41.63421, -41.77945, -41.92456, -42.06977, 
        -42.21399, -42.35935, -42.50511, -42.65121, -42.79739, -42.94202, 
        -43.08365, -43.22224, -43.35786, -43.49057, -43.62092, -43.74813, 
        -43.87204, -43.99237, -44.109, -44.22206, -44.3317, -44.44028, 
        -44.54823, -44.65599, -44.76411, -44.87262, -44.98085, -45.08828, 
        -45.19408, -45.29856, -45.40187, -45.50519, -45.60978, -45.71648, 
        -45.82659, -45.94042, -46.05821, -46.17957, -46.30663, -46.43867, 
        -46.57585, -46.71801, -46.86466, -47.01521, -47.17002, -47.32926, 
        -47.49312, -47.66193, -47.83497, -48.01291, -48.19663, -48.38711, 
        -48.58588, -48.79474, -49.01457, -49.24891, -49.49754, -49.75999, 
        -50.03479, -50.31832, -50.60485, -50.88702, -51.15674, -51.40556, 
        -51.62542, -51.80917, -51.95182, -52.04953, -52.1, -52.1038, 
        -52.06354, -51.98569, -51.87806, -51.75375, -51.62323, -51.49633, 
        -51.3812, -51.28252, -51.20137, -51.13618, -51.08544, -51.04486, 
        -51.0103, -50.97911, -50.9496, -50.92241, -50.89649, -50.87263, 
        -50.85314, -50.83897, -50.83112, -50.82928, -50.83252, -50.84176, 
        -50.85483, -50.87053, -50.88781, -50.90613, -50.92553, -50.94638, 
        -50.96891, -50.9933, -51.01924, -51.04562, -51.07165, -51.09607, 
        -51.11776, -51.13618, -51.15068, -51.16112, -51.1685, -51.17165, 
        -51.17052, -51.16375, -51.15266, -51.1366, -51.11445, -51.08637, 
        -51.05264, -51.01366, -50.97067, -50.92323, -50.87171, -50.81685, 
        -50.75911, -50.70029, -50.6399, -50.57833, -50.51596, -50.4526, 
        -50.38867, -50.32307, -50.2556, -50.18718, -50.11753, -50.04714, 
        -49.978, -49.91068, -49.84599, -49.78509, -49.72857, -49.67601, 
        -49.62666, -49.58085, -49.5379, -49.49792, -49.46027, -49.42475, 
        -49.3918, -49.36092, -49.33224, -49.30438, -49.27692, -49.25008, 
        -49.22425, -49.20005, -49.17671, -49.15555, -49.1366, -49.11992, 
        -49.10368, -49.09009, -49.077, -49.06316, -49.04791, -49.03085, 
        -49.01148, -48.9895, -48.96564, -48.93994, -48.91319, -48.88546, 
        -48.8573, -48.8291, -48.80109, -48.77334, -48.74473, -48.71449, 
        -48.68262, -48.6487, -48.6132, -48.57543, -48.53565, -48.49427, 
        -48.45137, -48.40724, -48.36193, -48.31553, -48.26732, -48.21954, 
        -48.17156, -48.12257, -48.07259, -48.02092, -47.9673, -47.91168, 
        -47.8537, -47.79309, -47.73032, -47.66579, -47.60069, -47.53502, 
        -47.46944, -47.4043, -47.33966, -47.27514, -47.20985, -47.14386, 
        -47.07693, -47.00845, -46.9385, -46.867, -46.79409, -46.71984, 
        -46.64429, -46.56759, -46.48906, -46.40679, -46.32074, -46.23008, 
        -46.13491, -46.03447, -45.93318, -45.83248, -45.736, -45.64742, 
        -45.56961, -45.50493, -45.45522, -45.42017, -45.39932, -45.39084, 
        -45.39277, -45.40301, -45.41993, -45.44199, -45.46823, -45.49747, 
        -45.52947, -45.56395, -45.59951, -45.63488, -45.66872, -45.69991, 
        -45.72794, -45.75318, -45.77644, -45.79902, -45.82177, -45.84639, 
        -45.87503, -45.9097, -45.95066, -45.99831, -46.05344, -46.11745, 
        -46.19002, -46.26962, -46.35381, -46.44124, -46.53075, -46.62114, 
        -46.71281, -46.80561, -46.90283, -47.00518, -47.11438, -47.2324, 
        -47.36106, -47.50162, -47.65463, -47.81997, -47.9964, -48.18233, 
        -48.37537,
  -38.52822, -38.62646, -38.73544, -38.85345, -38.95995, -39.05472, 
        -39.13063, -39.22042, -39.32724, -39.42305, -39.51237, -39.59806, 
        -39.6846, -39.76577, -39.86374, -39.95676, -40.06882, -40.17939, 
        -40.3037, -40.43836, -40.57072, -40.71954, -40.86456, -41.00678, 
        -41.15003, -41.2884, -41.42965, -41.57411, -41.71785, -41.86173, 
        -42.00465, -42.14854, -42.29231, -42.43739, -42.58278, -42.72682, 
        -42.86811, -43.00615, -43.14093, -43.27325, -43.40266, -43.52796, 
        -43.65068, -43.76946, -43.88408, -43.99522, -44.10361, -44.21025, 
        -44.31612, -44.42152, -44.52765, -44.63379, -44.73974, -44.84465, 
        -44.94812, -45.04983, -45.15025, -45.24927, -45.35007, -45.45271, 
        -45.55804, -45.66681, -45.77995, -45.89809, -46.022, -46.15221, 
        -46.28918, -46.43087, -46.57771, -46.72833, -46.88258, -47.04032, 
        -47.20264, -47.36975, -47.54052, -47.71772, -47.90071, -48.09034, 
        -48.28778, -48.49452, -48.71236, -48.94301, -49.18726, -49.44488, 
        -49.71454, -49.99298, -50.27415, -50.55067, -50.81443, -51.05675, 
        -51.26947, -51.44556, -51.57863, -51.66662, -51.70628, -51.69834, 
        -51.64533, -51.5546, -51.43582, -51.29997, -51.15911, -51.02368, 
        -50.90222, -50.79863, -50.71352, -50.6462, -50.59338, -50.55111, 
        -50.51515, -50.48286, -50.45285, -50.42374, -50.39772, -50.37453, 
        -50.35601, -50.34374, -50.33837, -50.34022, -50.34855, -50.36163, 
        -50.37818, -50.3965, -50.41556, -50.43467, -50.45374, -50.47308, 
        -50.49319, -50.51457, -50.53676, -50.55906, -50.58066, -50.59979, 
        -50.61731, -50.63124, -50.64199, -50.64923, -50.65332, -50.6543, 
        -50.65129, -50.64434, -50.63279, -50.61649, -50.59501, -50.56855, 
        -50.53662, -50.49998, -50.45943, -50.4149, -50.36652, -50.31495, 
        -50.26054, -50.20464, -50.14766, -50.08894, -50.03011, -49.97039, 
        -49.90949, -49.84708, -49.78291, -49.71699, -49.64998, -49.58276, 
        -49.516, -49.45029, -49.3871, -49.32737, -49.27163, -49.21986, 
        -49.1713, -49.12595, -49.08355, -49.04375, -49.00643, -48.97178, 
        -48.93957, -48.90974, -48.88197, -48.85445, -48.82876, -48.80358, 
        -48.7792, -48.75585, -48.73379, -48.71417, -48.69633, -48.67984, 
        -48.66563, -48.65287, -48.64027, -48.6272, -48.61306, -48.59705, 
        -48.57937, -48.55951, -48.53809, -48.51521, -48.49154, -48.46763, 
        -48.4439, -48.42044, -48.39733, -48.37426, -48.35053, -48.32506, 
        -48.29627, -48.26574, -48.23261, -48.19685, -48.15868, -48.11852, 
        -48.07684, -48.03387, -47.98969, -47.94482, -47.8992, -47.85329, 
        -47.80721, -47.76055, -47.71293, -47.66393, -47.61307, -47.56049, 
        -47.50597, -47.4495, -47.3912, -47.3317, -47.27166, -47.21146, 
        -47.15147, -47.09182, -47.03259, -46.97307, -46.91207, -46.84962, 
        -46.78555, -46.71851, -46.65015, -46.58012, -46.50813, -46.43502, 
        -46.36058, -46.28455, -46.20639, -46.12436, -46.03756, -45.9459, 
        -45.84897, -45.7482, -45.64624, -45.54591, -45.45123, -45.3658, 
        -45.29242, -45.23336, -45.18954, -45.1605, -45.1451, -45.14112, 
        -45.14643, -45.1586, -45.17607, -45.19766, -45.22249, -45.24942, 
        -45.27867, -45.3096, -45.34155, -45.3735, -45.40418, -45.4324, 
        -45.45793, -45.48119, -45.5041, -45.52609, -45.55065, -45.57807, 
        -45.61068, -45.64928, -45.69305, -45.74203, -45.79712, -45.85919, 
        -45.92856, -46.00373, -46.08416, -46.16873, -46.25686, -46.34788, 
        -46.44241, -46.54142, -46.64602, -46.75747, -46.87702, -47.00657, 
        -47.14791, -47.30201, -47.46904, -47.64798, -47.83716, -48.0334, 
        -48.23489,
  -38.4497, -38.5491, -38.65839, -38.76868, -38.86969, -38.95615, 
        -39.04072, -39.11885, -39.2136, -39.30618, -39.39793, -39.4851, 
        -39.56812, -39.6478, -39.73441, -39.83536, -39.93689, -40.04256, 
        -40.16063, -40.28119, -40.40665, -40.54643, -40.68659, -40.82551, 
        -40.96544, -41.10328, -41.2413, -41.38144, -41.52549, -41.67061, 
        -41.81387, -41.95564, -42.09871, -42.2416, -42.3856, -42.5276, 
        -42.66877, -42.80542, -42.93993, -43.07125, -43.19968, -43.32475, 
        -43.4461, -43.56307, -43.67591, -43.78529, -43.89224, -43.9969, 
        -44.1009, -44.20465, -44.30851, -44.41144, -44.51468, -44.61665, 
        -44.71715, -44.81606, -44.91322, -45.00947, -45.10622, -45.20427, 
        -45.30481, -45.40885, -45.51783, -45.63288, -45.75428, -45.88366, 
        -46.0198, -46.1618, -46.30832, -46.45908, -46.61251, -46.76884, 
        -46.92916, -47.0939, -47.26392, -47.43943, -47.62091, -47.80874, 
        -48.00391, -48.20773, -48.42179, -48.64756, -48.88626, -49.13794, 
        -49.40094, -49.67111, -49.94481, -50.21349, -50.46914, -50.70315, 
        -50.90726, -51.07461, -51.19959, -51.27802, -51.30756, -51.28859, 
        -51.22457, -51.12305, -50.99347, -50.8478, -50.69782, -50.55463, 
        -50.42709, -50.31813, -50.22792, -50.15704, -50.10104, -50.0561, 
        -50.0181, -49.98389, -49.95212, -49.92263, -49.89571, -49.87251, 
        -49.85494, -49.8442, -49.84149, -49.84664, -49.85907, -49.8764, 
        -49.8968, -49.91879, -49.94031, -49.96123, -49.98025, -49.99932, 
        -50.01807, -50.0371, -50.05634, -50.07532, -50.09334, -50.10964, 
        -50.12336, -50.1339, -50.14174, -50.14645, -50.14794, -50.14683, 
        -50.14231, -50.13442, -50.12239, -50.1057, -50.08405, -50.05813, 
        -50.02752, -49.99127, -49.95254, -49.91014, -49.86462, -49.81574, 
        -49.76461, -49.71164, -49.65755, -49.60326, -49.54792, -49.49135, 
        -49.43349, -49.37391, -49.31242, -49.24937, -49.18494, -49.12012, 
        -49.05544, -48.99226, -48.9312, -48.87311, -48.81865, -48.7678, 
        -48.71896, -48.67459, -48.63266, -48.59335, -48.55668, -48.52244, 
        -48.49125, -48.46263, -48.43636, -48.41174, -48.38795, -48.36516, 
        -48.34286, -48.32155, -48.30167, -48.28391, -48.26741, -48.25238, 
        -48.23871, -48.22622, -48.2139, -48.20131, -48.18778, -48.17282, 
        -48.15607, -48.13789, -48.11736, -48.09677, -48.07586, -48.05511, 
        -48.03497, -48.01553, -47.99649, -47.97749, -47.95777, -47.93614, 
        -47.91203, -47.88429, -47.85347, -47.81946, -47.78294, -47.74421, 
        -47.70376, -47.66198, -47.61922, -47.57611, -47.53276, -47.48939, 
        -47.44598, -47.40223, -47.35757, -47.31186, -47.2644, -47.21538, 
        -47.16476, -47.11161, -47.05836, -47.00425, -46.94968, -46.89503, 
        -46.84076, -46.78679, -46.7326, -46.67778, -46.62078, -46.56169, 
        -46.50014, -46.43614, -46.36967, -46.30082, -46.23051, -46.15877, 
        -46.08571, -46.01076, -45.93363, -45.85278, -45.76664, -45.67507, 
        -45.57835, -45.47817, -45.37706, -45.27903, -45.18736, -45.10598, 
        -45.0375, -44.98358, -44.94458, -44.92027, -44.90843, -44.90739, 
        -44.91316, -44.92525, -44.94211, -44.96252, -44.985, -45.00945, 
        -45.03581, -45.0637, -45.09251, -45.12104, -45.14875, -45.17465, 
        -45.19878, -45.22164, -45.24487, -45.26963, -45.29723, -45.32853, 
        -45.36526, -45.40733, -45.45369, -45.50425, -45.55949, -45.6199, 
        -45.68604, -45.75729, -45.83344, -45.91474, -46.00129, -46.09338, 
        -46.19036, -46.29512, -46.4078, -46.52868, -46.65844, -46.80033, 
        -46.95433, -47.12099, -47.30022, -47.49038, -47.68876, -47.89238, 
        -48.09725,
  -38.38452, -38.4837, -38.58629, -38.68767, -38.78387, -38.87305, 
        -38.95869, -39.04109, -39.12638, -39.2058, -39.29171, -39.37989, 
        -39.46236, -39.54032, -39.62303, -39.71764, -39.81532, -39.9206, 
        -40.02978, -40.14297, -40.2636, -40.39362, -40.52694, -40.66099, 
        -40.79518, -40.93072, -41.06751, -41.20638, -41.3475, -41.49374, 
        -41.63737, -41.7794, -41.92192, -42.06389, -42.20535, -42.34682, 
        -42.48698, -42.62284, -42.75566, -42.88586, -43.01346, -43.13703, 
        -43.25674, -43.37209, -43.48315, -43.59104, -43.69534, -43.79881, 
        -43.90132, -44.003, -44.10493, -44.20625, -44.30653, -44.40566, 
        -44.5029, -44.59813, -44.69194, -44.78467, -44.87723, -44.97076, 
        -45.06671, -45.16648, -45.27079, -45.38301, -45.50294, -45.6311, 
        -45.76717, -45.91013, -46.05767, -46.20831, -46.36074, -46.51505, 
        -46.6727, -46.83469, -47.00182, -47.17477, -47.35394, -47.53931, 
        -47.73159, -47.93059, -48.14008, -48.36009, -48.59225, -48.83659, 
        -49.09194, -49.35457, -49.61893, -49.87801, -50.12365, -50.3476, 
        -50.54194, -50.70006, -50.81597, -50.88529, -50.90573, -50.87747, 
        -50.80445, -50.69311, -50.55504, -50.40133, -50.24393, -50.09438, 
        -49.9607, -49.84598, -49.75156, -49.67593, -49.6152, -49.56577, 
        -49.52371, -49.48598, -49.45128, -49.4193, -49.39054, -49.36648, 
        -49.34925, -49.34007, -49.33961, -49.34707, -49.36284, -49.38434, 
        -49.40941, -49.43509, -49.46017, -49.48368, -49.50542, -49.52554, 
        -49.5438, -49.5615, -49.57864, -49.59504, -49.61018, -49.62332, 
        -49.63374, -49.6416, -49.64645, -49.64888, -49.64871, -49.64557, 
        -49.63894, -49.62971, -49.61705, -49.59971, -49.57799, -49.55191, 
        -49.52179, -49.48777, -49.44985, -49.40915, -49.36558, -49.3194, 
        -49.27117, -49.22097, -49.16975, -49.11802, -49.06563, -49.01231, 
        -48.95732, -48.90055, -48.84192, -48.78159, -48.71925, -48.65717, 
        -48.59541, -48.53506, -48.47659, -48.42086, -48.36816, -48.3185, 
        -48.27168, -48.22828, -48.18703, -48.14853, -48.11239, -48.07915, 
        -48.04898, -48.02188, -47.99742, -47.97518, -47.95421, -47.93431, 
        -47.91504, -47.89672, -47.87958, -47.86394, -47.84968, -47.83537, 
        -47.8228, -47.81054, -47.7984, -47.78598, -47.7727, -47.75822, 
        -47.74237, -47.72512, -47.70692, -47.68813, -47.6691, -47.65067, 
        -47.63331, -47.61677, -47.60085, -47.5848, -47.56809, -47.54924, 
        -47.5277, -47.50266, -47.47377, -47.44143, -47.4062, -47.36882, 
        -47.32981, -47.2896, -47.24877, -47.20697, -47.16647, -47.12635, 
        -47.08627, -47.04619, -47.00518, -46.96333, -46.92006, -46.87498, 
        -46.82864, -46.78106, -46.7328, -46.68413, -46.63516, -46.58631, 
        -46.53777, -46.48912, -46.44001, -46.38955, -46.33656, -46.28028, 
        -46.22112, -46.15934, -46.09457, -46.02752, -45.95889, -45.88877, 
        -45.81751, -45.74468, -45.66906, -45.5901, -45.50545, -45.41453, 
        -45.3198, -45.22168, -45.12344, -45.029, -44.9418, -44.86518, 
        -44.80183, -44.7525, -44.71754, -44.69612, -44.68623, -44.68585, 
        -44.69237, -44.70329, -44.71817, -44.73609, -44.75603, -44.77795, 
        -44.80139, -44.82635, -44.85218, -44.87804, -44.90348, -44.92786, 
        -44.95131, -44.97466, -44.99944, -45.0266, -45.05775, -45.09354, 
        -45.1336, -45.1787, -45.22764, -45.28031, -45.33593, -45.39475, 
        -45.4576, -45.52538, -45.59819, -45.67676, -45.76323, -45.85563, 
        -45.95725, -46.0681, -46.18856, -46.31955, -46.46127, -46.61456, 
        -46.77982, -46.9572, -47.14615, -47.34406, -47.54783, -47.75363, 
        -47.95814,
  -38.32653, -38.4231, -38.51878, -38.61415, -38.70675, -38.79591, 
        -38.87962, -38.96026, -39.04034, -39.12064, -39.19762, -39.28126, 
        -39.36285, -39.43953, -39.51806, -39.60943, -39.70779, -39.80651, 
        -39.91085, -40.01893, -40.13514, -40.25732, -40.38358, -40.51217, 
        -40.6426, -40.77269, -40.90892, -41.04661, -41.18575, -41.32935, 
        -41.47568, -41.61869, -41.76199, -41.90418, -42.04466, -42.18287, 
        -42.32184, -42.45672, -42.5881, -42.71694, -42.8418, -42.96383, 
        -43.08172, -43.19508, -43.3046, -43.41075, -43.51469, -43.6171, 
        -43.71791, -43.8179, -43.91758, -44.01615, -44.1135, -44.20948, 
        -44.30355, -44.39564, -44.48484, -44.57381, -44.6624, -44.75174, 
        -44.84338, -44.93942, -45.04171, -45.15151, -45.27032, -45.39792, 
        -45.53408, -45.67673, -45.82415, -45.97401, -46.1249, -46.27687, 
        -46.4312, -46.58866, -46.7524, -46.92219, -47.09803, -47.27951, 
        -47.46788, -47.66315, -47.86674, -48.08055, -48.30564, -48.54219, 
        -48.78851, -49.04129, -49.29466, -49.54223, -49.77635, -49.98915, 
        -50.17339, -50.32088, -50.42843, -50.49003, -50.503, -50.46775, 
        -50.38861, -50.27272, -50.12883, -49.96967, -49.80725, -49.6524, 
        -49.5124, -49.3907, -49.28969, -49.20713, -49.13957, -49.0837, 
        -49.0357, -48.99229, -48.95194, -48.9163, -48.88465, -48.85871, 
        -48.84088, -48.83236, -48.83391, -48.84469, -48.86351, -48.88859, 
        -48.9174, -48.94778, -48.97686, -49.00342, -49.0279, -49.04978, 
        -49.06873, -49.08599, -49.10187, -49.11565, -49.12728, -49.13799, 
        -49.14587, -49.15115, -49.15377, -49.15416, -49.15246, -49.14802, 
        -49.14087, -49.13055, -49.11654, -49.09843, -49.07613, -49.0493, 
        -49.01897, -48.98516, -48.94835, -48.90837, -48.86658, -48.82246, 
        -48.77676, -48.72961, -48.68021, -48.63111, -48.5815, -48.53112, 
        -48.47933, -48.42546, -48.3698, -48.31257, -48.25447, -48.19616, 
        -48.13809, -48.081, -48.0256, -47.97256, -47.92216, -47.87396, 
        -47.82895, -47.78612, -47.74622, -47.70823, -47.67314, -47.64046, 
        -47.61147, -47.58616, -47.56315, -47.54382, -47.52614, -47.50952, 
        -47.4942, -47.47964, -47.46597, -47.45345, -47.44141, -47.43015, 
        -47.41908, -47.40751, -47.39576, -47.38327, -47.36994, -47.35595, 
        -47.34038, -47.32368, -47.30614, -47.28841, -47.27101, -47.25423, 
        -47.23862, -47.22407, -47.20998, -47.19581, -47.18086, -47.16299, 
        -47.14314, -47.11975, -47.09277, -47.06185, -47.02794, -46.99187, 
        -46.95443, -46.91621, -46.87772, -46.83944, -46.80231, -46.76606, 
        -46.73019, -46.69442, -46.65801, -46.62038, -46.58168, -46.54128, 
        -46.49947, -46.45632, -46.41294, -46.36936, -46.32611, -46.28302, 
        -46.23992, -46.19655, -46.15205, -46.10579, -46.05638, -46.00211, 
        -45.94542, -45.88582, -45.82331, -45.75819, -45.69159, -45.62364, 
        -45.55433, -45.48406, -45.41097, -45.33421, -45.25233, -45.16504, 
        -45.07365, -44.9794, -44.88546, -44.79589, -44.71414, -44.64294, 
        -44.58462, -44.53971, -44.50771, -44.48801, -44.47823, -44.47684, 
        -44.48122, -44.48972, -44.50156, -44.51643, -44.5337, -44.55299, 
        -44.57395, -44.59658, -44.61981, -44.6437, -44.66729, -44.69068, 
        -44.71426, -44.73789, -44.76472, -44.79493, -44.82906, -44.86864, 
        -44.91302, -44.96065, -45.01196, -45.06573, -45.12161, -45.17899, 
        -45.23907, -45.3044, -45.37559, -45.45403, -45.54131, -45.63832, 
        -45.74507, -45.8643, -45.9931, -46.13479, -46.28818, -46.4534, 
        -46.62815, -46.81371, -47.00804, -47.20879, -47.41246, -47.61553, 
        -47.81445,
  -38.26963, -38.36381, -38.45409, -38.54482, -38.63369, -38.71923, 
        -38.80142, -38.87984, -38.9574, -39.03602, -39.11235, -39.19102, 
        -39.2724, -39.34907, -39.42633, -39.51068, -39.60594, -39.70243, 
        -39.80354, -39.90541, -40.01822, -40.13536, -40.25583, -40.37896, 
        -40.50388, -40.63293, -40.76658, -40.90361, -41.0423, -41.18321, 
        -41.32628, -41.47239, -41.61668, -41.75917, -41.89863, -42.03456, 
        -42.1712, -42.30523, -42.43474, -42.56167, -42.68587, -42.80615, 
        -42.92255, -43.03409, -43.1418, -43.24634, -43.34854, -43.44928, 
        -43.54855, -43.64705, -43.74481, -43.83997, -43.9347, -44.02781, 
        -44.11864, -44.20776, -44.2948, -44.37998, -44.46454, -44.54984, 
        -44.63768, -44.73067, -44.83067, -44.93921, -45.05687, -45.18381, 
        -45.31924, -45.46007, -45.60601, -45.75392, -45.90236, -46.05158, 
        -46.2024, -46.35715, -46.51678, -46.68217, -46.85363, -47.03079, 
        -47.2139, -47.40367, -47.60149, -47.80838, -48.02557, -48.25299, 
        -48.4891, -48.72928, -48.97033, -49.20513, -49.42674, -49.62774, 
        -49.80134, -49.94145, -50.04116, -50.09682, -50.10517, -50.06657, 
        -49.98497, -49.86679, -49.72131, -49.55969, -49.39372, -49.23418, 
        -49.08815, -48.95824, -48.84789, -48.75609, -48.67924, -48.61376, 
        -48.55784, -48.50658, -48.46089, -48.41983, -48.38421, -48.35519, 
        -48.33551, -48.32658, -48.32855, -48.34086, -48.36225, -48.39028, 
        -48.4227, -48.45686, -48.49006, -48.51972, -48.54662, -48.57027, 
        -48.59108, -48.60831, -48.62322, -48.63622, -48.6465, -48.65478, 
        -48.6606, -48.66427, -48.665, -48.66372, -48.66063, -48.65519, 
        -48.64681, -48.6352, -48.61982, -48.60065, -48.57742, -48.54942, 
        -48.51732, -48.48305, -48.44622, -48.4074, -48.36688, -48.32454, 
        -48.28101, -48.23666, -48.19142, -48.14516, -48.09827, -48.0508, 
        -48.00207, -47.95173, -47.89926, -47.84568, -47.79115, -47.7368, 
        -47.68283, -47.62973, -47.57792, -47.52798, -47.48014, -47.43308, 
        -47.38965, -47.34843, -47.30932, -47.27231, -47.2378, -47.20632, 
        -47.1785, -47.15499, -47.135, -47.11879, -47.10468, -47.09206, 
        -47.08073, -47.07056, -47.06086, -47.05188, -47.04269, -47.03411, 
        -47.0246, -47.01429, -47.00266, -46.99055, -46.97715, -46.96299, 
        -46.94737, -46.93014, -46.91319, -46.89622, -46.87968, -46.86407, 
        -46.84953, -46.83612, -46.8229, -46.80955, -46.7952, -46.77929, 
        -46.76042, -46.73825, -46.7126, -46.68332, -46.651, -46.61651, 
        -46.58076, -46.54453, -46.5087, -46.47377, -46.44005, -46.40801, 
        -46.37687, -46.34601, -46.31462, -46.28178, -46.2478, -46.21212, 
        -46.17405, -46.13581, -46.09698, -46.05832, -46.0203, -45.98255, 
        -45.94474, -45.90606, -45.86587, -45.82335, -45.77772, -45.72771, 
        -45.67375, -45.61679, -45.55681, -45.49443, -45.43004, -45.36522, 
        -45.29905, -45.23148, -45.16104, -45.08723, -45.0091, -44.92538, 
        -44.83805, -44.74887, -44.66049, -44.57657, -44.50066, -44.43525, 
        -44.38174, -44.3404, -44.31097, -44.29182, -44.28131, -44.27663, 
        -44.27823, -44.28334, -44.29142, -44.30285, -44.31727, -44.33416, 
        -44.35299, -44.37334, -44.39503, -44.41737, -44.44009, -44.46301, 
        -44.48718, -44.51339, -44.5425, -44.57542, -44.61297, -44.6553, 
        -44.70191, -44.75284, -44.80606, -44.86055, -44.91608, -44.97294, 
        -45.03261, -45.09705, -45.16857, -45.24908, -45.34007, -45.44389, 
        -45.55928, -45.68853, -45.82962, -45.98254, -46.14581, -46.31899, 
        -46.50063, -46.68968, -46.88422, -47.08191, -47.27966, -47.47424, 
        -47.6635,
  -38.21224, -38.30252, -38.3908, -38.47791, -38.56242, -38.64717, 
        -38.72823, -38.80518, -38.87963, -38.95695, -39.03143, -39.10939, 
        -39.18818, -39.2656, -39.34222, -39.42598, -39.51273, -39.6062, 
        -39.70428, -39.8044, -39.9125, -40.02568, -40.14208, -40.26183, 
        -40.38343, -40.50897, -40.6413, -40.77605, -40.91352, -41.05265, 
        -41.19373, -41.33606, -41.4828, -41.62551, -41.76465, -41.90075, 
        -42.03539, -42.16781, -42.29657, -42.42276, -42.54512, -42.66355, 
        -42.77784, -42.8875, -42.99343, -43.09523, -43.19571, -43.29445, 
        -43.39213, -43.48896, -43.58473, -43.67912, -43.77168, -43.86238, 
        -43.95068, -44.03643, -44.12012, -44.20209, -44.2829, -44.36454, 
        -44.44927, -44.53899, -44.63729, -44.74485, -44.86165, -44.98768, 
        -45.12152, -45.26123, -45.40444, -45.54914, -45.69407, -45.83976, 
        -45.98706, -46.13763, -46.29321, -46.45337, -46.61908, -46.79018, 
        -46.96625, -47.15028, -47.34155, -47.54154, -47.75042, -47.96811, 
        -48.19282, -48.42085, -48.64809, -48.86834, -49.07619, -49.26521, 
        -49.42903, -49.56044, -49.6544, -49.70595, -49.71263, -49.67401, 
        -49.5938, -49.47707, -49.3338, -49.17328, -49.0065, -48.8437, 
        -48.69197, -48.55433, -48.43331, -48.32917, -48.23983, -48.16292, 
        -48.09683, -48.03613, -47.98226, -47.93421, -47.89325, -47.86002, 
        -47.83756, -47.82665, -47.82679, -47.83946, -47.86199, -47.89202, 
        -47.92714, -47.96444, -48.00123, -48.03508, -48.06535, -48.09155, 
        -48.11312, -48.13072, -48.14539, -48.15686, -48.16555, -48.17153, 
        -48.17607, -48.17873, -48.17814, -48.17564, -48.17131, -48.16381, 
        -48.15448, -48.14162, -48.12494, -48.10425, -48.07934, -48.05022, 
        -48.01783, -47.98276, -47.94545, -47.90699, -47.868, -47.82745, 
        -47.7861, -47.74436, -47.70214, -47.6595, -47.61588, -47.57162, 
        -47.52609, -47.47882, -47.43034, -47.37945, -47.32883, -47.27867, 
        -47.22911, -47.1804, -47.1326, -47.08617, -47.0412, -46.99763, 
        -46.95649, -46.91671, -46.87847, -46.84256, -46.80933, -46.77858, 
        -46.75209, -46.72985, -46.71209, -46.6984, -46.68748, -46.67897, 
        -46.67207, -46.66594, -46.66047, -46.65556, -46.64923, -46.64313, 
        -46.63583, -46.62708, -46.6165, -46.6045, -46.591, -46.57639, 
        -46.56079, -46.54447, -46.52791, -46.51191, -46.49599, -46.48115, 
        -46.46758, -46.45456, -46.44168, -46.42829, -46.41397, -46.39833, 
        -46.37988, -46.3586, -46.3344, -46.30676, -46.27627, -46.24366, 
        -46.20969, -46.17467, -46.1415, -46.10981, -46.08006, -46.0523, 
        -46.0261, -46.00029, -45.97438, -45.94725, -45.91834, -45.88758, 
        -45.85512, -45.8213, -45.78713, -45.75291, -45.71943, -45.6865, 
        -45.65329, -45.61917, -45.58302, -45.54408, -45.50202, -45.45573, 
        -45.40521, -45.35148, -45.29473, -45.23554, -45.17455, -45.11269, 
        -45.05007, -44.9855, -44.91816, -44.84816, -44.77242, -44.69284, 
        -44.61067, -44.52743, -44.44551, -44.36813, -44.29847, -44.23866, 
        -44.18977, -44.15176, -44.12371, -44.10449, -44.09251, -44.08591, 
        -44.08395, -44.08541, -44.08987, -44.09819, -44.10964, -44.12425, 
        -44.14116, -44.16014, -44.18074, -44.20237, -44.22459, -44.248, 
        -44.27329, -44.30128, -44.33246, -44.36753, -44.40701, -44.45145, 
        -44.50021, -44.55241, -44.60697, -44.66261, -44.71902, -44.77688, 
        -44.838, -44.90471, -44.97954, -45.06425, -45.16281, -45.27572, 
        -45.40278, -45.54392, -45.69706, -45.86071, -46.03299, -46.21188, 
        -46.39588, -46.58359, -46.77255, -46.96114, -47.14746, -47.32837, 
        -47.50318,
  -38.15491, -38.24349, -38.33022, -38.41339, -38.49586, -38.57677, 
        -38.65649, -38.73415, -38.80634, -38.88222, -38.95643, -39.03354, 
        -39.11018, -39.18696, -39.26252, -39.34544, -39.43143, -39.52074, 
        -39.61582, -39.71332, -39.81741, -39.9257, -40.03812, -40.1545, 
        -40.2742, -40.40038, -40.5284, -40.66136, -40.79539, -40.93408, 
        -41.07426, -41.21535, -41.35806, -41.50245, -41.6416, -41.778, 
        -41.91133, -42.04317, -42.17146, -42.29585, -42.41723, -42.53446, 
        -42.64708, -42.75507, -42.85929, -42.96021, -43.05862, -43.15483, 
        -43.25021, -43.34477, -43.43842, -43.53093, -43.62199, -43.71064, 
        -43.7965, -43.87967, -43.95943, -44.03795, -44.11594, -44.19495, 
        -44.27753, -44.36669, -44.46383, -44.57005, -44.68517, -44.80923, 
        -44.94064, -45.07691, -45.21612, -45.3564, -45.49738, -45.63894, 
        -45.78164, -45.92825, -46.0791, -46.23374, -46.39307, -46.55758, 
        -46.7281, -46.90543, -47.08996, -47.28223, -47.48217, -47.68907, 
        -47.90123, -48.11516, -48.32728, -48.53268, -48.72673, -48.90318, 
        -49.05525, -49.17875, -49.26733, -49.31672, -49.3238, -49.28871, 
        -49.2135, -49.1039, -48.96679, -48.81132, -48.64703, -48.48329, 
        -48.32654, -48.18009, -48.04757, -47.92964, -47.82569, -47.73378, 
        -47.65474, -47.58202, -47.51817, -47.46153, -47.41388, -47.37529, 
        -47.34909, -47.33541, -47.33475, -47.3464, -47.36863, -47.39959, 
        -47.43605, -47.4752, -47.51417, -47.5507, -47.58347, -47.61132, 
        -47.63365, -47.65158, -47.66552, -47.67519, -47.68222, -47.68708, 
        -47.68937, -47.69105, -47.68964, -47.68614, -47.68088, -47.67346, 
        -47.66323, -47.64979, -47.63194, -47.60994, -47.5839, -47.5529, 
        -47.51992, -47.48396, -47.44638, -47.40803, -47.37036, -47.33168, 
        -47.2925, -47.25231, -47.21299, -47.17342, -47.13346, -47.09251, 
        -47.05035, -47.00681, -46.96185, -46.91605, -46.86978, -46.82387, 
        -46.77889, -46.7347, -46.69135, -46.64884, -46.60732, -46.56656, 
        -46.52784, -46.48982, -46.45315, -46.41835, -46.38605, -46.35625, 
        -46.33105, -46.30948, -46.2938, -46.28279, -46.2752, -46.27083, 
        -46.26796, -46.26641, -46.26485, -46.26386, -46.26213, -46.25888, 
        -46.2538, -46.24642, -46.23647, -46.22443, -46.21065, -46.19571, 
        -46.18003, -46.16371, -46.14772, -46.13208, -46.11738, -46.10359, 
        -46.09068, -46.07821, -46.06536, -46.05077, -46.03625, -46.02022, 
        -46.00229, -45.98183, -45.9587, -45.93267, -45.90408, -45.87369, 
        -45.84188, -45.81039, -45.78003, -45.75184, -45.72595, -45.70264, 
        -45.68108, -45.66033, -45.63974, -45.61803, -45.59437, -45.56873, 
        -45.54085, -45.51181, -45.48195, -45.45218, -45.42292, -45.39415, 
        -45.36503, -45.33466, -45.30238, -45.26731, -45.22783, -45.18582, 
        -45.13975, -45.0903, -45.03782, -44.983, -44.92623, -44.86826, 
        -44.80894, -44.74762, -44.68378, -44.61668, -44.54584, -44.47106, 
        -44.39378, -44.31643, -44.24092, -44.1702, -44.10653, -44.05225, 
        -44.0074, -43.97219, -43.94531, -43.92567, -43.91161, -43.9021, 
        -43.89647, -43.89432, -43.89547, -43.90088, -43.90946, -43.92179, 
        -43.93755, -43.95581, -43.97617, -43.99782, -44.02042, -44.04391, 
        -44.07072, -44.10023, -44.13322, -44.17005, -44.21113, -44.25714, 
        -44.30708, -44.36057, -44.41619, -44.47335, -44.53147, -44.59199, 
        -44.6572, -44.72938, -44.81143, -44.9062, -45.01564, -45.14124, 
        -45.28182, -45.43579, -45.60068, -45.77345, -45.95158, -46.13225, 
        -46.31375, -46.49449, -46.67264, -46.84744, -47.01749, -47.18179, 
        -47.33938,
  -38.09667, -38.18521, -38.27053, -38.35142, -38.42952, -38.50678, 
        -38.58487, -38.66475, -38.73972, -38.81343, -38.88667, -38.96329, 
        -39.03923, -39.11335, -39.19029, -39.27142, -39.35556, -39.44396, 
        -39.53601, -39.63107, -39.72953, -39.8325, -39.94157, -40.05508, 
        -40.17366, -40.29668, -40.42337, -40.55466, -40.68863, -40.82439, 
        -40.9639, -41.10499, -41.24606, -41.38869, -41.52698, -41.66288, 
        -41.79663, -41.92856, -42.05714, -42.18214, -42.30357, -42.42053, 
        -42.53168, -42.63818, -42.74062, -42.83973, -42.93573, -43.02943, 
        -43.12185, -43.21379, -43.30395, -43.39472, -43.48417, -43.57105, 
        -43.65551, -43.73632, -43.81398, -43.88976, -43.96524, -44.04223, 
        -44.12355, -44.21168, -44.30807, -44.41284, -44.52623, -44.64734, 
        -44.77347, -44.90487, -45.0386, -45.17364, -45.30969, -45.44751, 
        -45.58767, -45.73056, -45.87626, -46.02509, -46.17733, -46.33427, 
        -46.49759, -46.66781, -46.84534, -47.02974, -47.22029, -47.4154, 
        -47.61265, -47.81131, -48.00744, -48.19712, -48.37616, -48.53942, 
        -48.68165, -48.79725, -48.88119, -48.9292, -48.93889, -48.90957, 
        -48.84291, -48.74342, -48.61605, -48.46946, -48.31026, -48.14896, 
        -47.98719, -47.83187, -47.68713, -47.5541, -47.43385, -47.32637, 
        -47.23259, -47.14758, -47.07284, -47.00745, -46.95194, -46.90737, 
        -46.87666, -46.85971, -46.85637, -46.86577, -46.8865, -46.91652, 
        -46.95269, -46.99215, -47.031, -47.0688, -47.10298, -47.13196, 
        -47.15501, -47.17257, -47.18561, -47.19484, -47.20086, -47.20389, 
        -47.20464, -47.20617, -47.20415, -47.20054, -47.19469, -47.18629, 
        -47.17515, -47.16116, -47.14248, -47.11922, -47.09169, -47.05805, 
        -47.02367, -46.98734, -46.94954, -46.91133, -46.87498, -46.83788, 
        -46.80092, -46.76421, -46.72747, -46.69126, -46.65468, -46.61763, 
        -46.57911, -46.53912, -46.49812, -46.45614, -46.41413, -46.37248, 
        -46.33194, -46.29239, -46.25338, -46.21516, -46.17632, -46.13857, 
        -46.10249, -46.06641, -46.0316, -45.99819, -45.96699, -45.93813, 
        -45.91417, -45.89508, -45.88114, -45.87229, -45.86795, -45.86683, 
        -45.86789, -45.87001, -45.87249, -45.87503, -45.87636, -45.876, 
        -45.87305, -45.8671, -45.85781, -45.84583, -45.83174, -45.81628, 
        -45.79942, -45.78369, -45.76831, -45.75391, -45.74052, -45.72795, 
        -45.7162, -45.70432, -45.69186, -45.67842, -45.66365, -45.64775, 
        -45.63036, -45.61109, -45.58941, -45.56493, -45.53864, -45.51043, 
        -45.48119, -45.45252, -45.4251, -45.40038, -45.37843, -45.35938, 
        -45.34254, -45.32679, -45.31151, -45.29524, -45.27695, -45.25539, 
        -45.23236, -45.20756, -45.18208, -45.15649, -45.13116, -45.10584, 
        -45.0802, -45.05339, -45.02481, -44.99347, -44.95902, -44.92151, 
        -44.88046, -44.83601, -44.78878, -44.73895, -44.68696, -44.63324, 
        -44.57768, -44.51972, -44.45881, -44.39489, -44.32771, -44.25745, 
        -44.18521, -44.11337, -44.04398, -43.97957, -43.92189, -43.87238, 
        -43.83143, -43.79858, -43.77256, -43.75138, -43.73556, -43.72344, 
        -43.71486, -43.70963, -43.70805, -43.71045, -43.71692, -43.72799, 
        -43.74269, -43.76066, -43.7813, -43.80355, -43.82758, -43.85357, 
        -43.88219, -43.91354, -43.94793, -43.986, -44.02834, -44.07502, 
        -44.12597, -44.18041, -44.2377, -44.29679, -44.35894, -44.42414, 
        -44.4966, -44.57799, -44.67073, -44.77695, -44.89955, -45.03965, 
        -45.19535, -45.3626, -45.53773, -45.717, -45.89684, -46.07526, 
        -46.24932, -46.41801, -46.58068, -46.73737, -46.88793, -47.03275, 
        -47.16982,
  -38.03704, -38.12533, -38.21084, -38.29094, -38.36812, -38.44408, 
        -38.51928, -38.59718, -38.6758, -38.74878, -38.81991, -38.89814, 
        -38.97203, -39.04405, -39.12014, -39.20189, -39.28595, -39.37198, 
        -39.46267, -39.55764, -39.65376, -39.74982, -39.85292, -39.96138, 
        -40.07727, -40.19771, -40.32265, -40.45275, -40.58549, -40.72005, 
        -40.85827, -40.99865, -41.14144, -41.28303, -41.42102, -41.55722, 
        -41.69165, -41.82513, -41.95457, -42.08082, -42.2028, -42.31951, 
        -42.43031, -42.53606, -42.63613, -42.73296, -42.82632, -42.91694, 
        -43.00602, -43.0948, -43.18305, -43.2712, -43.35884, -43.44418, 
        -43.52643, -43.60545, -43.68115, -43.7551, -43.82874, -43.90442, 
        -43.98512, -44.07155, -44.16652, -44.26965, -44.37971, -44.49751, 
        -44.61958, -44.74506, -44.8727, -45.0019, -45.13285, -45.26667, 
        -45.40271, -45.54102, -45.68157, -45.82442, -45.96983, -46.11929, 
        -46.27392, -46.43663, -46.60605, -46.78164, -46.96151, -47.14432, 
        -47.32867, -47.5122, -47.69219, -47.86567, -48.02898, -48.17818, 
        -48.3083, -48.41477, -48.49345, -48.54014, -48.55285, -48.53028, 
        -48.47297, -48.38585, -48.27115, -48.13544, -47.98589, -47.828, 
        -47.66706, -47.50637, -47.35013, -47.20339, -47.0673, -46.94324, 
        -46.83411, -46.73547, -46.64886, -46.57401, -46.51064, -46.45974, 
        -46.4244, -46.40213, -46.39532, -46.40176, -46.41917, -46.44653, 
        -46.48021, -46.51794, -46.5567, -46.59356, -46.62775, -46.65653, 
        -46.67943, -46.69633, -46.70835, -46.71659, -46.7211, -46.72259, 
        -46.72214, -46.7226, -46.72042, -46.71618, -46.70911, -46.70029, 
        -46.68872, -46.67422, -46.65499, -46.63105, -46.60218, -46.56759, 
        -46.53276, -46.49598, -46.45835, -46.42081, -46.3856, -46.35015, 
        -46.31547, -46.2809, -46.24668, -46.21303, -46.17966, -46.14598, 
        -46.11086, -46.07436, -46.036, -45.99814, -45.96024, -45.92283, 
        -45.88663, -45.85143, -45.81707, -45.78329, -45.74904, -45.71436, 
        -45.68136, -45.64749, -45.61468, -45.58289, -45.55333, -45.52488, 
        -45.50225, -45.48463, -45.47213, -45.46505, -45.46339, -45.46535, 
        -45.4697, -45.47519, -45.4813, -45.48571, -45.49025, -45.49168, 
        -45.49074, -45.48553, -45.47629, -45.46447, -45.45016, -45.43494, 
        -45.41917, -45.40403, -45.39001, -45.37745, -45.36581, -45.35524, 
        -45.34487, -45.33448, -45.3231, -45.31024, -45.29603, -45.28069, 
        -45.26413, -45.24601, -45.22594, -45.20364, -45.1795, -45.15421, 
        -45.12694, -45.1015, -45.07771, -45.05656, -45.03877, -45.02379, 
        -45.01149, -45.0005, -44.99007, -44.97903, -44.966, -44.95043, 
        -44.93223, -44.91198, -44.89081, -44.86913, -44.84747, -44.8257, 
        -44.80329, -44.77996, -44.75474, -44.72709, -44.69695, -44.66423, 
        -44.62813, -44.58901, -44.54742, -44.50298, -44.45618, -44.40716, 
        -44.35559, -44.30096, -44.24164, -44.18052, -44.11645, -44.04998, 
        -43.98209, -43.91526, -43.85142, -43.79271, -43.74077, -43.69602, 
        -43.65876, -43.62828, -43.60312, -43.5825, -43.56509, -43.55085, 
        -43.53952, -43.53178, -43.52816, -43.52869, -43.53365, -43.54388, 
        -43.55852, -43.57703, -43.5985, -43.6223, -43.64853, -43.67655, 
        -43.70692, -43.73946, -43.77442, -43.81313, -43.85577, -43.90298, 
        -43.95525, -44.01083, -44.07074, -44.13433, -44.20143, -44.27483, 
        -44.35651, -44.45015, -44.55564, -44.67607, -44.81388, -44.96992, 
        -45.13991, -45.31848, -45.5012, -45.68323, -45.86089, -46.03205, 
        -46.1943, -46.34757, -46.49194, -46.62894, -46.75859, -46.88267, 
        -47.00087,
  -37.97752, -38.06516, -38.15293, -38.2331, -38.30891, -38.38391, 
        -38.45714, -38.53294, -38.60983, -38.68707, -38.75746, -38.83105, 
        -38.90269, -38.97696, -39.05494, -39.137, -39.22138, -39.30772, 
        -39.3965, -39.48739, -39.57658, -39.67032, -39.76872, -39.87209, 
        -39.98338, -40.10306, -40.22567, -40.35423, -40.48709, -40.62099, 
        -40.75765, -40.89756, -41.0416, -41.18667, -41.32444, -41.45975, 
        -41.59511, -41.73064, -41.86169, -41.98851, -42.112, -42.22942, 
        -42.34087, -42.44618, -42.54631, -42.64109, -42.73164, -42.81887, 
        -42.90414, -42.98893, -43.07414, -43.15988, -43.24513, -43.32883, 
        -43.40926, -43.48532, -43.55914, -43.63169, -43.70437, -43.77935, 
        -43.8596, -43.94596, -44.03985, -44.14024, -44.24705, -44.35985, 
        -44.47644, -44.59576, -44.71672, -44.84007, -44.9659, -45.09494, 
        -45.22577, -45.35952, -45.49467, -45.63067, -45.76892, -45.91109, 
        -46.05885, -46.21328, -46.37404, -46.53984, -46.70864, -46.879, 
        -47.04919, -47.21714, -47.38089, -47.53746, -47.6846, -47.81763, 
        -47.93389, -48.02935, -48.10125, -48.1456, -48.16082, -48.14533, 
        -48.09996, -48.0259, -47.9253, -47.80344, -47.66532, -47.51476, 
        -47.356, -47.19173, -47.02753, -46.8694, -46.71957, -46.57985, 
        -46.45573, -46.34385, -46.24551, -46.16128, -46.09108, -46.0341, 
        -45.99358, -45.96849, -45.95734, -45.95897, -45.972, -45.99458, 
        -46.02439, -46.05871, -46.09426, -46.12866, -46.16081, -46.18838, 
        -46.21031, -46.22649, -46.23662, -46.24323, -46.24643, -46.24689, 
        -46.2454, -46.24564, -46.24228, -46.23799, -46.2316, -46.22288, 
        -46.21094, -46.19565, -46.17582, -46.15097, -46.12123, -46.08527, 
        -46.04934, -46.0122, -45.97467, -45.93789, -45.90399, -45.87016, 
        -45.8357, -45.8033, -45.77158, -45.74014, -45.70908, -45.67796, 
        -45.64574, -45.61259, -45.57884, -45.54461, -45.51059, -45.4774, 
        -45.4455, -45.41469, -45.38464, -45.35481, -45.32459, -45.29379, 
        -45.26372, -45.2328, -45.20194, -45.17197, -45.14351, -45.11685, 
        -45.0944, -45.07722, -45.06574, -45.05981, -45.06035, -45.06442, 
        -45.07164, -45.08055, -45.08966, -45.09719, -45.10409, -45.10771, 
        -45.10803, -45.10284, -45.09452, -45.08303, -45.06836, -45.05259, 
        -45.03749, -45.02409, -45.01147, -45.0012, -44.9922, -44.98416, 
        -44.97599, -44.96772, -44.95706, -44.94623, -44.9332, -44.91909, 
        -44.90386, -44.88717, -44.86893, -44.84907, -44.82784, -44.80542, 
        -44.78289, -44.76118, -44.74128, -44.72429, -44.71036, -44.6995, 
        -44.69145, -44.6851, -44.67955, -44.67327, -44.66514, -44.65437, 
        -44.64162, -44.62622, -44.60907, -44.59141, -44.57328, -44.55492, 
        -44.53585, -44.5154, -44.49245, -44.46856, -44.44235, -44.41378, 
        -44.38251, -44.34874, -44.31263, -44.27393, -44.23255, -44.18793, 
        -44.14001, -44.08871, -44.03394, -43.97517, -43.91335, -43.84975, 
        -43.78547, -43.72306, -43.66442, -43.61107, -43.56442, -43.52417, 
        -43.49027, -43.46197, -43.43814, -43.41721, -43.39896, -43.38326, 
        -43.37043, -43.36097, -43.3558, -43.35519, -43.35989, -43.37006, 
        -43.38493, -43.4038, -43.42775, -43.45243, -43.48088, -43.51125, 
        -43.54353, -43.57712, -43.61271, -43.65142, -43.69432, -43.74227, 
        -43.79537, -43.85425, -43.91859, -43.98753, -44.06351, -44.14813, 
        -44.24302, -44.34961, -44.46925, -44.60575, -44.76066, -44.93165, 
        -45.11391, -45.30078, -45.4872, -45.6675, -45.8384, -45.99824, 
        -46.14536, -46.28062, -46.40508, -46.52108, -46.63028, -46.734, 
        -46.83219,
  -37.91904, -38.0087, -38.09562, -38.17427, -38.25255, -38.32792, 
        -38.40185, -38.47566, -38.54981, -38.62655, -38.69426, -38.76424, 
        -38.83773, -38.91317, -38.99247, -39.07435, -39.15828, -39.24392, 
        -39.32992, -39.41771, -39.5045, -39.59351, -39.68704, -39.78746, 
        -39.89572, -40.01208, -40.13662, -40.26417, -40.39467, -40.52806, 
        -40.66489, -40.80345, -40.94704, -41.09147, -41.23165, -41.36955, 
        -41.50543, -41.64293, -41.77667, -41.90678, -42.03189, -42.15076, 
        -42.26297, -42.3688, -42.46851, -42.56178, -42.64965, -42.73351, 
        -42.81546, -42.89552, -42.97758, -43.06036, -43.14332, -43.22483, 
        -43.3031, -43.37793, -43.44988, -43.52074, -43.59275, -43.66735, 
        -43.74704, -43.8325, -43.92409, -44.02201, -44.12547, -44.23292, 
        -44.34247, -44.4554, -44.57018, -44.68737, -44.80774, -44.93171, 
        -45.05811, -45.18649, -45.31563, -45.44508, -45.57603, -45.71035, 
        -45.85009, -45.99593, -46.1473, -46.3027, -46.46023, -46.61687, 
        -46.77276, -46.92537, -47.07253, -47.21243, -47.3415, -47.45906, 
        -47.56031, -47.64261, -47.70557, -47.74646, -47.76207, -47.75257, 
        -47.71696, -47.65569, -47.56968, -47.46232, -47.33685, -47.19552, 
        -47.04079, -46.87559, -46.70798, -46.54219, -46.3809, -46.23059, 
        -46.09644, -45.97314, -45.86541, -45.77358, -45.69823, -45.63718, 
        -45.59285, -45.56297, -45.54585, -45.54142, -45.54792, -45.56377, 
        -45.58887, -45.61672, -45.64751, -45.67694, -45.70568, -45.7307, 
        -45.75102, -45.76628, -45.77662, -45.78196, -45.78452, -45.78413, 
        -45.78251, -45.78262, -45.77908, -45.77456, -45.76793, -45.75886, 
        -45.74584, -45.72953, -45.7083, -45.68206, -45.64996, -45.61147, 
        -45.57429, -45.53611, -45.49863, -45.46217, -45.42994, -45.39686, 
        -45.36478, -45.3338, -45.30361, -45.27338, -45.24394, -45.2143, 
        -45.18447, -45.15424, -45.12417, -45.0935, -45.06352, -45.03458, 
        -45.00722, -44.98054, -44.95492, -44.92844, -44.90251, -44.8762, 
        -44.85069, -44.82247, -44.79444, -44.76675, -44.74004, -44.71289, 
        -44.69199, -44.67562, -44.66478, -44.66019, -44.66349, -44.66969, 
        -44.67944, -44.6912, -44.70331, -44.71322, -44.72128, -44.72569, 
        -44.72688, -44.72229, -44.71269, -44.70055, -44.6863, -44.67068, 
        -44.65642, -44.64361, -44.63318, -44.62518, -44.61918, -44.61446, 
        -44.61019, -44.6043, -44.59725, -44.58869, -44.57822, -44.56605, 
        -44.55204, -44.53725, -44.52127, -44.50449, -44.48642, -44.46762, 
        -44.44912, -44.43171, -44.41612, -44.40343, -44.39369, -44.38697, 
        -44.38311, -44.3811, -44.3798, -44.37721, -44.37444, -44.36866, 
        -44.36111, -44.35072, -44.33815, -44.32431, -44.30982, -44.29476, 
        -44.27873, -44.26117, -44.24207, -44.22125, -44.19848, -44.17371, 
        -44.14654, -44.11739, -44.08638, -44.05271, -44.01633, -43.97633, 
        -43.93233, -43.88395, -43.83149, -43.77467, -43.71457, -43.65326, 
        -43.59215, -43.53387, -43.48021, -43.43203, -43.39008, -43.35402, 
        -43.3237, -43.29662, -43.2738, -43.25324, -43.2348, -43.21851, 
        -43.20511, -43.19524, -43.18972, -43.1894, -43.19501, -43.20622, 
        -43.22241, -43.24295, -43.2682, -43.29705, -43.32787, -43.36044, 
        -43.39371, -43.42793, -43.46449, -43.50394, -43.54758, -43.59684, 
        -43.65301, -43.7165, -43.78661, -43.86422, -43.95045, -44.04714, 
        -44.15528, -44.27604, -44.41173, -44.56571, -44.73577, -44.91911, 
        -45.10929, -45.30016, -45.48577, -45.66003, -45.82048, -45.96524, 
        -46.09494, -46.21073, -46.31547, -46.41162, -46.50028, -46.58484, 
        -46.66466,
  -37.86575, -37.95483, -38.04022, -38.12111, -38.20029, -38.27664, 
        -38.35207, -38.42437, -38.49624, -38.56888, -38.63493, -38.70412, 
        -38.77698, -38.85068, -38.93034, -39.01281, -39.09567, -39.17876, 
        -39.26529, -39.35223, -39.43734, -39.5216, -39.61224, -39.70965, 
        -39.81488, -39.92838, -40.05038, -40.17922, -40.30929, -40.44157, 
        -40.57675, -40.71459, -40.85387, -40.99966, -41.14291, -41.2848, 
        -41.42468, -41.56381, -41.70045, -41.83283, -41.96012, -42.08071, 
        -42.19458, -42.30143, -42.40009, -42.49258, -42.57861, -42.65996, 
        -42.73862, -42.81679, -42.89552, -42.97576, -43.056, -43.13477, 
        -43.21019, -43.28239, -43.35237, -43.42171, -43.4924, -43.56619, 
        -43.64367, -43.72767, -43.81696, -43.91177, -44.0113, -44.11366, 
        -44.21885, -44.32544, -44.43421, -44.54552, -44.66016, -44.77795, 
        -44.89816, -45.01992, -45.14225, -45.26525, -45.38908, -45.51493, 
        -45.64652, -45.78349, -45.92493, -46.06939, -46.21502, -46.35989, 
        -46.50171, -46.6386, -46.76939, -46.89114, -47.00261, -47.10114, 
        -47.18525, -47.25343, -47.30574, -47.33995, -47.35482, -47.34786, 
        -47.32003, -47.26987, -47.1971, -47.1038, -46.991, -46.86005, 
        -46.71344, -46.55259, -46.38543, -46.21549, -46.04725, -45.88863, 
        -45.74529, -45.61393, -45.49842, -45.40163, -45.32275, -45.25921, 
        -45.21142, -45.17659, -45.15301, -45.14061, -45.13818, -45.14558, 
        -45.16247, -45.18602, -45.21189, -45.23582, -45.26017, -45.28213, 
        -45.30034, -45.3146, -45.32351, -45.3287, -45.33031, -45.32912, 
        -45.3271, -45.32695, -45.32397, -45.31758, -45.31003, -45.30011, 
        -45.2865, -45.26907, -45.24678, -45.21854, -45.18621, -45.14696, 
        -45.11029, -45.07267, -45.03452, -44.99828, -44.96662, -44.93368, 
        -44.90239, -44.87179, -44.84247, -44.81227, -44.78323, -44.7544, 
        -44.72526, -44.69733, -44.67056, -44.6437, -44.61775, -44.59283, 
        -44.56951, -44.54692, -44.52553, -44.50425, -44.48252, -44.45984, 
        -44.43801, -44.41349, -44.38848, -44.36346, -44.33915, -44.3136, 
        -44.29367, -44.2778, -44.26717, -44.26289, -44.26703, -44.27415, 
        -44.28534, -44.29744, -44.31076, -44.32194, -44.33125, -44.33708, 
        -44.33811, -44.33458, -44.32586, -44.31441, -44.30142, -44.28765, 
        -44.27525, -44.26545, -44.25792, -44.25317, -44.25058, -44.24973, 
        -44.24924, -44.24755, -44.2438, -44.23808, -44.23038, -44.22041, 
        -44.20937, -44.19675, -44.18349, -44.1699, -44.15577, -44.14061, 
        -44.12651, -44.11353, -44.10283, -44.09453, -44.08932, -44.08665, 
        -44.08654, -44.08858, -44.09166, -44.0949, -44.09685, -44.09621, 
        -44.09391, -44.08843, -44.08069, -44.07103, -44.06001, -44.04817, 
        -44.03503, -44.02021, -44.00336, -43.9848, -43.96444, -43.94212, 
        -43.91808, -43.89241, -43.8651, -43.83574, -43.80361, -43.7678, 
        -43.7277, -43.68198, -43.63234, -43.57788, -43.52068, -43.46206, 
        -43.40406, -43.34961, -43.30037, -43.25718, -43.21983, -43.18805, 
        -43.161, -43.13759, -43.11638, -43.09677, -43.07855, -43.06237, 
        -43.04903, -43.03952, -43.03483, -43.03574, -43.04307, -43.05613, 
        -43.07426, -43.09753, -43.12458, -43.15561, -43.18761, -43.22231, 
        -43.2571, -43.29271, -43.33058, -43.37106, -43.41595, -43.46812, 
        -43.52797, -43.59848, -43.67739, -43.76571, -43.86291, -43.97218, 
        -44.09406, -44.23055, -44.38356, -44.55155, -44.73296, -44.92391, 
        -45.11764, -45.30705, -45.48604, -45.65003, -45.79631, -45.92459, 
        -46.03615, -46.13335, -46.21972, -46.29787, -46.37016, -46.43719, 
        -46.50039,
  -37.82333, -37.91127, -37.99621, -38.07734, -38.15685, -38.23398, 
        -38.30854, -38.37943, -38.44945, -38.51851, -38.58031, -38.64792, 
        -38.71888, -38.79189, -38.87115, -38.95202, -39.03333, -39.11535, 
        -39.19994, -39.28596, -39.37114, -39.45288, -39.54388, -39.63949, 
        -39.74287, -39.85359, -39.97234, -40.09647, -40.22662, -40.3604, 
        -40.49723, -40.63472, -40.77369, -40.91606, -41.06357, -41.20797, 
        -41.35077, -41.49253, -41.63018, -41.76506, -41.89421, -42.01669, 
        -42.13245, -42.24049, -42.34105, -42.43365, -42.5193, -42.59937, 
        -42.67637, -42.75214, -42.8287, -42.90611, -42.98338, -43.0588, 
        -43.13013, -43.19912, -43.26623, -43.33361, -43.40218, -43.47411, 
        -43.55027, -43.63174, -43.71846, -43.80988, -43.90542, -44.00363, 
        -44.10347, -44.20467, -44.30755, -44.41301, -44.5214, -44.63162, 
        -44.7448, -44.85937, -44.97429, -45.08996, -45.20665, -45.32589, 
        -45.44916, -45.57691, -45.70814, -45.84145, -45.9752, -46.10695, 
        -46.23456, -46.35588, -46.46951, -46.5732, -46.66492, -46.74269, 
        -46.8085, -46.86095, -46.9005, -46.92695, -46.93864, -46.93457, 
        -46.91283, -46.87147, -46.80932, -46.72777, -46.62645, -46.5057, 
        -46.36737, -46.21211, -46.04759, -45.87817, -45.70897, -45.54549, 
        -45.39772, -45.26039, -45.13968, -45.03716, -44.95168, -44.88724, 
        -44.83857, -44.80094, -44.77166, -44.75196, -44.74105, -44.739, 
        -44.74631, -44.76266, -44.77957, -44.79818, -44.81711, -44.83619, 
        -44.85316, -44.86593, -44.87475, -44.87906, -44.88126, -44.88032, 
        -44.87844, -44.8788, -44.8762, -44.87157, -44.86442, -44.85308, 
        -44.83673, -44.8176, -44.79258, -44.76223, -44.73043, -44.69088, 
        -44.65471, -44.6174, -44.57896, -44.54255, -44.5117, -44.47813, 
        -44.44679, -44.41593, -44.386, -44.3536, -44.32242, -44.29247, 
        -44.26493, -44.24099, -44.21825, -44.19617, -44.17493, -44.15477, 
        -44.13551, -44.11666, -44.09917, -44.08224, -44.06558, -44.04721, 
        -44.02932, -44.00831, -43.98684, -43.96489, -43.94339, -43.91898, 
        -43.90057, -43.88584, -43.87588, -43.87178, -43.87595, -43.88315, 
        -43.89468, -43.90808, -43.9216, -43.93249, -43.94224, -43.94859, 
        -43.95055, -43.94825, -43.94129, -43.93158, -43.92024, -43.90867, 
        -43.89871, -43.89212, -43.8882, -43.88733, -43.88908, -43.89244, 
        -43.8963, -43.89758, -43.89793, -43.89574, -43.89109, -43.88428, 
        -43.87598, -43.86662, -43.85677, -43.847, -43.83726, -43.82751, 
        -43.81851, -43.81054, -43.80455, -43.80111, -43.80009, -43.80176, 
        -43.80572, -43.81196, -43.81929, -43.8269, -43.8334, -43.83785, 
        -43.84003, -43.83943, -43.83607, -43.83054, -43.8231, -43.81431, 
        -43.80385, -43.79021, -43.77525, -43.75845, -43.73954, -43.7186, 
        -43.69642, -43.67295, -43.64817, -43.62186, -43.59303, -43.56078, 
        -43.52446, -43.48338, -43.4371, -43.38646, -43.33231, -43.27702, 
        -43.22292, -43.17271, -43.12765, -43.08913, -43.05642, -43.02877, 
        -43.0051, -42.98451, -42.96514, -42.9467, -42.92941, -42.91384, 
        -42.90129, -42.8928, -42.88961, -42.89301, -42.90297, -42.91868, 
        -42.93923, -42.9625, -42.99253, -43.02554, -43.06006, -43.09674, 
        -43.13504, -43.17294, -43.21145, -43.25417, -43.30256, -43.35668, 
        -43.41488, -43.50227, -43.59387, -43.69218, -43.80289, -43.92792, 
        -44.06504, -44.21643, -44.3817, -44.55958, -44.74711, -44.93954, 
        -45.13045, -45.31275, -45.48085, -45.63084, -45.76136, -45.87287, 
        -45.96738, -46.04795, -46.118, -46.18065, -46.23787, -46.2899, 
        -46.33796,
  -37.7943, -37.87973, -37.96462, -38.04452, -38.12348, -38.19941, 
        -38.27295, -38.34113, -38.40893, -38.46922, -38.53125, -38.59607, 
        -38.6644, -38.73595, -38.81283, -38.89267, -38.97256, -39.0521, 
        -39.13362, -39.21674, -39.30211, -39.38916, -39.47805, -39.57494, 
        -39.67807, -39.78875, -39.90622, -40.02979, -40.15741, -40.2888, 
        -40.423, -40.55958, -40.70161, -40.84524, -40.99273, -41.13913, 
        -41.28419, -41.42705, -41.56794, -41.70438, -41.83511, -41.95965, 
        -42.07681, -42.18671, -42.28932, -42.38312, -42.46944, -42.54974, 
        -42.62633, -42.69998, -42.77492, -42.84983, -42.92395, -42.99545, 
        -43.06382, -43.12875, -43.19256, -43.25684, -43.32281, -43.39199, 
        -43.46522, -43.5437, -43.62698, -43.71499, -43.80686, -43.89976, 
        -43.99492, -44.09109, -44.18862, -44.28787, -44.38972, -44.49337, 
        -44.59862, -44.70545, -44.81274, -44.92078, -45.03003, -45.14177, 
        -45.25677, -45.37503, -45.49579, -45.61758, -45.73792, -45.8564, 
        -45.96978, -46.07594, -46.1725, -46.25754, -46.32949, -46.38832, 
        -46.43468, -46.47001, -46.49582, -46.51249, -46.51984, -46.51506, 
        -46.49724, -46.46143, -46.40737, -46.33526, -46.24427, -46.13163, 
        -46.00143, -45.85328, -45.69537, -45.53074, -45.364, -45.2019, 
        -45.05431, -44.91431, -44.78811, -44.67763, -44.59547, -44.53036, 
        -44.48073, -44.44099, -44.40834, -44.38315, -44.36376, -44.35294, 
        -44.34834, -44.35106, -44.35735, -44.36544, -44.37615, -44.39429, 
        -44.41159, -44.42279, -44.43373, -44.44044, -44.44562, -44.44447, 
        -44.44209, -44.44302, -44.44109, -44.43699, -44.42875, -44.41631, 
        -44.39943, -44.37856, -44.35161, -44.31916, -44.28619, -44.24706, 
        -44.21114, -44.17452, -44.13527, -44.09743, -44.06656, -44.03316, 
        -43.99964, -43.96713, -43.93488, -43.90108, -43.86779, -43.83833, 
        -43.81312, -43.79144, -43.77273, -43.75439, -43.7368, -43.72117, 
        -43.70617, -43.69154, -43.67731, -43.6652, -43.65344, -43.63997, 
        -43.62592, -43.6092, -43.59125, -43.57227, -43.55323, -43.53234, 
        -43.5159, -43.50377, -43.49564, -43.49236, -43.49644, -43.5027, 
        -43.5145, -43.52717, -43.53839, -43.54756, -43.55695, -43.56359, 
        -43.56689, -43.56649, -43.56266, -43.55446, -43.54602, -43.53764, 
        -43.53082, -43.52788, -43.52835, -43.53173, -43.53791, -43.54581, 
        -43.55402, -43.56086, -43.56547, -43.56722, -43.56599, -43.56246, 
        -43.55724, -43.55144, -43.54522, -43.53965, -43.53461, -43.53028, 
        -43.5266, -43.52405, -43.52302, -43.52438, -43.52769, -43.53365, 
        -43.54134, -43.55088, -43.56102, -43.57246, -43.5831, -43.59174, 
        -43.59792, -43.60166, -43.60254, -43.60092, -43.597, -43.59122, 
        -43.58331, -43.57286, -43.5597, -43.54373, -43.52551, -43.50518, 
        -43.48378, -43.46131, -43.43785, -43.41367, -43.38759, -43.35872, 
        -43.32615, -43.289, -43.24659, -43.20021, -43.15001, -43.09909, 
        -43.04946, -43.00374, -42.96283, -42.92895, -42.90084, -42.8773, 
        -42.85604, -42.83815, -42.82026, -42.80309, -42.78715, -42.77298, 
        -42.76217, -42.7552, -42.75388, -42.75948, -42.7724, -42.79094, 
        -42.81323, -42.83943, -42.87148, -42.90772, -42.93961, -42.98376, 
        -43.02774, -43.07081, -43.11294, -43.15997, -43.21422, -43.27189, 
        -43.32937, -43.43769, -43.54144, -43.65495, -43.77838, -43.91399, 
        -44.06315, -44.22492, -44.39854, -44.58135, -44.76919, -44.95708, 
        -45.139, -45.30876, -45.46171, -45.59517, -45.70893, -45.80438, 
        -45.88414, -45.95013, -46.00762, -46.05827, -46.1034, -46.14357, 
        -46.17935,
  -37.78122, -37.8641, -37.94673, -38.02445, -38.10406, -38.17805, 
        -38.24688, -38.31287, -38.37284, -38.43067, -38.48985, -38.55134, 
        -38.61573, -38.68405, -38.75642, -38.83319, -38.90932, -38.98573, 
        -39.07033, -39.15298, -39.2366, -39.32474, -39.4165, -39.51096, 
        -39.61386, -39.72601, -39.84567, -39.97059, -40.09946, -40.23157, 
        -40.365, -40.50011, -40.64028, -40.7837, -40.93332, -41.0796, 
        -41.22659, -41.37077, -41.51148, -41.64939, -41.78201, -41.90907, 
        -42.02855, -42.13924, -42.24353, -42.33949, -42.42719, -42.50853, 
        -42.58556, -42.66035, -42.73405, -42.80697, -42.87791, -42.94547, 
        -43.00969, -43.07077, -43.13074, -43.19162, -43.25402, -43.31882, 
        -43.38813, -43.46277, -43.54236, -43.62617, -43.71394, -43.8036, 
        -43.89437, -43.9856, -44.07777, -44.17112, -44.26576, -44.36189, 
        -44.45893, -44.55751, -44.65697, -44.75742, -44.85784, -44.96119, 
        -45.0676, -45.17599, -45.28617, -45.39631, -45.50549, -45.61072, 
        -45.70985, -45.80083, -45.88045, -45.94695, -45.99985, -46.03926, 
        -46.06748, -46.08574, -46.09867, -46.10431, -46.10446, -46.0979, 
        -46.0796, -46.0479, -45.99893, -45.93329, -45.84943, -45.7451, 
        -45.6227, -45.48224, -45.33196, -45.17373, -45.01287, -44.85548, 
        -44.71177, -44.57328, -44.44476, -44.33296, -44.24771, -44.18068, 
        -44.12847, -44.08737, -44.05299, -44.02536, -44.00146, -43.98439, 
        -43.97306, -43.96732, -43.96503, -43.96198, -43.96451, -43.9729, 
        -43.98418, -43.99474, -44.00445, -44.01141, -44.01881, -44.01864, 
        -44.01609, -44.01771, -44.01304, -44.0063, -43.99869, -43.98814, 
        -43.97066, -43.94922, -43.92182, -43.88991, -43.85578, -43.81574, 
        -43.77898, -43.74206, -43.70456, -43.6681, -43.63526, -43.59879, 
        -43.56093, -43.52488, -43.49238, -43.45823, -43.4265, -43.39807, 
        -43.37453, -43.35471, -43.33836, -43.32187, -43.3069, -43.29558, 
        -43.28436, -43.27519, -43.26701, -43.26044, -43.2537, -43.24452, 
        -43.23398, -43.22093, -43.20583, -43.18941, -43.17348, -43.15557, 
        -43.14265, -43.13274, -43.12773, -43.1261, -43.13018, -43.13628, 
        -43.14531, -43.15546, -43.16362, -43.16875, -43.1757, -43.18127, 
        -43.18572, -43.18985, -43.19166, -43.18883, -43.1846, -43.18036, 
        -43.17834, -43.17989, -43.18434, -43.1929, -43.20434, -43.21654, 
        -43.22878, -43.24034, -43.24911, -43.25465, -43.25718, -43.2569, 
        -43.255, -43.25259, -43.25096, -43.25012, -43.24879, -43.24968, 
        -43.25134, -43.25399, -43.25788, -43.26377, -43.27144, -43.28095, 
        -43.29219, -43.30541, -43.31952, -43.33361, -43.34719, -43.3592, 
        -43.36902, -43.37638, -43.381, -43.38275, -43.38231, -43.37981, 
        -43.37492, -43.36647, -43.35472, -43.33978, -43.32203, -43.30166, 
        -43.28049, -43.25813, -43.23518, -43.2126, -43.18856, -43.16152, 
        -43.13259, -43.0997, -43.06168, -43.02118, -42.97579, -42.92954, 
        -42.88538, -42.84473, -42.8084, -42.77914, -42.7546, -42.73524, 
        -42.71907, -42.70347, -42.684, -42.66671, -42.65362, -42.64415, 
        -42.63662, -42.63174, -42.63186, -42.63861, -42.65289, -42.67304, 
        -42.69697, -42.72668, -42.75766, -42.80359, -42.84389, -42.89403, 
        -42.94178, -42.99061, -43.03798, -43.09169, -43.15428, -43.22503, 
        -43.30777, -43.41322, -43.52532, -43.64735, -43.78022, -43.92562, 
        -44.082, -44.2495, -44.42543, -44.60677, -44.78843, -44.966, 
        -45.13404, -45.2877, -45.42311, -45.53954, -45.63713, -45.71848, 
        -45.78569, -45.84222, -45.89042, -45.93245, -45.96877, -46.00029, 
        -46.02699,
  -37.78857, -37.86806, -37.94913, -38.02562, -38.09889, -38.16832, 
        -38.23238, -38.29333, -38.34857, -38.40369, -38.45934, -38.51641, 
        -38.57784, -38.64037, -38.70979, -38.78137, -38.85479, -38.93053, 
        -39.01218, -39.09513, -39.17823, -39.26187, -39.35013, -39.4485, 
        -39.55303, -39.66498, -39.78897, -39.91785, -40.04971, -40.18217, 
        -40.31831, -40.45399, -40.59314, -40.73428, -40.88235, -41.03169, 
        -41.17822, -41.32092, -41.46272, -41.59977, -41.73507, -41.86363, 
        -41.98538, -42.09957, -42.2058, -42.30366, -42.39296, -42.47594, 
        -42.55416, -42.6294, -42.70265, -42.77373, -42.84184, -42.90588, 
        -42.9649, -43.02207, -43.07847, -43.1355, -43.19427, -43.25586, 
        -43.32104, -43.39098, -43.46582, -43.54537, -43.62841, -43.71374, 
        -43.80009, -43.88658, -43.9732, -44.06014, -44.14676, -44.23505, 
        -44.32396, -44.41405, -44.50537, -44.59755, -44.69118, -44.78615, 
        -44.88348, -44.98187, -45.081, -45.17966, -45.27635, -45.36873, 
        -45.45403, -45.52996, -45.59386, -45.64299, -45.67681, -45.69873, 
        -45.70897, -45.71266, -45.713, -45.70992, -45.70341, -45.69266, 
        -45.67285, -45.64161, -45.59615, -45.53413, -45.45452, -45.35513, 
        -45.23891, -45.10513, -44.96237, -44.81159, -44.65867, -44.50785, 
        -44.37105, -44.23914, -44.11579, -43.99832, -43.91043, -43.84223, 
        -43.79007, -43.7464, -43.70961, -43.6772, -43.64802, -43.62526, 
        -43.6095, -43.59718, -43.58866, -43.57949, -43.57677, -43.57799, 
        -43.58075, -43.5864, -43.5933, -43.59779, -43.60245, -43.60412, 
        -43.60189, -43.59898, -43.59222, -43.58303, -43.5744, -43.56545, 
        -43.54837, -43.5263, -43.49796, -43.46491, -43.42677, -43.39212, 
        -43.35433, -43.31892, -43.28439, -43.24936, -43.21668, -43.17852, 
        -43.1363, -43.09879, -43.06293, -43.0278, -42.99747, -42.9705, 
        -42.94864, -42.93026, -42.91619, -42.90235, -42.89133, -42.88262, 
        -42.87802, -42.87436, -42.87176, -42.86831, -42.86506, -42.85896, 
        -42.85057, -42.84118, -42.82906, -42.81459, -42.8004, -42.78903, 
        -42.77906, -42.77165, -42.76788, -42.76929, -42.77393, -42.77818, 
        -42.7867, -42.79395, -42.79868, -42.79697, -42.80261, -42.80639, 
        -42.80962, -42.81434, -42.82229, -42.8276, -42.83065, -42.83415, 
        -42.83943, -42.84711, -42.85787, -42.87216, -42.88868, -42.9059, 
        -42.92256, -42.93816, -42.95164, -42.96121, -42.96736, -42.97011, 
        -42.97149, -42.97316, -42.97524, -42.97879, -42.98317, -42.98965, 
        -42.99625, -43.00374, -43.01228, -43.02221, -43.03373, -43.04665, 
        -43.06082, -43.0769, -43.09321, -43.1095, -43.12528, -43.13919, 
        -43.15151, -43.16168, -43.17, -43.17552, -43.17836, -43.17924, 
        -43.17582, -43.17002, -43.15997, -43.14608, -43.12902, -43.10843, 
        -43.08707, -43.06484, -43.04238, -43.02076, -42.99971, -42.97699, 
        -42.95263, -42.92459, -42.89275, -42.8585, -42.81908, -42.77868, 
        -42.73989, -42.70449, -42.67132, -42.6459, -42.62537, -42.60986, 
        -42.59666, -42.58254, -42.56228, -42.53566, -42.52752, -42.52964, 
        -42.52575, -42.52325, -42.5224, -42.52581, -42.53506, -42.56105, 
        -42.58892, -42.62122, -42.65924, -42.71799, -42.77254, -42.82454, 
        -42.88017, -42.93331, -42.98759, -43.04922, -43.12135, -43.20771, 
        -43.30558, -43.41615, -43.53746, -43.66799, -43.80784, -43.95792, 
        -44.11709, -44.2844, -44.45668, -44.63025, -44.80042, -44.96292, 
        -45.11321, -45.2483, -45.36541, -45.4649, -45.54837, -45.61795, 
        -45.67593, -45.7255, -45.76819, -45.80499, -45.83638, -45.86207, 
        -45.88261,
  -37.81939, -37.89603, -37.97256, -38.04601, -38.11452, -38.17736, 
        -38.23627, -38.29016, -38.33891, -38.3887, -38.43921, -38.49141, 
        -38.5478, -38.60697, -38.67009, -38.73722, -38.80988, -38.88117, 
        -38.95802, -39.04046, -39.12265, -39.20645, -39.29592, -39.39376, 
        -39.50005, -39.6137, -39.73573, -39.86715, -40.0024, -40.13773, 
        -40.27394, -40.41461, -40.55438, -40.6968, -40.84423, -40.99177, 
        -41.13746, -41.28053, -41.42204, -41.56068, -41.69631, -41.82695, 
        -41.95061, -42.0669, -42.17469, -42.27385, -42.36465, -42.44886, 
        -42.52736, -42.60323, -42.6763, -42.74623, -42.81165, -42.87281, 
        -42.92965, -42.98334, -43.0359, -43.08898, -43.14385, -43.20132, 
        -43.26191, -43.32674, -43.39603, -43.47039, -43.54694, -43.6278, 
        -43.70954, -43.79077, -43.87191, -43.95251, -44.03301, -44.11356, 
        -44.19419, -44.27591, -44.35901, -44.44275, -44.52795, -44.61426, 
        -44.70184, -44.79043, -44.87875, -44.96614, -45.04997, -45.12988, 
        -45.20199, -45.26363, -45.31269, -45.34668, -45.36547, -45.37122, 
        -45.36852, -45.35957, -45.34853, -45.33689, -45.32401, -45.30833, 
        -45.28613, -45.25371, -45.20836, -45.14737, -45.06779, -44.97104, 
        -44.85891, -44.7299, -44.59463, -44.45291, -44.30928, -44.16974, 
        -44.04333, -43.92299, -43.80779, -43.69636, -43.59982, -43.52857, 
        -43.47218, -43.42556, -43.38536, -43.34841, -43.31365, -43.28537, 
        -43.25949, -43.23965, -43.22555, -43.2129, -43.20171, -43.19613, 
        -43.19431, -43.19429, -43.19568, -43.19547, -43.19659, -43.1973, 
        -43.19475, -43.19094, -43.18238, -43.17179, -43.16153, -43.15572, 
        -43.13955, -43.11501, -43.08347, -43.04594, -43.01139, -42.9748, 
        -42.93963, -42.90631, -42.87296, -42.84, -42.80901, -42.77283, 
        -42.73291, -42.69092, -42.65072, -42.61235, -42.58066, -42.55331, 
        -42.53103, -42.51543, -42.50344, -42.49136, -42.48185, -42.47925, 
        -42.48023, -42.48278, -42.48704, -42.48896, -42.48876, -42.48602, 
        -42.48126, -42.4761, -42.46843, -42.45623, -42.44526, -42.43637, 
        -42.42786, -42.42247, -42.42102, -42.42141, -42.42734, -42.43161, 
        -42.43801, -42.44281, -42.44635, -42.44382, -42.44967, -42.45412, 
        -42.45861, -42.46505, -42.47606, -42.48469, -42.49475, -42.50602, 
        -42.51892, -42.5337, -42.55038, -42.57062, -42.59247, -42.61478, 
        -42.63623, -42.65689, -42.67391, -42.68742, -42.69691, -42.70401, 
        -42.71048, -42.71539, -42.72174, -42.72896, -42.73829, -42.74844, 
        -42.75992, -42.77192, -42.78493, -42.79827, -42.81297, -42.82864, 
        -42.84541, -42.86203, -42.87983, -42.89747, -42.91433, -42.92963, 
        -42.94381, -42.95643, -42.96785, -42.97683, -42.98373, -42.98789, 
        -42.98917, -42.98597, -42.97826, -42.96591, -42.9497, -42.929, 
        -42.9073, -42.88442, -42.86201, -42.84062, -42.8208, -42.801, 
        -42.78065, -42.75771, -42.73148, -42.70456, -42.67105, -42.63684, 
        -42.60426, -42.57613, -42.5484, -42.52881, -42.51223, -42.50101, 
        -42.49176, -42.48096, -42.46617, -42.45082, -42.44028, -42.4371, 
        -42.43383, -42.43165, -42.42829, -42.41815, -42.43099, -42.46881, 
        -42.49897, -42.54567, -42.60728, -42.66835, -42.72636, -42.78427, 
        -42.84596, -42.90311, -42.96541, -43.0369, -43.11843, -43.21793, 
        -43.32723, -43.44724, -43.57624, -43.71231, -43.85564, -44.00559, 
        -44.16188, -44.32246, -44.48498, -44.64512, -44.79879, -44.94248, 
        -45.07333, -45.18896, -45.28844, -45.37286, -45.4448, -45.50527, 
        -45.55792, -45.60354, -45.6441, -45.67905, -45.70829, -45.73119, 
        -45.74827,
  -37.86591, -37.94178, -38.0158, -38.0859, -38.1493, -38.2058, -38.2584, 
        -38.30363, -38.34604, -38.38869, -38.4339, -38.47979, -38.52871, 
        -38.58253, -38.64017, -38.70256, -38.76832, -38.83735, -38.911, 
        -38.99002, -39.07246, -39.15758, -39.24718, -39.3464, -39.4544, 
        -39.56863, -39.69324, -39.8234, -39.95864, -40.09252, -40.22952, 
        -40.37028, -40.51955, -40.66709, -40.81227, -40.95981, -41.1042, 
        -41.24826, -41.39109, -41.53093, -41.66805, -41.7994, -41.9232, 
        -42.04015, -42.14831, -42.2477, -42.33915, -42.42404, -42.50437, 
        -42.5809, -42.65361, -42.7224, -42.78626, -42.84536, -42.89944, 
        -42.95007, -42.99938, -43.04878, -43.09956, -43.15176, -43.208, 
        -43.26751, -43.33106, -43.39902, -43.47103, -43.54567, -43.6226, 
        -43.69799, -43.77311, -43.84766, -43.92132, -43.99456, -44.06778, 
        -44.14124, -44.2158, -44.2909, -44.36621, -44.44355, -44.52146, 
        -44.59966, -44.67757, -44.75431, -44.82822, -44.89622, -44.95598, 
        -45.00491, -45.04053, -45.06132, -45.06797, -45.06188, -45.04731, 
        -45.02884, -45.00974, -44.99129, -44.97225, -44.95214, -44.92638, 
        -44.89158, -44.84449, -44.78217, -44.70284, -44.6065, -44.49508, 
        -44.37032, -44.23891, -44.10624, -43.97241, -43.84462, -43.72946, 
        -43.61938, -43.51474, -43.41153, -43.31855, -43.2382, -43.17698, 
        -43.12534, -43.08027, -43.03819, -42.99508, -42.96081, -42.92995, 
        -42.90355, -42.88349, -42.866, -42.85044, -42.83607, -42.826, 
        -42.81676, -42.81169, -42.80276, -42.80137, -42.80017, -42.79622, 
        -42.78899, -42.77917, -42.76722, -42.75524, -42.74626, -42.73671, 
        -42.71078, -42.67164, -42.63785, -42.60427, -42.56817, -42.53645, 
        -42.50418, -42.47263, -42.43695, -42.40363, -42.36929, -42.33696, 
        -42.29141, -42.25191, -42.21322, -42.18157, -42.15252, -42.13153, 
        -42.11241, -42.09654, -42.09015, -42.08981, -42.08958, -42.09256, 
        -42.09848, -42.10938, -42.11653, -42.11769, -42.11941, -42.11954, 
        -42.12057, -42.11916, -42.11296, -42.10376, -42.09415, -42.08753, 
        -42.084, -42.08438, -42.08417, -42.08883, -42.09382, -42.09937, 
        -42.10445, -42.10849, -42.10731, -42.11506, -42.11961, -42.1268, 
        -42.13611, -42.15249, -42.16511, -42.17851, -42.19612, -42.21442, 
        -42.23548, -42.25906, -42.28573, -42.31439, -42.34267, -42.3696, 
        -42.39503, -42.41714, -42.4348, -42.44881, -42.46071, -42.47114, 
        -42.48088, -42.4887, -42.4994, -42.5117, -42.52622, -42.5414, 
        -42.55702, -42.57333, -42.59003, -42.60741, -42.62527, -42.64394, 
        -42.66255, -42.68077, -42.69889, -42.71618, -42.73291, -42.74887, 
        -42.76382, -42.77783, -42.79041, -42.80137, -42.80967, -42.81514, 
        -42.81524, -42.80995, -42.79963, -42.78476, -42.76452, -42.743, 
        -42.7198, -42.69713, -42.67641, -42.65588, -42.63915, -42.62285, 
        -42.60562, -42.58566, -42.56672, -42.53961, -42.51086, -42.48502, 
        -42.46335, -42.44124, -42.4271, -42.41774, -42.41164, -42.40583, 
        -42.40091, -42.39209, -42.38169, -42.37243, -42.36629, -42.36399, 
        -42.36245, -42.35149, -42.34484, -42.38548, -42.43423, -42.47504, 
        -42.52279, -42.58342, -42.6476, -42.71389, -42.77511, -42.83641, 
        -42.90099, -42.97283, -43.05546, -43.15055, -43.25792, -43.37648, 
        -43.50309, -43.63717, -43.77534, -43.91721, -44.06227, -44.20992, 
        -44.3585, -44.50536, -44.64747, -44.78122, -44.90399, -45.01454, 
        -45.11208, -45.19605, -45.26899, -45.3329, -45.38959, -45.43957, 
        -45.48478, -45.52544, -45.56125, -45.59024, -45.6125, -45.62803,
  -37.9226, -37.99601, -38.06715, -38.13454, -38.1952, -38.24823, 
        -38.29571, -38.33435, -38.36883, -38.4056, -38.44273, -38.48095, 
        -38.52364, -38.57071, -38.62259, -38.67831, -38.73818, -38.80209, 
        -38.87008, -38.94496, -39.02432, -39.10974, -39.20107, -39.30326, 
        -39.41425, -39.53463, -39.66336, -39.79406, -39.92761, -40.0611, 
        -40.19697, -40.33625, -40.48547, -40.64007, -40.78782, -40.93544, 
        -41.08191, -41.2262, -41.37001, -41.51143, -41.64894, -41.78004, 
        -41.9044, -42.02055, -42.12755, -42.22583, -42.31691, -42.402, 
        -42.48233, -42.55875, -42.6309, -42.69857, -42.76106, -42.81728, 
        -42.86946, -42.91733, -42.96393, -43.00986, -43.05707, -43.10627, 
        -43.15798, -43.21262, -43.27036, -43.33233, -43.39783, -43.46617, 
        -43.53645, -43.60635, -43.67509, -43.74384, -43.81007, -43.8764, 
        -43.94227, -44.00792, -44.07367, -44.13995, -44.20722, -44.27519, 
        -44.3435, -44.41153, -44.47918, -44.5457, -44.60889, -44.66591, 
        -44.71485, -44.75278, -44.77736, -44.78702, -44.78412, -44.76995, 
        -44.74749, -44.72216, -44.6978, -44.67451, -44.65217, -44.62844, 
        -44.59963, -44.56138, -44.51171, -44.44705, -44.36602, -44.26861, 
        -44.157, -44.03336, -43.90678, -43.77897, -43.6544, -43.53682, 
        -43.43033, -43.3301, -43.23652, -43.14629, -43.06178, -42.98539, 
        -42.9188, -42.86084, -42.80384, -42.75269, -42.70349, -42.66166, 
        -42.62208, -42.58735, -42.56128, -42.5413, -42.51774, -42.49347, 
        -42.47241, -42.45495, -42.44176, -42.42919, -42.42238, -42.41745, 
        -42.40839, -42.39797, -42.38965, -42.37772, -42.36631, -42.34948, 
        -42.33705, -42.31995, -42.27945, -42.24637, -42.21386, -42.1773, 
        -42.14578, -42.11455, -42.08126, -42.04478, -42.01182, -41.97616, 
        -41.9509, -41.90454, -41.86587, -41.83022, -41.80038, -41.77559, 
        -41.7533, -41.729, -41.71338, -41.70493, -41.70213, -41.70648, 
        -41.71476, -41.72464, -41.73857, -41.75128, -41.75625, -41.76258, 
        -41.7685, -41.77607, -41.78191, -41.78106, -41.77328, -41.76734, 
        -41.76139, -41.75924, -41.75891, -41.75891, -41.76289, -41.76874, 
        -41.77628, -41.7841, -41.79215, -41.79258, -41.80065, -41.80935, 
        -41.8197, -41.8311, -41.85061, -41.86612, -41.88283, -41.90216, 
        -41.92416, -41.94988, -41.97951, -42.01278, -42.04844, -42.08281, 
        -42.1174, -42.15017, -42.17831, -42.20184, -42.22017, -42.23807, 
        -42.25521, -42.27008, -42.28157, -42.29492, -42.30967, -42.32575, 
        -42.34341, -42.3621, -42.3811, -42.40036, -42.42023, -42.43962, 
        -42.4586, -42.47713, -42.49555, -42.51369, -42.53171, -42.54902, 
        -42.5664, -42.58383, -42.60107, -42.61766, -42.63156, -42.64429, 
        -42.65446, -42.6584, -42.65653, -42.64862, -42.63548, -42.61673, 
        -42.59631, -42.57436, -42.5527, -42.53315, -42.51491, -42.50163, 
        -42.48892, -42.47504, -42.46044, -42.4482, -42.42935, -42.40566, 
        -42.38581, -42.36999, -42.35318, -42.34369, -42.33899, -42.33656, 
        -42.33497, -42.33401, -42.32852, -42.32065, -42.31437, -42.31081, 
        -42.30951, -42.3111, -42.301, -42.32114, -42.37222, -42.41745, 
        -42.46537, -42.52071, -42.58403, -42.65062, -42.71733, -42.78442, 
        -42.85363, -42.92777, -43.01043, -43.10424, -43.20883, -43.32503, 
        -43.45033, -43.58215, -43.71769, -43.85426, -43.99068, -44.12637, 
        -44.26049, -44.39202, -44.51884, -44.63895, -44.75042, -44.85194, 
        -44.94301, -45.02502, -45.09789, -45.16334, -45.22281, -45.27805, 
        -45.32895, -45.37593, -45.41875, -45.45576, -45.48581, -45.50787, 
        -45.52222,
  -37.98428, -38.05616, -38.12391, -38.18875, -38.24704, -38.29667, 
        -38.33979, -38.37586, -38.40815, -38.43932, -38.46804, -38.49622, 
        -38.52976, -38.56887, -38.61292, -38.66103, -38.71355, -38.77131, 
        -38.83279, -38.90182, -38.97738, -39.06108, -39.15483, -39.26452, 
        -39.38483, -39.51039, -39.64078, -39.7728, -39.90544, -40.03925, 
        -40.17506, -40.31295, -40.45953, -40.61856, -40.77049, -40.91875, 
        -41.06799, -41.21614, -41.36134, -41.50316, -41.63997, -41.76956, 
        -41.89206, -42.0057, -42.10986, -42.20596, -42.29547, -42.37894, 
        -42.45866, -42.53459, -42.60592, -42.6723, -42.7333, -42.78903, 
        -42.83941, -42.8855, -42.92928, -42.97226, -43.016, -43.06122, 
        -43.10831, -43.15759, -43.20979, -43.26543, -43.32352, -43.38516, 
        -43.44815, -43.51155, -43.57473, -43.63755, -43.69868, -43.75893, 
        -43.818, -43.87627, -43.9338, -43.99142, -44.04929, -44.10822, 
        -44.16672, -44.22491, -44.28249, -44.33772, -44.39071, -44.43768, 
        -44.47727, -44.50562, -44.52106, -44.52369, -44.51495, -44.49551, 
        -44.46891, -44.43614, -44.41232, -44.38667, -44.36177, -44.33615, 
        -44.30459, -44.26426, -44.21213, -44.14377, -44.05972, -43.96128, 
        -43.84806, -43.72324, -43.59755, -43.47356, -43.35677, -43.24727, 
        -43.14837, -43.05436, -42.96815, -42.88476, -42.80527, -42.73325, 
        -42.66747, -42.60676, -42.55046, -42.49577, -42.44218, -42.39464, 
        -42.34692, -42.30255, -42.26667, -42.2301, -42.19895, -42.1733, 
        -42.14248, -42.11601, -42.09543, -42.07556, -42.05817, -42.05104, 
        -42.03485, -42.02547, -42.01717, -42.00748, -41.99667, -41.97726, 
        -41.95944, -41.94925, -41.90659, -41.87143, -41.83732, -41.80075, 
        -41.7682, -41.73719, -41.70355, -41.66952, -41.63612, -41.6016, 
        -41.57839, -41.54609, -41.5003, -41.46689, -41.44008, -41.41823, 
        -41.39674, -41.36989, -41.34993, -41.34661, -41.33759, -41.3437, 
        -41.35433, -41.36663, -41.38169, -41.39916, -41.40968, -41.41943, 
        -41.42757, -41.4411, -41.45378, -41.46022, -41.4591, -41.45517, 
        -41.45224, -41.45132, -41.45125, -41.45178, -41.45322, -41.46009, 
        -41.47005, -41.48349, -41.49356, -41.49656, -41.5069, -41.51805, 
        -41.52855, -41.53888, -41.55967, -41.57742, -41.59737, -41.61986, 
        -41.64571, -41.67441, -41.70937, -41.752, -41.79319, -41.8362, 
        -41.87766, -41.91896, -41.95521, -41.98583, -42.01065, -42.03659, 
        -42.06152, -42.08126, -42.09753, -42.11264, -42.12909, -42.1466, 
        -42.16515, -42.18552, -42.20647, -42.22808, -42.24956, -42.26957, 
        -42.28773, -42.30576, -42.32306, -42.3418, -42.36086, -42.3795, 
        -42.39833, -42.41842, -42.43908, -42.45985, -42.47943, -42.49693, 
        -42.51214, -42.52044, -42.52213, -42.51695, -42.50625, -42.48981, 
        -42.47216, -42.4534, -42.43397, -42.41724, -42.40113, -42.39037, 
        -42.38016, -42.36713, -42.35429, -42.34963, -42.33699, -42.32303, 
        -42.30883, -42.29592, -42.28305, -42.27623, -42.27544, -42.27629, 
        -42.27687, -42.27797, -42.27394, -42.26664, -42.26579, -42.26844, 
        -42.27137, -42.28528, -42.30139, -42.33379, -42.37558, -42.42302, 
        -42.47827, -42.53907, -42.6054, -42.67458, -42.74795, -42.82254, 
        -42.9022, -42.98703, -43.07989, -43.1834, -43.29603, -43.418, 
        -43.54645, -43.67875, -43.81195, -43.94302, -44.07017, -44.19294, 
        -44.3104, -44.42159, -44.5256, -44.62164, -44.71011, -44.79047, 
        -44.86427, -44.9338, -44.99948, -45.06127, -45.12094, -45.17779, 
        -45.23145, -45.28123, -45.32582, -45.36391, -45.39404, -45.41538, 
        -45.42796,
  -38.04875, -38.11844, -38.18586, -38.24889, -38.30456, -38.35236, 
        -38.3922, -38.4252, -38.45319, -38.47906, -38.50183, -38.51933, 
        -38.54094, -38.56984, -38.60736, -38.64823, -38.69596, -38.74685, 
        -38.80222, -38.86682, -38.93888, -39.02155, -39.11822, -39.23394, 
        -39.3595, -39.49015, -39.62387, -39.75633, -39.88885, -40.02223, 
        -40.16029, -40.29858, -40.4465, -40.60477, -40.76069, -40.91225, 
        -41.06416, -41.21497, -41.36201, -41.50225, -41.63747, -41.76546, 
        -41.8833, -41.99279, -42.09361, -42.18701, -42.27449, -42.35747, 
        -42.43591, -42.51059, -42.58043, -42.64492, -42.70422, -42.75799, 
        -42.80617, -42.85007, -42.89105, -42.93095, -42.97013, -43.01157, 
        -43.05432, -43.09895, -43.14611, -43.19607, -43.24863, -43.30335, 
        -43.35953, -43.41643, -43.47386, -43.53086, -43.58692, -43.64124, 
        -43.69393, -43.74524, -43.79469, -43.84259, -43.89151, -43.94088, 
        -43.98985, -44.03815, -44.08547, -44.13153, -44.17431, -44.21201, 
        -44.24262, -44.26281, -44.27157, -44.26854, -44.25546, -44.23294, 
        -44.20419, -44.17449, -44.14571, -44.11847, -44.09177, -44.06517, 
        -44.03166, -43.99037, -43.93838, -43.86964, -43.78385, -43.68417, 
        -43.57097, -43.44525, -43.3163, -43.19186, -43.08006, -42.97438, 
        -42.87864, -42.78759, -42.70293, -42.62254, -42.54105, -42.47444, 
        -42.40583, -42.34887, -42.29266, -42.23997, -42.18317, -42.12801, 
        -42.07917, -42.03259, -41.98708, -41.94231, -41.89977, -41.8698, 
        -41.8359, -41.80124, -41.76733, -41.74145, -41.72145, -41.70835, 
        -41.68705, -41.67824, -41.66993, -41.65754, -41.64545, -41.6268, 
        -41.60741, -41.60082, -41.56008, -41.51923, -41.48349, -41.44559, 
        -41.41282, -41.38021, -41.3454, -41.31001, -41.27915, -41.24628, 
        -41.21949, -41.20211, -41.1607, -41.13064, -41.1053, -41.08247, 
        -41.06153, -41.03126, -41.0108, -41.00515, -40.99929, -41.00272, 
        -41.01073, -41.0219, -41.03999, -41.06296, -41.07681, -41.08832, 
        -41.09995, -41.11809, -41.13457, -41.14717, -41.15431, -41.15919, 
        -41.15892, -41.15471, -41.15531, -41.15668, -41.15755, -41.16589, 
        -41.17825, -41.18921, -41.20003, -41.20534, -41.21769, -41.23277, 
        -41.24619, -41.25677, -41.28056, -41.30111, -41.32556, -41.35147, 
        -41.37935, -41.41488, -41.46036, -41.50401, -41.55286, -41.60205, 
        -41.64914, -41.69766, -41.7424, -41.78144, -41.81463, -41.85257, 
        -41.88435, -41.90838, -41.92862, -41.94849, -41.96794, -41.98754, 
        -42.00794, -42.02898, -42.0504, -42.07304, -42.09548, -42.11684, 
        -42.1362, -42.15378, -42.16993, -42.18799, -42.20739, -42.22781, 
        -42.2484, -42.27144, -42.29497, -42.31943, -42.34364, -42.36744, 
        -42.3885, -42.40092, -42.40616, -42.40425, -42.39646, -42.38269, 
        -42.36825, -42.35268, -42.33756, -42.32221, -42.304, -42.2923, 
        -42.28022, -42.25853, -42.24925, -42.25141, -42.25433, -42.24628, 
        -42.24078, -42.23573, -42.22952, -42.2292, -42.23227, -42.23577, 
        -42.23634, -42.24018, -42.2374, -42.23436, -42.23699, -42.24848, 
        -42.26348, -42.28667, -42.31558, -42.3517, -42.3979, -42.44731, 
        -42.50746, -42.57439, -42.64698, -42.72452, -42.80759, -42.89224, 
        -42.98048, -43.07603, -43.17769, -43.28778, -43.4056, -43.52884, 
        -43.65726, -43.78693, -43.91434, -44.03653, -44.15174, -44.25866, 
        -44.35666, -44.44569, -44.52566, -44.59807, -44.66456, -44.72662, 
        -44.78727, -44.84843, -44.91109, -44.97395, -45.03649, -45.09655, 
        -45.15343, -45.20506, -45.2504, -45.28735, -45.31537, -45.33414, 
        -45.34356,
  -38.12023, -38.18838, -38.25416, -38.31519, -38.36842, -38.41344, 
        -38.44923, -38.47869, -38.50291, -38.52262, -38.53898, -38.55344, 
        -38.56595, -38.58329, -38.60758, -38.63994, -38.67955, -38.72562, 
        -38.77685, -38.83866, -38.90783, -38.98915, -39.0872, -39.20357, 
        -39.33593, -39.47214, -39.61131, -39.74944, -39.884, -40.01876, 
        -40.15381, -40.29448, -40.44415, -40.60386, -40.76081, -40.91617, 
        -41.07095, -41.22212, -41.36821, -41.50758, -41.64004, -41.76435, 
        -41.87934, -41.98449, -42.0813, -42.17151, -42.25652, -42.3373, 
        -42.41419, -42.48684, -42.55446, -42.61667, -42.67243, -42.72347, 
        -42.76904, -42.81002, -42.84788, -42.88407, -42.92054, -42.95746, 
        -42.99587, -43.03595, -43.07827, -43.12287, -43.16942, -43.21776, 
        -43.26733, -43.31832, -43.37023, -43.42122, -43.47193, -43.52119, 
        -43.56811, -43.61188, -43.65359, -43.69415, -43.73425, -43.77433, 
        -43.81354, -43.8522, -43.88932, -43.92529, -43.9584, -43.98711, 
        -44.00932, -44.02286, -44.02601, -44.01857, -44.00213, -43.97902, 
        -43.95086, -43.91972, -43.89059, -43.86425, -43.83745, -43.81013, 
        -43.77756, -43.73712, -43.68538, -43.61651, -43.53239, -43.43089, 
        -43.31836, -43.19435, -43.06495, -42.93539, -42.82, -42.71374, 
        -42.61556, -42.52367, -42.43925, -42.36273, -42.28242, -42.21801, 
        -42.15618, -42.09545, -42.03933, -41.98653, -41.93001, -41.87848, 
        -41.82591, -41.76248, -41.70653, -41.65652, -41.61275, -41.57374, 
        -41.53067, -41.49347, -41.45704, -41.42878, -41.40683, -41.38718, 
        -41.36318, -41.35274, -41.34022, -41.32751, -41.31513, -41.29238, 
        -41.27091, -41.25643, -41.23483, -41.18602, -41.15047, -41.11167, 
        -41.0737, -41.03833, -41.00342, -40.96748, -40.93687, -40.90454, 
        -40.8779, -40.86623, -40.84206, -40.80691, -40.78478, -40.76237, 
        -40.73723, -40.71032, -40.69195, -40.68373, -40.68349, -40.68037, 
        -40.69157, -40.70012, -40.71409, -40.7406, -40.75614, -40.7704, 
        -40.78327, -40.80112, -40.82204, -40.8417, -40.85609, -40.86783, 
        -40.87223, -40.87392, -40.87876, -40.88165, -40.8842, -40.9013, 
        -40.91332, -40.92103, -40.92851, -40.93766, -40.94823, -40.97056, 
        -40.98674, -40.99663, -41.02166, -41.04368, -41.06845, -41.09489, 
        -41.12362, -41.1563, -41.21925, -41.27158, -41.3297, -41.38537, 
        -41.4384, -41.49393, -41.55003, -41.59578, -41.64214, -41.68894, 
        -41.72711, -41.75715, -41.78159, -41.80591, -41.82832, -41.8506, 
        -41.87259, -41.89454, -41.91684, -41.93932, -41.96286, -41.98561, 
        -42.00603, -42.02364, -42.04027, -42.05758, -42.07649, -42.09759, 
        -42.11988, -42.14507, -42.17174, -42.1991, -42.22821, -42.25695, 
        -42.28431, -42.30114, -42.31036, -42.31257, -42.30867, -42.29935, 
        -42.28986, -42.27972, -42.27028, -42.26143, -42.23844, -42.22641, 
        -42.22002, -42.2015, -42.18756, -42.19125, -42.19481, -42.18864, 
        -42.18517, -42.1885, -42.1937, -42.19818, -42.20221, -42.20587, 
        -42.20422, -42.20372, -42.19318, -42.19072, -42.1995, -42.22948, 
        -42.25964, -42.29092, -42.33087, -42.37677, -42.4306, -42.48679, 
        -42.55254, -42.62962, -42.71182, -42.80129, -42.89494, -42.98963, 
        -43.08674, -43.18799, -43.29515, -43.40883, -43.52787, -43.65148, 
        -43.77659, -43.90095, -44.02032, -44.13177, -44.233, -44.32287, 
        -44.40059, -44.46694, -44.52418, -44.57443, -44.62106, -44.66919, 
        -44.72028, -44.77721, -44.83971, -44.90559, -44.97186, -45.03646, 
        -45.09361, -45.14465, -45.18774, -45.22086, -45.24406, -45.2576, 
        -45.26191,
  -38.19852, -38.26371, -38.32715, -38.38531, -38.43544, -38.47731, 
        -38.51061, -38.53619, -38.55588, -38.57085, -38.58131, -38.59029, 
        -38.59644, -38.60129, -38.61674, -38.64068, -38.67016, -38.70934, 
        -38.75589, -38.81719, -38.8871, -38.97131, -39.07147, -39.18849, 
        -39.32282, -39.46185, -39.60486, -39.74685, -39.88692, -40.02374, 
        -40.16214, -40.3069, -40.45781, -40.61339, -40.77116, -40.93109, 
        -41.08733, -41.24006, -41.38382, -41.52121, -41.64926, -41.76902, 
        -41.87928, -41.98043, -42.07355, -42.16027, -42.24247, -42.32003, 
        -42.39468, -42.46474, -42.52945, -42.58854, -42.64198, -42.68948, 
        -42.73141, -42.76842, -42.80239, -42.83405, -42.86564, -42.89812, 
        -42.93147, -42.96645, -43.0036, -43.04145, -43.08243, -43.12496, 
        -43.16853, -43.21435, -43.2612, -43.30861, -43.35538, -43.39893, 
        -43.4403, -43.47788, -43.51198, -43.54432, -43.57568, -43.60671, 
        -43.63647, -43.66561, -43.69168, -43.71859, -43.74231, -43.7626, 
        -43.77765, -43.78493, -43.78364, -43.77383, -43.75593, -43.73164, 
        -43.70323, -43.67369, -43.64401, -43.61676, -43.59046, -43.56307, 
        -43.53145, -43.49164, -43.44129, -43.37451, -43.29188, -43.19412, 
        -43.08368, -42.96333, -42.83801, -42.71324, -42.58818, -42.47115, 
        -42.36597, -42.26995, -42.18581, -42.11217, -42.0388, -41.97355, 
        -41.9077, -41.84437, -41.78444, -41.73199, -41.674, -41.62442, 
        -41.5746, -41.52031, -41.45972, -41.39723, -41.34242, -41.29456, 
        -41.24663, -41.20324, -41.1678, -41.13604, -41.11274, -41.09018, 
        -41.06834, -41.05285, -41.03751, -41.02101, -41.00135, -40.98098, 
        -40.96082, -40.94167, -40.93144, -40.87774, -40.83256, -40.79348, 
        -40.75048, -40.71152, -40.67481, -40.6404, -40.61111, -40.58141, 
        -40.55651, -40.54644, -40.53243, -40.49525, -40.4743, -40.44981, 
        -40.41962, -40.39845, -40.38192, -40.37379, -40.37409, -40.37531, 
        -40.37365, -40.38692, -40.40404, -40.4309, -40.45576, -40.47395, 
        -40.48611, -40.50143, -40.52236, -40.5485, -40.57127, -40.58579, 
        -40.60094, -40.60624, -40.61576, -40.62412, -40.62893, -40.65232, 
        -40.66659, -40.6777, -40.67799, -40.68954, -40.70225, -40.72622, 
        -40.74323, -40.75534, -40.77404, -40.79353, -40.81408, -40.83108, 
        -40.85825, -40.8997, -40.97317, -41.05046, -41.11919, -41.18125, 
        -41.23927, -41.30921, -41.3801, -41.4402, -41.49386, -41.54639, 
        -41.59053, -41.62716, -41.65721, -41.68377, -41.70958, -41.73385, 
        -41.758, -41.78082, -41.80302, -41.82633, -41.8503, -41.87426, 
        -41.89582, -41.91483, -41.93092, -41.94896, -41.96604, -41.9868, 
        -42.00928, -42.03737, -42.06815, -42.10103, -42.13474, -42.16802, 
        -42.2019, -42.22319, -42.23607, -42.24221, -42.24311, -42.23939, 
        -42.23647, -42.23261, -42.22991, -42.22673, -42.2149, -42.2128, 
        -42.20934, -42.20274, -42.19671, -42.20225, -42.19822, -42.18276, 
        -42.1731, -42.17429, -42.17257, -42.18257, -42.18852, -42.19077, 
        -42.18845, -42.17869, -42.17289, -42.17784, -42.19178, -42.22181, 
        -42.26933, -42.3124, -42.35927, -42.4171, -42.48126, -42.54766, 
        -42.62709, -42.71335, -42.80524, -42.90479, -43.00727, -43.1087, 
        -43.21128, -43.31626, -43.42468, -43.53846, -43.6555, -43.77467, 
        -43.89452, -44.01107, -44.12088, -44.221, -44.30796, -44.38012, 
        -44.43906, -44.48517, -44.52166, -44.55295, -44.5846, -44.62228, 
        -44.66791, -44.72271, -44.7878, -44.8577, -44.92614, -44.99151, 
        -45.04835, -45.09509, -45.13201, -45.15763, -45.17314, -45.17902, 
        -45.17695,
  -38.28151, -38.34485, -38.4047, -38.459, -38.50523, -38.54327, 
        -38.57243, -38.59371, -38.60891, -38.6186, -38.62331, -38.62468, 
        -38.62346, -38.62354, -38.63218, -38.64795, -38.66988, -38.70371, 
        -38.74792, -38.8061, -38.87659, -38.9631, -39.0672, -39.18784, 
        -39.32235, -39.46386, -39.60754, -39.75202, -39.89528, -40.03694, 
        -40.18008, -40.32727, -40.48065, -40.63963, -40.80097, -40.95975, 
        -41.11773, -41.26723, -41.40778, -41.54095, -41.66463, -41.77863, 
        -41.88466, -41.98196, -42.07158, -42.15518, -42.23436, -42.31033, 
        -42.38214, -42.44927, -42.51057, -42.56582, -42.61504, -42.65778, 
        -42.69497, -42.72722, -42.75611, -42.78127, -42.8067, -42.83291, 
        -42.86025, -42.88916, -42.92019, -42.95311, -42.98842, -43.02555, 
        -43.0646, -43.1054, -43.14896, -43.19239, -43.23438, -43.27347, 
        -43.30886, -43.34044, -43.36687, -43.39169, -43.41491, -43.4371, 
        -43.45801, -43.47775, -43.49668, -43.5146, -43.53002, -43.54266, 
        -43.55069, -43.55241, -43.54704, -43.53465, -43.51534, -43.49012, 
        -43.46132, -43.43092, -43.39997, -43.37161, -43.34415, -43.31621, 
        -43.28525, -43.24705, -43.19964, -43.1376, -43.05915, -42.96564, 
        -42.86025, -42.74403, -42.62487, -42.50191, -42.38042, -42.26103, 
        -42.14621, -42.04234, -41.96136, -41.88607, -41.80811, -41.73727, 
        -41.66201, -41.59423, -41.53306, -41.48058, -41.4273, -41.37612, 
        -41.3243, -41.2724, -41.21658, -41.15612, -41.09256, -41.03839, 
        -40.98726, -40.93647, -40.89456, -40.86109, -40.83626, -40.80944, 
        -40.78573, -40.77346, -40.75608, -40.73654, -40.71768, -40.70191, 
        -40.6846, -40.66801, -40.64798, -40.60602, -40.55231, -40.5071, 
        -40.46314, -40.41853, -40.37152, -40.33521, -40.30546, -40.28088, 
        -40.261, -40.24361, -40.22513, -40.20392, -40.18166, -40.14571, 
        -40.11454, -40.09052, -40.07577, -40.0657, -40.06369, -40.06458, 
        -40.06742, -40.08137, -40.10342, -40.13103, -40.16348, -40.19001, 
        -40.20413, -40.21639, -40.24663, -40.27543, -40.30273, -40.31821, 
        -40.34251, -40.35778, -40.36924, -40.38375, -40.40394, -40.42463, 
        -40.43632, -40.4496, -40.46342, -40.46511, -40.48, -40.50484, 
        -40.52632, -40.52905, -40.52975, -40.55586, -40.56926, -40.58195, 
        -40.60442, -40.66437, -40.76293, -40.851, -40.92971, -41.00414, 
        -41.07933, -41.16388, -41.24052, -41.30725, -41.36461, -41.42237, 
        -41.47254, -41.51625, -41.55141, -41.58206, -41.61026, -41.63821, 
        -41.66289, -41.68624, -41.70942, -41.734, -41.75963, -41.78522, 
        -41.80787, -41.82819, -41.84504, -41.86359, -41.88193, -41.89971, 
        -41.92085, -41.95035, -41.98242, -42.02557, -42.06423, -42.10301, 
        -42.13972, -42.16417, -42.18066, -42.19111, -42.19751, -42.20017, 
        -42.20384, -42.20681, -42.21132, -42.21562, -42.21098, -42.21457, 
        -42.21719, -42.21736, -42.2134, -42.21886, -42.21252, -42.20122, 
        -42.18854, -42.1884, -42.18735, -42.18885, -42.19381, -42.197, 
        -42.19764, -42.19952, -42.20302, -42.21465, -42.23274, -42.25685, 
        -42.29778, -42.34774, -42.40475, -42.47215, -42.54865, -42.62619, 
        -42.71798, -42.81789, -42.92201, -43.02744, -43.13586, -43.2412, 
        -43.34548, -43.44972, -43.55556, -43.66406, -43.77597, -43.88866, 
        -44.00038, -44.10794, -44.20749, -44.2957, -44.36934, -44.42616, 
        -44.46852, -44.4974, -44.51809, -44.5361, -44.55819, -44.5895, 
        -44.63324, -44.69014, -44.75695, -44.82821, -44.89742, -44.95938, 
        -45.01163, -45.05098, -45.07837, -45.09396, -45.0992, -45.09613, 
        -45.08659,
  -38.36907, -38.4283, -38.48385, -38.53324, -38.57458, -38.60713, 
        -38.63036, -38.64726, -38.65756, -38.66218, -38.66227, -38.65821, 
        -38.65186, -38.64722, -38.64846, -38.65763, -38.67466, -38.70369, 
        -38.74613, -38.80465, -38.87868, -38.96701, -39.07393, -39.19897, 
        -39.33404, -39.47656, -39.62297, -39.77052, -39.91663, -40.06225, 
        -40.20963, -40.35937, -40.51552, -40.6775, -40.83987, -41.00038, 
        -41.15452, -41.30143, -41.43944, -41.56776, -41.68715, -41.79771, 
        -41.89965, -41.99329, -42.07978, -42.16055, -42.23704, -42.3103, 
        -42.37922, -42.44283, -42.50039, -42.55122, -42.59444, -42.63166, 
        -42.66295, -42.68886, -42.71046, -42.72945, -42.74771, -42.76651, 
        -42.78617, -42.80725, -42.83076, -42.85672, -42.88578, -42.91726, 
        -42.95152, -42.98909, -43.02696, -43.06631, -43.10428, -43.13988, 
        -43.1708, -43.19718, -43.21964, -43.23884, -43.2556, -43.27085, 
        -43.28436, -43.29644, -43.30738, -43.31728, -43.32486, -43.33038, 
        -43.33155, -43.32794, -43.31711, -43.30198, -43.28061, -43.25376, 
        -43.22383, -43.19232, -43.16073, -43.13023, -43.10089, -43.07141, 
        -43.0399, -43.00326, -42.95844, -42.89935, -42.82635, -42.73872, 
        -42.63932, -42.52921, -42.41672, -42.29971, -42.18285, -42.0662, 
        -41.96215, -41.86439, -41.77755, -41.69276, -41.60329, -41.5239, 
        -41.44325, -41.36398, -41.30109, -41.24731, -41.19022, -41.13425, 
        -41.08138, -41.02847, -40.97268, -40.92175, -40.86494, -40.80596, 
        -40.74322, -40.69405, -40.6433, -40.60138, -40.57603, -40.55043, 
        -40.52468, -40.51447, -40.49181, -40.47565, -40.46276, -40.46009, 
        -40.45069, -40.41452, -40.37185, -40.33522, -40.27612, -40.2217, 
        -40.16677, -40.12589, -40.08746, -40.05064, -40.02433, -40.00396, 
        -39.97812, -39.95585, -39.94259, -39.91795, -39.89526, -39.85999, 
        -39.82813, -39.79266, -39.77192, -39.75751, -39.7534, -39.75286, 
        -39.76246, -39.77311, -39.80595, -39.84871, -39.88654, -39.91973, 
        -39.93586, -39.94606, -39.96412, -40.00364, -40.04579, -40.07283, 
        -40.09975, -40.1266, -40.15719, -40.18407, -40.20406, -40.21565, 
        -40.22846, -40.23784, -40.25833, -40.26949, -40.29187, -40.32116, 
        -40.33267, -40.33406, -40.33842, -40.34765, -40.36724, -40.38236, 
        -40.42514, -40.4991, -40.5942, -40.66837, -40.76046, -40.8632, 
        -40.9629, -41.0503, -41.12425, -41.19227, -41.25388, -41.31829, 
        -41.37409, -41.4223, -41.4631, -41.49797, -41.53031, -41.55895, 
        -41.58509, -41.60981, -41.63522, -41.66069, -41.68734, -41.71441, 
        -41.73997, -41.76201, -41.7803, -41.79992, -41.81946, -41.8431, 
        -41.8681, -41.8985, -41.92892, -41.97144, -42.01485, -42.0554, 
        -42.09359, -42.12063, -42.14112, -42.15636, -42.16861, -42.17794, 
        -42.18878, -42.20027, -42.21239, -42.22442, -42.22631, -42.23579, 
        -42.24342, -42.24775, -42.24827, -42.25389, -42.24729, -42.23651, 
        -42.22738, -42.22153, -42.21793, -42.21814, -42.21974, -42.22292, 
        -42.22624, -42.23376, -42.24145, -42.2557, -42.27761, -42.30878, 
        -42.3473, -42.39977, -42.46573, -42.54365, -42.63151, -42.72268, 
        -42.82736, -42.93732, -43.04919, -43.15994, -43.27065, -43.37578, 
        -43.4777, -43.57745, -43.67752, -43.77969, -43.88327, -43.98729, 
        -44.08941, -44.18659, -44.27515, -44.35155, -44.4128, -44.45745, 
        -44.48695, -44.50467, -44.51574, -44.52703, -44.5451, -44.57501, 
        -44.61811, -44.67541, -44.74116, -44.81035, -44.87516, -44.93088, 
        -44.97411, -45.0034, -45.01928, -45.02353, -45.01822, -45.00602, 
        -44.98872,
  -38.45714, -38.51036, -38.56032, -38.60364, -38.63839, -38.66511, 
        -38.68376, -38.69545, -38.70126, -38.70111, -38.69639, -38.68823, 
        -38.67777, -38.67005, -38.66412, -38.66673, -38.67956, -38.70841, 
        -38.75275, -38.81005, -38.88649, -38.98029, -39.09107, -39.217, 
        -39.3531, -39.49769, -39.64697, -39.7977, -39.94864, -40.09883, 
        -40.24896, -40.40273, -40.562, -40.72595, -40.88931, -41.04895, 
        -41.20208, -41.34638, -41.48086, -41.60592, -41.72107, -41.82752, 
        -41.92572, -42.01624, -42.10003, -42.17844, -42.2517, -42.32246, 
        -42.38838, -42.4484, -42.50158, -42.5472, -42.58556, -42.61622, 
        -42.64017, -42.65775, -42.67071, -42.68106, -42.69059, -42.69999, 
        -42.71032, -42.72232, -42.73709, -42.75432, -42.77647, -42.80259, 
        -42.83286, -42.86633, -42.90186, -42.93738, -42.97139, -43.00299, 
        -43.0304, -43.05339, -43.07202, -43.08691, -43.09912, -43.10902, 
        -43.11647, -43.12217, -43.12561, -43.12858, -43.12932, -43.12776, 
        -43.12305, -43.11419, -43.10039, -43.08131, -43.0574, -43.02844, 
        -42.99614, -42.9621, -42.92726, -42.89272, -42.85903, -42.82609, 
        -42.7926, -42.7561, -42.71342, -42.65853, -42.59057, -42.50991, 
        -42.41758, -42.31222, -42.20719, -42.10062, -41.99192, -41.88436, 
        -41.78485, -41.68545, -41.59266, -41.50267, -41.41513, -41.33468, 
        -41.25292, -41.16964, -41.10286, -41.04026, -40.97136, -40.91156, 
        -40.8537, -40.80041, -40.74546, -40.69471, -40.64075, -40.58121, 
        -40.51309, -40.46124, -40.41363, -40.36367, -40.3344, -40.30259, 
        -40.27797, -40.2609, -40.24446, -40.23349, -40.22976, -40.23218, 
        -40.21806, -40.16574, -40.11213, -40.0772, -40.0098, -39.94457, 
        -39.891, -39.84053, -39.80484, -39.77646, -39.75663, -39.73903, 
        -39.72264, -39.69323, -39.67714, -39.63353, -39.60147, -39.57663, 
        -39.5463, -39.52235, -39.50449, -39.478, -39.46766, -39.46465, 
        -39.47521, -39.49567, -39.52369, -39.5575, -39.59665, -39.64737, 
        -39.68111, -39.68555, -39.70638, -39.74931, -39.79415, -39.8237, 
        -39.85781, -39.9001, -39.94575, -39.99002, -40.02374, -40.05135, 
        -40.07102, -40.08708, -40.09601, -40.11452, -40.13937, -40.17257, 
        -40.187, -40.18391, -40.18233, -40.18229, -40.20066, -40.24009, 
        -40.30696, -40.37648, -40.447, -40.54912, -40.66323, -40.77488, 
        -40.87182, -40.94648, -41.01952, -41.09995, -41.16969, -41.2356, 
        -41.29355, -41.34501, -41.39086, -41.43071, -41.46634, -41.49724, 
        -41.52497, -41.5516, -41.57755, -41.60291, -41.63179, -41.66047, 
        -41.68776, -41.71226, -41.73344, -41.7554, -41.77831, -41.80309, 
        -41.83016, -41.86118, -41.89746, -41.93997, -41.98286, -42.02398, 
        -42.06153, -42.09172, -42.11687, -42.1381, -42.15706, -42.1744, 
        -42.19289, -42.21279, -42.23354, -42.25351, -42.265, -42.27982, 
        -42.29134, -42.29854, -42.30002, -42.30223, -42.2941, -42.283, 
        -42.27266, -42.26565, -42.26165, -42.26027, -42.26031, -42.26184, 
        -42.26447, -42.27312, -42.28325, -42.30007, -42.32506, -42.35998, 
        -42.40423, -42.46475, -42.54007, -42.62745, -42.72818, -42.83274, 
        -42.94843, -43.06665, -43.1834, -43.29563, -43.40405, -43.50478, 
        -43.60012, -43.69189, -43.78278, -43.87526, -43.96871, -44.06246, 
        -44.15411, -44.24013, -44.31824, -44.38448, -44.43569, -44.47145, 
        -44.49343, -44.50542, -44.51329, -44.52364, -44.54329, -44.57506, 
        -44.61872, -44.67418, -44.73671, -44.79869, -44.85429, -44.89911, 
        -44.93019, -44.94692, -44.95037, -44.94308, -44.92804, -44.90754, 
        -44.88355,
  -38.54168, -38.59054, -38.63404, -38.67014, -38.69781, -38.71737, 
        -38.73037, -38.7364, -38.73672, -38.7319, -38.7219, -38.70993, 
        -38.69651, -38.68527, -38.67628, -38.67683, -38.68821, -38.71629, 
        -38.76001, -38.82021, -38.90009, -38.99596, -39.10992, -39.23714, 
        -39.37467, -39.51962, -39.67106, -39.82541, -39.98026, -40.13509, 
        -40.29108, -40.44993, -40.61284, -40.77719, -40.94104, -41.10053, 
        -41.25294, -41.39658, -41.52987, -41.65303, -41.76588, -41.86831, 
        -41.96368, -42.05164, -42.13322, -42.21001, -42.28219, -42.35089, 
        -42.41371, -42.46991, -42.51798, -42.55785, -42.58975, -42.6129, 
        -42.62817, -42.63605, -42.63907, -42.63805, -42.63658, -42.63489, 
        -42.63404, -42.63523, -42.63962, -42.64859, -42.66325, -42.683, 
        -42.70852, -42.73761, -42.76966, -42.80159, -42.83319, -42.8617, 
        -42.88706, -42.90849, -42.9244, -42.93739, -42.94718, -42.95384, 
        -42.95714, -42.95834, -42.95797, -42.95502, -42.95012, -42.94266, 
        -42.93221, -42.91839, -42.90005, -42.87814, -42.85072, -42.81854, 
        -42.7827, -42.74467, -42.70398, -42.66398, -42.62532, -42.58802, 
        -42.5515, -42.51321, -42.47205, -42.42087, -42.3584, -42.28362, 
        -42.19763, -42.09887, -42.00121, -41.90129, -41.80076, -41.70033, 
        -41.60142, -41.5013, -41.40235, -41.30904, -41.22203, -41.14087, 
        -41.0541, -40.9712, -40.89588, -40.81766, -40.73938, -40.68162, 
        -40.63193, -40.57782, -40.53123, -40.48272, -40.43217, -40.37164, 
        -40.31385, -40.25002, -40.19772, -40.14444, -40.1035, -40.06981, 
        -40.04029, -40.0192, -40.00812, -40.01479, -40.02987, -40.03602, 
        -40.01564, -39.96945, -39.90752, -39.86139, -39.76986, -39.69176, 
        -39.63768, -39.58383, -39.54655, -39.51562, -39.49187, -39.4919, 
        -39.47722, -39.44377, -39.43206, -39.39288, -39.3474, -39.30896, 
        -39.27527, -39.26471, -39.23866, -39.22829, -39.21194, -39.20751, 
        -39.22206, -39.23862, -39.26505, -39.30103, -39.34546, -39.39925, 
        -39.43228, -39.44458, -39.47821, -39.52502, -39.56985, -39.60103, 
        -39.64392, -39.69738, -39.75064, -39.80641, -39.85287, -39.89294, 
        -39.9265, -39.9529, -39.97648, -40.00351, -40.02532, -40.0415, 
        -40.05306, -40.0588, -40.06947, -40.0784, -40.10042, -40.15268, 
        -40.23513, -40.30384, -40.36407, -40.464, -40.59719, -40.71058, 
        -40.794, -40.86467, -40.94197, -41.02692, -41.09948, -41.16489, 
        -41.22468, -41.27998, -41.32948, -41.37369, -41.4125, -41.44486, 
        -41.47449, -41.50191, -41.52871, -41.55745, -41.5879, -41.61868, 
        -41.64832, -41.67527, -41.69796, -41.7233, -41.74942, -41.77746, 
        -41.80654, -41.84048, -41.87773, -41.91839, -41.96165, -42.00168, 
        -42.04168, -42.07579, -42.10654, -42.13409, -42.1601, -42.18523, 
        -42.21166, -42.23975, -42.26902, -42.29622, -42.31527, -42.33537, 
        -42.35113, -42.36079, -42.36355, -42.36618, -42.35985, -42.34998, 
        -42.34095, -42.33392, -42.33022, -42.32737, -42.32582, -42.32602, 
        -42.32778, -42.33632, -42.34771, -42.3666, -42.3954, -42.43525, 
        -42.48544, -42.55351, -42.63727, -42.73449, -42.84276, -42.95719, 
        -43.07856, -43.20005, -43.31672, -43.42556, -43.5275, -43.61959, 
        -43.70493, -43.78575, -43.86407, -43.94444, -44.02617, -44.10866, 
        -44.18902, -44.26502, -44.33315, -44.39072, -44.43521, -44.46646, 
        -44.48621, -44.4986, -44.50904, -44.52353, -44.54792, -44.58318, 
        -44.62735, -44.68032, -44.73593, -44.78814, -44.83158, -44.86267, 
        -44.87943, -44.88182, -44.87301, -44.8555, -44.8319, -44.80486, 
        -44.77633,
  -38.62148, -38.66398, -38.7004, -38.72926, -38.74922, -38.76077, 
        -38.76657, -38.76664, -38.76168, -38.75245, -38.7398, -38.72516, 
        -38.7104, -38.696, -38.68644, -38.68714, -38.69659, -38.72553, 
        -38.76865, -38.83089, -38.91187, -39.0094, -39.12405, -39.25212, 
        -39.3897, -39.53564, -39.68793, -39.84466, -40.00428, -40.16486, 
        -40.32714, -40.49142, -40.65794, -40.82497, -40.99003, -41.14999, 
        -41.30373, -41.44829, -41.58252, -41.70651, -41.81914, -41.92178, 
        -42.01564, -42.10193, -42.18216, -42.25759, -42.32874, -42.39513, 
        -42.45477, -42.50661, -42.54953, -42.58213, -42.60644, -42.621, 
        -42.62651, -42.62447, -42.6163, -42.60448, -42.59031, -42.57582, 
        -42.56219, -42.55079, -42.54364, -42.54256, -42.54843, -42.56153, 
        -42.58105, -42.60575, -42.63329, -42.66262, -42.69173, -42.71894, 
        -42.74381, -42.76503, -42.78217, -42.79487, -42.80418, -42.80956, 
        -42.81077, -42.80929, -42.80526, -42.79813, -42.78856, -42.7769, 
        -42.76205, -42.74268, -42.72031, -42.69361, -42.66217, -42.6263, 
        -42.58608, -42.54257, -42.4966, -42.45, -42.40422, -42.36085, 
        -42.31945, -42.27841, -42.23644, -42.18704, -42.1286, -42.05925, 
        -41.97974, -41.88741, -41.79533, -41.70176, -41.60723, -41.51222, 
        -41.41806, -41.31711, -41.21804, -41.12366, -41.03587, -40.95296, 
        -40.85572, -40.77316, -40.69093, -40.61194, -40.52948, -40.46719, 
        -40.41413, -40.36151, -40.30886, -40.26303, -40.22679, -40.17962, 
        -40.128, -40.07052, -40.0122, -39.9447, -39.89423, -39.85274, 
        -39.82492, -39.80381, -39.78988, -39.8029, -39.8296, -39.83276, 
        -39.81052, -39.77836, -39.72758, -39.67213, -39.57717, -39.47798, 
        -39.41655, -39.35843, -39.32035, -39.2847, -39.26105, -39.25573, 
        -39.25027, -39.22047, -39.20292, -39.18534, -39.13839, -39.08758, 
        -39.05799, -39.0429, -39.01292, -38.99389, -38.97935, -38.98589, 
        -38.9998, -39.018, -39.04546, -39.0833, -39.13187, -39.19153, 
        -39.2258, -39.23532, -39.27209, -39.32281, -39.37527, -39.41974, 
        -39.47739, -39.54033, -39.60445, -39.66143, -39.71473, -39.75658, 
        -39.78908, -39.82136, -39.85307, -39.89561, -39.93232, -39.95993, 
        -39.97961, -39.98984, -40.01685, -40.04935, -40.07816, -40.12716, 
        -40.2199, -40.29947, -40.35475, -40.45836, -40.56329, -40.66154, 
        -40.74084, -40.8132, -40.88469, -40.97047, -41.04058, -41.10672, 
        -41.1684, -41.22647, -41.28109, -41.32801, -41.36903, -41.40283, 
        -41.43295, -41.46109, -41.49016, -41.52146, -41.55432, -41.58722, 
        -41.61866, -41.6478, -41.67275, -41.69985, -41.72727, -41.75718, 
        -41.78951, -41.82442, -41.86288, -41.90403, -41.94629, -41.9884, 
        -42.03151, -42.07132, -42.10896, -42.14405, -42.17831, -42.21293, 
        -42.24945, -42.28676, -42.3239, -42.35799, -42.38361, -42.40943, 
        -42.42961, -42.44206, -42.44719, -42.45107, -42.44679, -42.43932, 
        -42.43159, -42.42508, -42.42088, -42.41654, -42.41366, -42.41214, 
        -42.41307, -42.42097, -42.43295, -42.4541, -42.48632, -42.53147, 
        -42.58741, -42.66236, -42.75248, -42.85628, -42.97051, -43.08831, 
        -43.21075, -43.3298, -43.44115, -43.54174, -43.63319, -43.71325, 
        -43.78583, -43.8534, -43.91939, -43.98667, -44.05541, -44.12584, 
        -44.19624, -44.263, -44.32349, -44.37502, -44.41575, -44.44601, 
        -44.46831, -44.48647, -44.5041, -44.52653, -44.55727, -44.59644, 
        -44.64161, -44.6894, -44.73561, -44.77473, -44.80305, -44.81823, 
        -44.8197, -44.80883, -44.78849, -44.76183, -44.73211, -44.70113, 
        -44.67002,
  -38.69169, -38.72759, -38.75677, -38.77804, -38.79098, -38.79642, 
        -38.79569, -38.78955, -38.77894, -38.76562, -38.74961, -38.73296, 
        -38.71624, -38.70181, -38.69202, -38.69069, -38.70284, -38.73171, 
        -38.77657, -38.83858, -38.9197, -39.01829, -39.13203, -39.25893, 
        -39.39485, -39.53924, -39.69032, -39.84843, -40.01161, -40.17837, 
        -40.34621, -40.51688, -40.68885, -40.86097, -41.03006, -41.19543, 
        -41.35296, -41.5008, -41.63875, -41.76612, -41.8806, -41.9844, 
        -42.0787, -42.16492, -42.24486, -42.31985, -42.38869, -42.45258, 
        -42.50929, -42.55662, -42.59404, -42.62085, -42.63697, -42.64249, 
        -42.63773, -42.62457, -42.6043, -42.57942, -42.55152, -42.52287, 
        -42.49499, -42.47005, -42.44944, -42.43698, -42.43353, -42.43897, 
        -42.45237, -42.47243, -42.4979, -42.52464, -42.55196, -42.57943, 
        -42.60534, -42.62753, -42.64602, -42.65998, -42.66986, -42.67538, 
        -42.67641, -42.6732, -42.66747, -42.65746, -42.64532, -42.63071, 
        -42.61278, -42.59117, -42.56512, -42.53405, -42.49805, -42.4569, 
        -42.41068, -42.36052, -42.30712, -42.25323, -42.19931, -42.14877, 
        -42.10134, -42.05589, -42.0123, -41.96321, -41.90664, -41.84099, 
        -41.76721, -41.68086, -41.59494, -41.5078, -41.41927, -41.33029, 
        -41.24061, -41.14484, -41.04708, -40.95288, -40.86242, -40.78152, 
        -40.68372, -40.59666, -40.50966, -40.42388, -40.34198, -40.27243, 
        -40.21561, -40.1579, -40.1054, -40.07278, -40.03932, -39.98598, 
        -39.93075, -39.88393, -39.82936, -39.78004, -39.7204, -39.66801, 
        -39.6384, -39.60977, -39.58216, -39.59127, -39.62063, -39.62968, 
        -39.60473, -39.57636, -39.5358, -39.48549, -39.42168, -39.32866, 
        -39.24969, -39.18875, -39.1332, -39.09253, -39.07122, -39.06538, 
        -39.04847, -39.01052, -39.00883, -38.98853, -38.92792, -38.8914, 
        -38.87573, -38.86357, -38.84192, -38.82069, -38.79588, -38.79574, 
        -38.80999, -38.8428, -38.87556, -38.91486, -38.96511, -39.02058, 
        -39.04583, -39.06011, -39.09358, -39.1454, -39.19406, -39.24323, 
        -39.30358, -39.37465, -39.45794, -39.52611, -39.58212, -39.62851, 
        -39.66383, -39.69388, -39.7294, -39.78518, -39.83657, -39.88369, 
        -39.91845, -39.95515, -39.99211, -40.03497, -40.07512, -40.12234, 
        -40.20645, -40.3041, -40.38268, -40.4632, -40.55172, -40.63567, 
        -40.71275, -40.7812, -40.85774, -40.93023, -40.99709, -41.06228, 
        -41.12563, -41.18695, -41.24386, -41.29206, -41.3334, -41.3677, 
        -41.39844, -41.42771, -41.45747, -41.49221, -41.52773, -41.56277, 
        -41.59629, -41.62745, -41.65374, -41.68183, -41.71038, -41.74107, 
        -41.77514, -41.813, -41.85356, -41.89667, -41.94147, -41.98777, 
        -42.03659, -42.08309, -42.12845, -42.17258, -42.21667, -42.26181, 
        -42.30858, -42.35526, -42.40087, -42.44271, -42.47543, -42.50627, 
        -42.53022, -42.54554, -42.55453, -42.55997, -42.55836, -42.55187, 
        -42.54597, -42.54024, -42.53611, -42.53129, -42.52696, -42.52394, 
        -42.52378, -42.53061, -42.54282, -42.56514, -42.60075, -42.65023, 
        -42.71281, -42.79271, -42.88727, -42.99396, -43.10878, -43.22485, 
        -43.34216, -43.45312, -43.55424, -43.64236, -43.71922, -43.78461, 
        -43.84195, -43.89452, -43.94571, -43.99936, -44.05576, -44.11501, 
        -44.17596, -44.23546, -44.29111, -44.34035, -44.38166, -44.41474, 
        -44.44337, -44.47038, -44.49776, -44.52941, -44.56574, -44.60812, 
        -44.65239, -44.69444, -44.7303, -44.75651, -44.76938, -44.76926, 
        -44.75525, -44.73139, -44.7, -44.66619, -44.63224, -44.59951, 
        -44.56853,
  -38.75176, -38.78139, -38.80407, -38.81831, -38.82449, -38.8235, 
        -38.81653, -38.80459, -38.78921, -38.77184, -38.7525, -38.73386, 
        -38.71594, -38.69963, -38.68991, -38.6914, -38.70546, -38.73608, 
        -38.78297, -38.84405, -38.92369, -39.01985, -39.12954, -39.25178, 
        -39.38285, -39.52225, -39.67174, -39.83061, -39.99652, -40.16859, 
        -40.34467, -40.52349, -40.70359, -40.88327, -41.05986, -41.23116, 
        -41.39488, -41.55016, -41.69473, -41.82671, -41.94502, -42.05239, 
        -42.14924, -42.23738, -42.31816, -42.39305, -42.46205, -42.52381, 
        -42.57673, -42.61966, -42.65094, -42.67027, -42.67811, -42.67394, 
        -42.6585, -42.63367, -42.59946, -42.56087, -42.5189, -42.4751, 
        -42.43239, -42.39291, -42.35959, -42.33551, -42.32235, -42.32001, 
        -42.32711, -42.34179, -42.36435, -42.3898, -42.41722, -42.44503, 
        -42.473, -42.49671, -42.51722, -42.5334, -42.5451, -42.55209, 
        -42.55417, -42.55188, -42.54556, -42.53564, -42.52216, -42.50605, 
        -42.48631, -42.46247, -42.43305, -42.39792, -42.35666, -42.30933, 
        -42.25624, -42.19753, -42.13625, -42.07328, -42.01139, -41.95319, 
        -41.89991, -41.85036, -41.80362, -41.75318, -41.69747, -41.63466, 
        -41.56433, -41.48327, -41.40333, -41.32172, -41.23919, -41.15622, 
        -41.07372, -40.98503, -40.89273, -40.80119, -40.71076, -40.62553, 
        -40.52822, -40.43963, -40.34978, -40.26446, -40.17253, -40.09918, 
        -40.0317, -39.97961, -39.93837, -39.90311, -39.857, -39.79714, 
        -39.73497, -39.70316, -39.66336, -39.60599, -39.56588, -39.51784, 
        -39.47614, -39.44416, -39.4164, -39.40765, -39.42885, -39.44118, 
        -39.41143, -39.37472, -39.34422, -39.30951, -39.26264, -39.19928, 
        -39.13159, -39.06396, -38.99841, -38.92628, -38.88762, -38.8974, 
        -38.87201, -38.83453, -38.81822, -38.81366, -38.76662, -38.73148, 
        -38.72183, -38.70188, -38.67855, -38.66682, -38.6494, -38.64957, 
        -38.66862, -38.70103, -38.74892, -38.79752, -38.84049, -38.86589, 
        -38.88519, -38.89473, -38.93066, -38.98092, -39.02731, -39.07803, 
        -39.13536, -39.22242, -39.31142, -39.38538, -39.44677, -39.49839, 
        -39.54521, -39.58745, -39.63404, -39.68721, -39.74756, -39.80305, 
        -39.854, -39.90285, -39.94933, -39.99878, -40.05697, -40.12608, 
        -40.20841, -40.29677, -40.38063, -40.4616, -40.541, -40.61926, 
        -40.69671, -40.77074, -40.84192, -40.90863, -40.97343, -41.03844, 
        -41.10001, -41.16013, -41.21815, -41.26412, -41.30509, -41.33875, 
        -41.36945, -41.39971, -41.43409, -41.47178, -41.51032, -41.54836, 
        -41.58438, -41.61718, -41.64437, -41.67312, -41.70229, -41.73376, 
        -41.76939, -41.80961, -41.85327, -41.90005, -41.94967, -42.00205, 
        -42.05751, -42.11213, -42.16711, -42.22178, -42.27695, -42.33229, 
        -42.38941, -42.44601, -42.50047, -42.55023, -42.59033, -42.62615, 
        -42.65388, -42.67313, -42.68484, -42.69302, -42.69444, -42.69187, 
        -42.68813, -42.68391, -42.68023, -42.67498, -42.66974, -42.66499, 
        -42.663, -42.668, -42.67982, -42.70332, -42.74077, -42.7933, 
        -42.85985, -42.94238, -43.03717, -43.14196, -43.25212, -43.36106, 
        -43.46758, -43.56544, -43.65119, -43.72311, -43.78297, -43.83149, 
        -43.87136, -43.9082, -43.94497, -43.98533, -44.03038, -44.08043, 
        -44.13428, -44.18935, -44.24278, -44.29301, -44.3379, -44.37795, 
        -44.4153, -44.4517, -44.48976, -44.5306, -44.57437, -44.61893, 
        -44.66085, -44.6963, -44.72195, -44.7348, -44.73361, -44.71823, 
        -44.69034, -44.655, -44.61499, -44.5758, -44.53959, -44.50765, -44.479,
  -38.79949, -38.82362, -38.84074, -38.84898, -38.84961, -38.84253, 
        -38.83014, -38.81324, -38.79386, -38.77303, -38.75252, -38.73314, 
        -38.71434, -38.69802, -38.68984, -38.69187, -38.70707, -38.73932, 
        -38.7847, -38.84563, -38.92076, -39.01221, -39.11541, -39.22918, 
        -39.35366, -39.48882, -39.63353, -39.79101, -39.9592, -40.13662, 
        -40.32039, -40.50877, -40.69874, -40.8882, -41.0746, -41.25438, 
        -41.42745, -41.59149, -41.74422, -41.88424, -42.01048, -42.12404, 
        -42.22581, -42.31739, -42.40063, -42.4761, -42.54392, -42.60357, 
        -42.65269, -42.69022, -42.71471, -42.7255, -42.72474, -42.71094, 
        -42.68455, -42.64767, -42.60134, -42.54858, -42.49212, -42.4331, 
        -42.37514, -42.3207, -42.27373, -42.23787, -42.21469, -42.20354, 
        -42.20488, -42.2137, -42.23275, -42.25681, -42.28518, -42.31666, 
        -42.34744, -42.37547, -42.39886, -42.41785, -42.43228, -42.44154, 
        -42.44523, -42.44447, -42.4395, -42.43022, -42.41721, -42.401, 
        -42.38036, -42.35416, -42.32188, -42.28255, -42.2357, -42.1817, 
        -42.12112, -42.05487, -41.98463, -41.91327, -41.84318, -41.77767, 
        -41.71785, -41.66344, -41.61249, -41.55927, -41.5032, -41.44152, 
        -41.37449, -41.29731, -41.22281, -41.14648, -41.06993, -40.99187, 
        -40.91473, -40.83437, -40.74826, -40.66096, -40.57065, -40.48441, 
        -40.39561, -40.30826, -40.21616, -40.12841, -40.03841, -39.95409, 
        -39.8815, -39.82096, -39.78872, -39.74076, -39.69016, -39.63265, 
        -39.57391, -39.54723, -39.50193, -39.45638, -39.42201, -39.37293, 
        -39.34418, -39.30616, -39.26799, -39.25975, -39.27876, -39.26638, 
        -39.2546, -39.20988, -39.16872, -39.1453, -39.1118, -39.05973, 
        -38.98702, -38.917, -38.85782, -38.80294, -38.75008, -38.75641, 
        -38.7173, -38.69585, -38.67641, -38.67777, -38.64909, -38.6113, 
        -38.5941, -38.56821, -38.54777, -38.54067, -38.52448, -38.53374, 
        -38.548, -38.57806, -38.6165, -38.67557, -38.71181, -38.72499, 
        -38.73553, -38.74895, -38.78331, -38.83041, -38.87922, -38.93317, 
        -38.99733, -39.07822, -39.16071, -39.24577, -39.30947, -39.36024, 
        -39.41746, -39.48844, -39.55293, -39.60907, -39.66351, -39.72826, 
        -39.78403, -39.84194, -39.89573, -39.94994, -40.01454, -40.09219, 
        -40.17966, -40.27276, -40.36155, -40.45183, -40.53517, -40.61258, 
        -40.69066, -40.7682, -40.83927, -40.90686, -40.97302, -41.03275, 
        -41.09361, -41.15208, -41.20437, -41.24847, -41.28765, -41.32194, 
        -41.35361, -41.38635, -41.42485, -41.46677, -41.50847, -41.5495, 
        -41.58765, -41.62209, -41.64944, -41.6783, -41.70813, -41.74112, 
        -41.77726, -41.82021, -41.86747, -41.91953, -41.9753, -42.03455, 
        -42.09803, -42.16224, -42.22816, -42.29423, -42.36139, -42.42891, 
        -42.49685, -42.56419, -42.62832, -42.68605, -42.73462, -42.7765, 
        -42.80867, -42.83172, -42.84726, -42.8578, -42.86229, -42.86246, 
        -42.86083, -42.85776, -42.85329, -42.84723, -42.84064, -42.83361, 
        -42.8288, -42.83043, -42.841, -42.86411, -42.90088, -42.95475, 
        -43.02249, -43.10411, -43.19613, -43.29386, -43.39456, -43.49135, 
        -43.58224, -43.6624, -43.7298, -43.783, -43.82403, -43.85467, 
        -43.87881, -43.90039, -43.92379, -43.95244, -43.98827, -44.03092, 
        -44.08095, -44.13402, -44.18913, -44.24271, -44.29335, -44.34184, 
        -44.38932, -44.43636, -44.48392, -44.53281, -44.58144, -44.6266, 
        -44.66516, -44.6949, -44.71088, -44.71186, -44.69728, -44.66867, 
        -44.62969, -44.58442, -44.53785, -44.49461, -44.45799, -44.42815, 
        -44.40345,
  -38.83424, -38.85369, -38.86597, -38.87021, -38.86717, -38.85686, 
        -38.8403, -38.82023, -38.79813, -38.77533, -38.75362, -38.73343, 
        -38.7148, -38.69886, -38.6895, -38.69262, -38.70939, -38.74031, 
        -38.78423, -38.84221, -38.91283, -38.99606, -39.09065, -39.1966, 
        -39.31296, -39.44109, -39.58163, -39.73623, -39.90477, -40.0862, 
        -40.27641, -40.47388, -40.67472, -40.87574, -41.07374, -41.26611, 
        -41.45055, -41.62526, -41.78863, -41.93816, -42.07386, -42.19514, 
        -42.30336, -42.39962, -42.48554, -42.5611, -42.62849, -42.68567, 
        -42.7307, -42.76276, -42.78099, -42.7856, -42.77611, -42.75259, 
        -42.71531, -42.6663, -42.6072, -42.54077, -42.46947, -42.39635, 
        -42.32383, -42.25507, -42.19402, -42.14618, -42.11305, -42.09346, 
        -42.08881, -42.09518, -42.11194, -42.13523, -42.16277, -42.1973, 
        -42.2323, -42.26435, -42.2924, -42.31464, -42.33142, -42.34265, 
        -42.34923, -42.34982, -42.34675, -42.33921, -42.32787, -42.31224, 
        -42.29171, -42.26447, -42.22942, -42.18637, -42.13447, -42.07407, 
        -42.00541, -41.9306, -41.85158, -41.77145, -41.69365, -41.62132, 
        -41.55523, -41.49391, -41.43811, -41.38229, -41.325, -41.26384, 
        -41.1991, -41.12718, -41.0568, -40.98558, -40.91389, -40.84174, 
        -40.76939, -40.69464, -40.61079, -40.52517, -40.43728, -40.34845, 
        -40.25819, -40.17836, -40.0975, -40.01242, -39.92812, -39.83419, 
        -39.75764, -39.69452, -39.64559, -39.59245, -39.53139, -39.48571, 
        -39.42744, -39.3955, -39.36254, -39.31882, -39.29055, -39.24537, 
        -39.2146, -39.17912, -39.16238, -39.15086, -39.142, -39.10958, 
        -39.10109, -39.07915, -39.04413, -39.00401, -38.9728, -38.91463, 
        -38.8386, -38.77127, -38.72443, -38.6826, -38.64494, -38.64963, 
        -38.62223, -38.60414, -38.59123, -38.57827, -38.57193, -38.5416, 
        -38.5097, -38.48014, -38.4653, -38.45714, -38.44886, -38.45429, 
        -38.46928, -38.49067, -38.52758, -38.56969, -38.59385, -38.5981, 
        -38.60434, -38.6376, -38.66615, -38.70772, -38.75209, -38.80594, 
        -38.86959, -38.94488, -39.03394, -39.11238, -39.17636, -39.23462, 
        -39.31065, -39.39196, -39.46846, -39.53561, -39.59555, -39.66237, 
        -39.73053, -39.79557, -39.85373, -39.91798, -39.98814, -40.07925, 
        -40.17125, -40.26336, -40.35967, -40.45301, -40.53972, -40.62003, 
        -40.69874, -40.77453, -40.8469, -40.91496, -40.9808, -41.04094, 
        -41.09892, -41.15149, -41.19847, -41.24016, -41.27896, -41.31371, 
        -41.34875, -41.38513, -41.42617, -41.47168, -41.51508, -41.55838, 
        -41.59883, -41.63505, -41.66484, -41.69615, -41.7284, -41.76307, 
        -41.8036, -41.85018, -41.90293, -41.96138, -42.02442, -42.09246, 
        -42.16481, -42.23954, -42.3163, -42.39378, -42.47216, -42.55087, 
        -42.62952, -42.70653, -42.77914, -42.84421, -42.8997, -42.94622, 
        -42.9826, -43.00951, -43.02821, -43.04159, -43.04843, -43.05164, 
        -43.05234, -43.05125, -43.04791, -43.04244, -43.03473, -43.02586, 
        -43.01897, -43.01839, -43.02699, -43.04848, -43.08548, -43.13764, 
        -43.20304, -43.27935, -43.36364, -43.45037, -43.53603, -43.61563, 
        -43.68699, -43.74648, -43.79262, -43.82553, -43.8471, -43.85988, 
        -43.86821, -43.87615, -43.88758, -43.90736, -43.93657, -43.97606, 
        -44.02411, -44.07805, -44.13688, -44.19606, -44.25446, -44.31193, 
        -44.36891, -44.42529, -44.47982, -44.53426, -44.58588, -44.63116, 
        -44.66634, -44.6897, -44.69758, -44.68873, -44.66383, -44.62528, 
        -44.577, -44.52436, -44.47265, -44.42692, -44.39062, -44.36357, 
        -44.34325,
  -38.85939, -38.87497, -38.88396, -38.88554, -38.8799, -38.86779, 
        -38.84926, -38.8275, -38.80403, -38.77978, -38.75772, -38.73743, 
        -38.71931, -38.70526, -38.69545, -38.69904, -38.71481, -38.74392, 
        -38.78561, -38.83802, -38.90103, -38.97612, -39.06173, -39.15833, 
        -39.26569, -39.38648, -39.52103, -39.67164, -39.83945, -40.02309, 
        -40.21977, -40.42564, -40.63679, -40.84978, -41.06051, -41.26583, 
        -41.46284, -41.64965, -41.82471, -41.98564, -42.13, -42.26079, 
        -42.37651, -42.47836, -42.56777, -42.64581, -42.71231, -42.76699, 
        -42.80836, -42.83547, -42.84782, -42.84548, -42.82782, -42.7948, 
        -42.74695, -42.68694, -42.61505, -42.53617, -42.4518, -42.36506, 
        -42.27895, -42.19684, -42.12426, -42.06497, -42.02227, -41.99548, 
        -41.98336, -41.98641, -42.00045, -42.02448, -42.05544, -42.09192, 
        -42.13004, -42.16537, -42.19718, -42.22287, -42.24256, -42.2567, 
        -42.26515, -42.26963, -42.26896, -42.2637, -42.25406, -42.23942, 
        -42.2186, -42.19011, -42.15324, -42.10674, -42.04981, -41.98284, 
        -41.90679, -41.82234, -41.73479, -41.6467, -41.56172, -41.48283, 
        -41.41099, -41.34538, -41.28516, -41.22584, -41.16713, -41.10672, 
        -41.04368, -40.97512, -40.90783, -40.84007, -40.77219, -40.70454, 
        -40.63634, -40.56561, -40.48822, -40.40762, -40.32668, -40.24657, 
        -40.16198, -40.08714, -40.00471, -39.91897, -39.82148, -39.72564, 
        -39.64606, -39.58025, -39.53426, -39.47865, -39.42304, -39.36931, 
        -39.31611, -39.27762, -39.24743, -39.201, -39.1631, -39.12774, 
        -39.09775, -39.06946, -39.04758, -39.03707, -39.03896, -39.01009, 
        -38.97454, -38.96202, -38.93959, -38.90815, -38.86573, -38.80853, 
        -38.74701, -38.68336, -38.63711, -38.60717, -38.58599, -38.5918, 
        -38.58111, -38.56904, -38.58011, -38.5587, -38.53955, -38.50837, 
        -38.47626, -38.44875, -38.43518, -38.41311, -38.40247, -38.40405, 
        -38.41547, -38.4327, -38.45267, -38.4861, -38.50384, -38.51271, 
        -38.5059, -38.5301, -38.56432, -38.59937, -38.63866, -38.6867, 
        -38.74204, -38.81012, -38.8879, -38.97442, -39.05226, -39.1249, 
        -39.21849, -39.30792, -39.38783, -39.45481, -39.51869, -39.59917, 
        -39.67582, -39.75246, -39.82415, -39.90215, -39.97937, -40.06899, 
        -40.16463, -40.26306, -40.36596, -40.46212, -40.55304, -40.63504, 
        -40.71537, -40.78978, -40.86138, -40.92825, -40.99248, -41.05003, 
        -41.10605, -41.15641, -41.20138, -41.24289, -41.28304, -41.32056, 
        -41.35983, -41.40202, -41.44724, -41.49545, -41.54041, -41.58424, 
        -41.6264, -41.66684, -41.70064, -41.73555, -41.7715, -41.81062, 
        -41.85452, -41.90614, -41.96589, -42.03164, -42.10328, -42.18017, 
        -42.26186, -42.34621, -42.43338, -42.52156, -42.60904, -42.69788, 
        -42.78571, -42.87123, -42.95039, -43.0218, -43.08363, -43.13478, 
        -43.17484, -43.20565, -43.22787, -43.24379, -43.25428, -43.25997, 
        -43.26285, -43.2634, -43.26097, -43.25549, -43.24706, -43.23704, 
        -43.22834, -43.2254, -43.23149, -43.25052, -43.28432, -43.3322, 
        -43.39148, -43.45945, -43.53153, -43.60326, -43.67072, -43.72979, 
        -43.779, -43.81596, -43.83998, -43.85199, -43.85463, -43.85004, 
        -43.84459, -43.84133, -43.84456, -43.85791, -43.88341, -43.92217, 
        -43.97126, -44.0286, -44.09201, -44.15792, -44.22432, -44.29007, 
        -44.35513, -44.41869, -44.48003, -44.53789, -44.59024, -44.63446, 
        -44.66649, -44.68468, -44.68642, -44.67064, -44.63856, -44.59304, 
        -44.5385, -44.48055, -44.42506, -44.37763, -44.34143, -44.31652, 
        -44.29998,
  -38.87606, -38.88888, -38.89592, -38.89638, -38.8903, -38.87635, 
        -38.85819, -38.83678, -38.81387, -38.79142, -38.77013, -38.75004, 
        -38.73303, -38.72032, -38.71352, -38.71632, -38.72964, -38.75506, 
        -38.7918, -38.83829, -38.89404, -38.96091, -39.03779, -39.12423, 
        -39.22254, -39.33671, -39.46544, -39.61067, -39.77517, -39.95858, 
        -40.15784, -40.36958, -40.58971, -40.81359, -41.03577, -41.25412, 
        -41.4645, -41.66447, -41.85182, -42.02432, -42.18052, -42.32038, 
        -42.44416, -42.55211, -42.6452, -42.72475, -42.79082, -42.84309, 
        -42.88064, -42.90363, -42.91054, -42.9019, -42.87667, -42.83514, 
        -42.77786, -42.70777, -42.62647, -42.53721, -42.44161, -42.34336, 
        -42.24498, -42.15111, -42.0673, -41.99763, -41.9461, -41.91224, 
        -41.89536, -41.89292, -41.90577, -41.92863, -41.96093, -41.99955, 
        -42.04047, -42.08073, -42.11685, -42.14631, -42.16924, -42.18618, 
        -42.19733, -42.20371, -42.20454, -42.20114, -42.19286, -42.17913, 
        -42.15714, -42.12798, -42.08958, -42.03983, -41.97852, -41.90556, 
        -41.82248, -41.73195, -41.63653, -41.5415, -41.4502, -41.36515, 
        -41.2877, -41.217, -41.15258, -41.09055, -41.03021, -40.97042, 
        -40.9088, -40.84188, -40.77665, -40.711, -40.64536, -40.58022, 
        -40.51513, -40.44927, -40.37821, -40.30443, -40.22897, -40.15544, 
        -40.08051, -40.00737, -39.93099, -39.84708, -39.74645, -39.65535, 
        -39.56997, -39.49742, -39.44452, -39.39882, -39.35373, -39.30106, 
        -39.24916, -39.20253, -39.16709, -39.12733, -39.07944, -39.03455, 
        -38.99833, -38.97314, -38.95278, -38.94985, -38.94374, -38.9339, 
        -38.90248, -38.88482, -38.87263, -38.86617, -38.83229, -38.79818, 
        -38.75122, -38.69942, -38.64343, -38.60753, -38.59378, -38.59649, 
        -38.62124, -38.6166, -38.61602, -38.59562, -38.56355, -38.53668, 
        -38.49408, -38.46963, -38.45677, -38.42352, -38.38636, -38.37482, 
        -38.37273, -38.37762, -38.38385, -38.40172, -38.43564, -38.44373, 
        -38.44907, -38.4627, -38.48852, -38.5157, -38.54784, -38.5918, 
        -38.63872, -38.68045, -38.75698, -38.85729, -38.94237, -39.01936, 
        -39.12926, -39.23023, -39.31124, -39.38982, -39.4537, -39.53636, 
        -39.62188, -39.71033, -39.7981, -39.89353, -39.98906, -40.08141, 
        -40.17604, -40.2774, -40.38102, -40.48105, -40.57389, -40.65822, 
        -40.73952, -40.81432, -40.88522, -40.9521, -41.01493, -41.07132, 
        -41.12543, -41.17457, -41.21928, -41.26145, -41.30368, -41.34605, 
        -41.3915, -41.43846, -41.4871, -41.53759, -41.58089, -41.62505, 
        -41.67032, -41.7179, -41.75915, -41.80048, -41.84171, -41.88499, 
        -41.93555, -41.99418, -42.06154, -42.13548, -42.21569, -42.30097, 
        -42.39079, -42.48367, -42.57921, -42.67586, -42.77248, -42.86941, 
        -42.96435, -43.05572, -43.14078, -43.21688, -43.28307, -43.33845, 
        -43.38247, -43.41607, -43.44145, -43.45973, -43.47233, -43.47993, 
        -43.48406, -43.48537, -43.48307, -43.4777, -43.46868, -43.45744, 
        -43.44702, -43.44129, -43.44471, -43.45924, -43.48813, -43.52897, 
        -43.5793, -43.63538, -43.69281, -43.7464, -43.79322, -43.83007, 
        -43.8562, -43.87, -43.87198, -43.86432, -43.84962, -43.83197, 
        -43.81575, -43.80478, -43.80309, -43.81414, -43.83955, -43.87919, 
        -43.93083, -43.99239, -44.06064, -44.13271, -44.20565, -44.27795, 
        -44.34922, -44.41747, -44.4819, -44.54121, -44.59324, -44.63542, 
        -44.66476, -44.67939, -44.67722, -44.65741, -44.62165, -44.57243, 
        -44.51416, -44.45305, -44.39519, -44.34645, -44.31011, -44.28626, 
        -44.26984,
  -38.88608, -38.89731, -38.90358, -38.90432, -38.89885, -38.8873, 
        -38.87139, -38.8521, -38.83164, -38.81125, -38.79164, -38.773, 
        -38.75709, -38.74542, -38.73914, -38.7418, -38.75352, -38.77534, 
        -38.80768, -38.84888, -38.89896, -38.95886, -39.02858, -39.10746, 
        -39.19791, -39.30214, -39.42381, -39.56196, -39.72104, -39.90023, 
        -40.09907, -40.31349, -40.5394, -40.77209, -41.00638, -41.23741, 
        -41.46087, -41.67333, -41.87313, -42.05691, -42.2234, -42.37233, 
        -42.50364, -42.61725, -42.71413, -42.79395, -42.85932, -42.91043, 
        -42.94608, -42.96553, -42.96896, -42.95558, -42.92412, -42.87521, 
        -42.80989, -42.73146, -42.64177, -42.54394, -42.43927, -42.33204, 
        -42.22415, -42.11926, -42.026, -41.9477, -41.88873, -41.84776, 
        -41.82698, -41.82243, -41.83226, -41.85425, -41.88649, -41.92621, 
        -41.96943, -42.01257, -42.0521, -42.08551, -42.11181, -42.13133, 
        -42.14357, -42.15125, -42.15334, -42.15046, -42.14256, -42.12893, 
        -42.10775, -42.07806, -42.03819, -41.98593, -41.92097, -41.84332, 
        -41.7546, -41.65788, -41.55639, -41.45577, -41.35871, -41.26834, 
        -41.18475, -41.10924, -41.04052, -40.97621, -40.91451, -40.85473, 
        -40.79401, -40.72981, -40.66573, -40.60077, -40.53607, -40.47145, 
        -40.40746, -40.3447, -40.27734, -40.21542, -40.14592, -40.08179, 
        -40.01116, -39.9381, -39.86651, -39.78677, -39.70889, -39.62788, 
        -39.54694, -39.47774, -39.42631, -39.38631, -39.35024, -39.29211, 
        -39.24862, -39.20288, -39.1506, -39.10615, -39.05658, -39.00632, 
        -38.96714, -38.93691, -38.90859, -38.90128, -38.88625, -38.86923, 
        -38.85215, -38.85963, -38.86617, -38.85069, -38.84359, -38.8327, 
        -38.79731, -38.77073, -38.72578, -38.67897, -38.662, -38.66338, 
        -38.69308, -38.68922, -38.66603, -38.6435, -38.60529, -38.5706, 
        -38.53313, -38.51716, -38.49223, -38.45397, -38.41288, -38.3806, 
        -38.36557, -38.35488, -38.34774, -38.34672, -38.36195, -38.39196, 
        -38.40153, -38.41589, -38.43468, -38.45554, -38.48588, -38.52137, 
        -38.5559, -38.5971, -38.66039, -38.75328, -38.84576, -38.95445, 
        -39.06517, -39.16883, -39.25269, -39.33389, -39.40842, -39.49616, 
        -39.5923, -39.69067, -39.78726, -39.89194, -39.99779, -40.10085, 
        -40.20415, -40.30706, -40.41042, -40.51169, -40.60638, -40.69304, 
        -40.77754, -40.85423, -40.92573, -40.99227, -41.05415, -41.10929, 
        -41.1618, -41.20947, -41.25291, -41.29596, -41.34221, -41.3894, 
        -41.43677, -41.48723, -41.5396, -41.59451, -41.6418, -41.68921, 
        -41.7402, -41.79467, -41.84464, -41.89354, -41.94152, -41.99218, 
        -42.05449, -42.12097, -42.19632, -42.27805, -42.36593, -42.45834, 
        -42.55458, -42.65351, -42.7547, -42.8567, -42.95862, -43.06046, 
        -43.15983, -43.25481, -43.34307, -43.42236, -43.49166, -43.54958, 
        -43.59649, -43.63287, -43.65975, -43.67986, -43.69401, -43.7025, 
        -43.70694, -43.70774, -43.70521, -43.6993, -43.68949, -43.67701, 
        -43.66491, -43.65676, -43.65677, -43.66773, -43.68986, -43.72157, 
        -43.76039, -43.80221, -43.84246, -43.87651, -43.9016, -43.91607, 
        -43.9191, -43.91111, -43.89241, -43.86677, -43.83751, -43.80895, 
        -43.78559, -43.77078, -43.76799, -43.7796, -43.80682, -43.84911, 
        -43.90367, -43.96838, -44.04093, -44.11716, -44.19504, -44.27128, 
        -44.34571, -44.41558, -44.48131, -44.54033, -44.5909, -44.63118, 
        -44.6586, -44.67134, -44.66762, -44.646, -44.60921, -44.55898, 
        -44.50068, -44.43834, -44.37958, -44.3298, -44.29257, -44.26785, 
        -44.25198,
  -38.89541, -38.90625, -38.91306, -38.91475, -38.91092, -38.90237, 
        -38.8898, -38.87436, -38.85752, -38.83943, -38.82204, -38.80568, 
        -38.79204, -38.78264, -38.77797, -38.78023, -38.79138, -38.80989, 
        -38.83717, -38.87331, -38.91787, -38.97107, -39.03365, -39.10661, 
        -39.18972, -39.28659, -39.39982, -39.53181, -39.68393, -39.85848, 
        -40.05399, -40.2675, -40.49601, -40.73433, -40.97766, -41.21926, 
        -41.45432, -41.67904, -41.88968, -42.08274, -42.25837, -42.41533, 
        -42.55313, -42.67141, -42.77174, -42.85443, -42.92058, -42.97067, 
        -43.00526, -43.02273, -43.02312, -43.00568, -42.96931, -42.91531, 
        -42.84356, -42.75766, -42.66148, -42.55657, -42.44454, -42.33, 
        -42.21479, -42.10406, -42.00354, -41.9181, -41.85103, -41.80135, 
        -41.77737, -41.77254, -41.77893, -41.80347, -41.83371, -41.872, 
        -41.91512, -41.96044, -42.0029, -42.03984, -42.06947, -42.09138, 
        -42.10594, -42.11444, -42.11657, -42.11319, -42.10501, -42.09102, 
        -42.0694, -42.03886, -41.99761, -41.94349, -41.87572, -41.79464, 
        -41.70093, -41.5997, -41.49371, -41.38856, -41.28713, -41.19208, 
        -41.10479, -41.02504, -40.95231, -40.88504, -40.8224, -40.76175, 
        -40.70121, -40.63841, -40.57469, -40.51006, -40.44424, -40.37926, 
        -40.31468, -40.25199, -40.18964, -40.12792, -40.07105, -40.00929, 
        -39.94568, -39.88059, -39.81287, -39.74548, -39.67619, -39.61019, 
        -39.54831, -39.49622, -39.44854, -39.39835, -39.3633, -39.30289, 
        -39.27775, -39.24697, -39.19967, -39.15042, -39.09557, -39.03648, 
        -38.99951, -38.9777, -38.91824, -38.88819, -38.87534, -38.87685, 
        -38.86792, -38.86774, -38.88251, -38.88335, -38.86161, -38.86301, 
        -38.85709, -38.83025, -38.80547, -38.78218, -38.7714, -38.76847, 
        -38.76924, -38.74768, -38.71532, -38.68899, -38.63667, -38.61554, 
        -38.58188, -38.55997, -38.55244, -38.52074, -38.48065, -38.43538, 
        -38.3969, -38.36944, -38.34225, -38.32653, -38.32096, -38.33311, 
        -38.35025, -38.3656, -38.38177, -38.39964, -38.42289, -38.45117, 
        -38.47318, -38.50736, -38.56651, -38.65129, -38.76842, -38.88806, 
        -39.00885, -39.11718, -39.20664, -39.29869, -39.38534, -39.48612, 
        -39.5915, -39.69674, -39.80166, -39.91105, -40.02801, -40.14209, 
        -40.2523, -40.35582, -40.45817, -40.55922, -40.65465, -40.7451, 
        -40.83363, -40.91415, -40.987, -41.0528, -41.11392, -41.16841, 
        -41.21826, -41.26311, -41.30577, -41.34847, -41.39449, -41.44183, 
        -41.49616, -41.55449, -41.61657, -41.67852, -41.73536, -41.79076, 
        -41.84663, -41.9073, -41.96581, -42.02474, -42.08195, -42.14299, 
        -42.21079, -42.28576, -42.36826, -42.45743, -42.55193, -42.6497, 
        -42.75005, -42.85215, -42.95578, -43.05843, -43.1619, -43.26484, 
        -43.36512, -43.46093, -43.54987, -43.62975, -43.69986, -43.75908, 
        -43.80754, -43.84578, -43.87563, -43.89772, -43.91281, -43.92135, 
        -43.92567, -43.92661, -43.92329, -43.91584, -43.90465, -43.89072, 
        -43.87736, -43.86721, -43.8633, -43.86814, -43.88203, -43.903, 
        -43.92783, -43.9536, -43.97549, -43.98946, -43.99289, -43.98503, 
        -43.96619, -43.93752, -43.90091, -43.86007, -43.81861, -43.78255, 
        -43.75531, -43.74, -43.73862, -43.75308, -43.78296, -43.82653, 
        -43.88334, -43.95052, -44.02512, -44.10389, -44.18364, -44.26232, 
        -44.33777, -44.4091, -44.47437, -44.53232, -44.58149, -44.62019, 
        -44.64663, -44.65866, -44.65494, -44.63461, -44.59859, -44.55072, 
        -44.49357, -44.43321, -44.37469, -44.32446, -44.28576, -44.2584, 
        -44.23988,
  -38.90746, -38.91932, -38.92733, -38.93061, -38.92826, -38.92356, 
        -38.91529, -38.90431, -38.89193, -38.87831, -38.86405, -38.85087, 
        -38.83985, -38.83222, -38.82907, -38.83112, -38.84012, -38.85614, 
        -38.87963, -38.91018, -38.94955, -38.99818, -39.05549, -39.12243, 
        -39.20186, -39.29349, -39.40048, -39.52518, -39.67049, -39.83805, 
        -40.02774, -40.23807, -40.46571, -40.70758, -40.95478, -41.20472, 
        -41.44923, -41.68333, -41.9037, -42.10604, -42.28923, -42.45243, 
        -42.5954, -42.71772, -42.82127, -42.90631, -42.97385, -43.02437, 
        -43.05855, -43.07508, -43.07253, -43.05233, -43.01291, -42.95556, 
        -42.8801, -42.7914, -42.69032, -42.58066, -42.46382, -42.345, 
        -42.22535, -42.11012, -42.00504, -41.91349, -41.83876, -41.78409, 
        -41.75315, -41.74405, -41.75172, -41.76997, -41.8019, -41.83816, 
        -41.88126, -41.92719, -41.97162, -42.0108, -42.04337, -42.06716, 
        -42.08303, -42.09181, -42.09336, -42.08928, -42.08001, -42.06469, 
        -42.04096, -42.00942, -41.96709, -41.91175, -41.8426, -41.75961, 
        -41.66432, -41.55986, -41.45181, -41.34336, -41.23839, -41.13969, 
        -41.04811, -40.96336, -40.88638, -40.81623, -40.75127, -40.68881, 
        -40.62628, -40.56347, -40.49963, -40.43417, -40.36699, -40.30072, 
        -40.23584, -40.17319, -40.11363, -40.06024, -40.00467, -39.94541, 
        -39.88749, -39.8292, -39.77281, -39.71815, -39.66576, -39.60931, 
        -39.5612, -39.51747, -39.47588, -39.43424, -39.39056, -39.34188, 
        -39.31158, -39.28564, -39.25723, -39.20876, -39.15298, -39.09046, 
        -39.06228, -39.02608, -38.96756, -38.93249, -38.9259, -38.92476, 
        -38.94796, -38.93796, -38.93791, -38.93315, -38.91978, -38.90761, 
        -38.907, -38.91177, -38.89482, -38.86676, -38.85625, -38.8529, 
        -38.84332, -38.81285, -38.7822, -38.74791, -38.70552, -38.68216, 
        -38.65787, -38.63142, -38.61682, -38.58751, -38.547, -38.50665, 
        -38.46438, -38.42289, -38.37261, -38.34668, -38.32128, -38.3177, 
        -38.31413, -38.32801, -38.33899, -38.34483, -38.37374, -38.41286, 
        -38.43712, -38.47246, -38.53283, -38.61214, -38.71634, -38.82597, 
        -38.96236, -39.08022, -39.1825, -39.28416, -39.38869, -39.49926, 
        -39.61618, -39.73152, -39.8446, -39.96168, -40.0794, -40.19711, 
        -40.30806, -40.41246, -40.51535, -40.61815, -40.71882, -40.81638, 
        -40.91071, -40.99646, -41.07383, -41.14153, -41.20211, -41.25608, 
        -41.30519, -41.34909, -41.38977, -41.4311, -41.48497, -41.54396, 
        -41.60152, -41.66845, -41.73246, -41.79745, -41.85912, -41.92332, 
        -41.98808, -42.05415, -42.11956, -42.18634, -42.25254, -42.32502, 
        -42.40145, -42.48395, -42.57372, -42.66924, -42.76831, -42.86954, 
        -42.97099, -43.07298, -43.17557, -43.27796, -43.37976, -43.48085, 
        -43.57932, -43.67311, -43.76074, -43.84033, -43.90959, -43.9687, 
        -44.01746, -44.05713, -44.08771, -44.10984, -44.12477, -44.13298, 
        -44.13646, -44.13486, -44.12919, -44.11972, -44.10627, -44.09043, 
        -44.0739, -44.06047, -44.05088, -44.04819, -44.05247, -44.06155, 
        -44.07205, -44.08117, -44.08416, -44.07808, -44.06077, -44.03259, 
        -43.99425, -43.94743, -43.89585, -43.84382, -43.79533, -43.75494, 
        -43.72631, -43.71258, -43.71355, -43.72926, -43.7609, -43.80653, 
        -43.86457, -43.93153, -44.00655, -44.08532, -44.16545, -44.24406, 
        -44.31981, -44.39056, -44.45488, -44.51157, -44.55962, -44.59755, 
        -44.62367, -44.63572, -44.63354, -44.61586, -44.58334, -44.53892, 
        -44.48578, -44.42816, -44.37208, -44.32173, -44.28031, -44.24971, 
        -44.22697,
  -38.9266, -38.93998, -38.9497, -38.95603, -38.95807, -38.95713, 
        -38.95307, -38.94657, -38.93869, -38.92891, -38.91773, -38.90723, 
        -38.89904, -38.89293, -38.88959, -38.89141, -38.89906, -38.91298, 
        -38.93382, -38.96242, -38.99865, -39.04336, -39.09712, -39.16051, 
        -39.23524, -39.32228, -39.42373, -39.54276, -39.68186, -39.84132, 
        -40.02433, -40.22967, -40.45477, -40.69638, -40.94718, -41.2009, 
        -41.4512, -41.69204, -41.91946, -42.12791, -42.31668, -42.48476, 
        -42.63144, -42.75735, -42.86265, -42.95004, -43.01958, -43.07132, 
        -43.10614, -43.12225, -43.11959, -43.09795, -43.05752, -42.99964, 
        -42.92252, -42.8322, -42.72903, -42.61667, -42.49741, -42.37625, 
        -42.25465, -42.13607, -42.02769, -41.93258, -41.85316, -41.7953, 
        -41.76118, -41.74643, -41.74995, -41.76384, -41.79153, -41.8245, 
        -41.86557, -41.91146, -41.95608, -41.99713, -42.03066, -42.0563, 
        -42.07219, -42.08112, -42.0821, -42.07673, -42.06593, -42.04884, 
        -42.02464, -41.99192, -41.94869, -41.89318, -41.82382, -41.7406, 
        -41.64457, -41.54004, -41.43007, -41.31979, -41.21224, -41.10981, 
        -41.01257, -40.92339, -40.84177, -40.76756, -40.69903, -40.63391, 
        -40.57046, -40.50708, -40.44231, -40.37577, -40.30777, -40.23991, 
        -40.17424, -40.11139, -40.05313, -39.99764, -39.94056, -39.8822, 
        -39.82645, -39.77625, -39.73262, -39.69025, -39.65251, -39.6095, 
        -39.57156, -39.53758, -39.50329, -39.47015, -39.42681, -39.388, 
        -39.36431, -39.33602, -39.31063, -39.26554, -39.22481, -39.19135, 
        -39.15849, -39.11593, -39.06424, -39.03742, -39.03927, -39.02897, 
        -39.03844, -39.0375, -39.03157, -39.02184, -39.01125, -39.00166, 
        -38.98831, -38.99405, -38.98987, -38.96944, -38.95424, -38.93456, 
        -38.92376, -38.87636, -38.8281, -38.80845, -38.79279, -38.76523, 
        -38.73391, -38.70972, -38.68046, -38.64905, -38.60803, -38.56786, 
        -38.52409, -38.48324, -38.43756, -38.39605, -38.37696, -38.35543, 
        -38.31679, -38.3116, -38.32512, -38.3322, -38.35799, -38.39738, 
        -38.43504, -38.47788, -38.54768, -38.64286, -38.72214, -38.81785, 
        -38.94388, -39.06625, -39.17921, -39.29351, -39.40928, -39.53646, 
        -39.66986, -39.79141, -39.90868, -40.02631, -40.13843, -40.25564, 
        -40.37308, -40.48118, -40.58871, -40.6969, -40.80528, -40.91037, 
        -41.01146, -41.1026, -41.18423, -41.25438, -41.31657, -41.37052, 
        -41.42017, -41.46646, -41.51253, -41.56084, -41.61574, -41.67947, 
        -41.74106, -41.80624, -41.87173, -41.94118, -42.01009, -42.08081, 
        -42.15332, -42.22614, -42.29898, -42.37449, -42.45329, -42.53574, 
        -42.62154, -42.71157, -42.80753, -42.90685, -43.00819, -43.10952, 
        -43.21027, -43.31009, -43.40915, -43.50752, -43.60485, -43.70165, 
        -43.79631, -43.88687, -43.97104, -44.04758, -44.11507, -44.17288, 
        -44.22081, -44.25928, -44.28927, -44.31116, -44.32534, -44.33222, 
        -44.33345, -44.32919, -44.32033, -44.30741, -44.29058, -44.27149, 
        -44.25165, -44.23339, -44.21857, -44.20808, -44.20156, -44.19693, 
        -44.19254, -44.18438, -44.1688, -44.14336, -44.10657, -44.05967, 
        -44.00438, -43.94307, -43.87971, -43.81917, -43.76571, -43.72299, 
        -43.69413, -43.68094, -43.68274, -43.69997, -43.73204, -43.77708, 
        -43.83338, -43.89931, -43.97245, -44.05062, -44.1301, -44.20764, 
        -44.28288, -44.35321, -44.41698, -44.47301, -44.52036, -44.55778, 
        -44.58381, -44.59732, -44.59735, -44.58333, -44.55595, -44.51669, 
        -44.46871, -44.41547, -44.36193, -44.31258, -44.27031, -44.23602, 
        -44.20839,
  -38.95953, -38.97492, -38.98714, -38.99608, -39.00157, -39.00412, 
        -39.00421, -39.00203, -38.9976, -38.98977, -38.98171, -38.97366, 
        -38.96743, -38.96302, -38.96095, -38.96272, -38.96928, -38.98166, 
        -39.00098, -39.02766, -39.0622, -39.10498, -39.1566, -39.21659, 
        -39.28839, -39.37217, -39.47007, -39.58429, -39.71799, -39.87243, 
        -40.04956, -40.24911, -40.46946, -40.70694, -40.95641, -41.21098, 
        -41.46315, -41.70701, -41.93759, -42.14901, -42.34157, -42.51258, 
        -42.66187, -42.7907, -42.89968, -42.98943, -43.06058, -43.11391, 
        -43.14917, -43.16567, -43.16386, -43.14307, -43.10302, -43.0457, 
        -42.96998, -42.87881, -42.77628, -42.66419, -42.54442, -42.42356, 
        -42.30222, -42.18459, -42.07516, -41.97832, -41.8995, -41.83767, 
        -41.79466, -41.77252, -41.7713, -41.78145, -41.80059, -41.83056, 
        -41.86765, -41.9101, -41.95397, -41.9947, -42.02914, -42.05595, 
        -42.07339, -42.08271, -42.08271, -42.07592, -42.06326, -42.04436, 
        -42.01873, -41.98512, -41.94176, -41.88677, -41.81847, -41.73545, 
        -41.64112, -41.53738, -41.42817, -41.31676, -41.20673, -41.10049, 
        -40.99949, -40.90524, -40.81863, -40.73941, -40.66616, -40.59757, 
        -40.53147, -40.46645, -40.40094, -40.33369, -40.26471, -40.19613, 
        -40.12894, -40.06615, -40.00489, -39.94577, -39.88299, -39.82333, 
        -39.77347, -39.7303, -39.69629, -39.66591, -39.63786, -39.60612, 
        -39.58157, -39.55559, -39.5279, -39.50106, -39.47068, -39.44266, 
        -39.42365, -39.40416, -39.37395, -39.34965, -39.30951, -39.27378, 
        -39.25457, -39.22848, -39.19607, -39.17048, -39.16518, -39.15765, 
        -39.15224, -39.14246, -39.13942, -39.1318, -39.12402, -39.11437, 
        -39.10973, -39.10525, -39.09516, -39.08345, -39.06594, -39.04249, 
        -39.01486, -38.96829, -38.92698, -38.89666, -38.88259, -38.85076, 
        -38.81264, -38.78706, -38.75422, -38.70805, -38.66179, -38.62039, 
        -38.5787, -38.53759, -38.50032, -38.48407, -38.45947, -38.40767, 
        -38.36562, -38.36712, -38.37912, -38.37334, -38.37097, -38.41297, 
        -38.46289, -38.51883, -38.60899, -38.70644, -38.78149, -38.85949, 
        -38.96182, -39.08038, -39.20007, -39.32527, -39.45461, -39.58323, 
        -39.71564, -39.84461, -39.96651, -40.08976, -40.21157, -40.33322, 
        -40.45235, -40.56598, -40.68002, -40.79573, -40.91143, -41.02394, 
        -41.13246, -41.22896, -41.31359, -41.38658, -41.45025, -41.50513, 
        -41.5563, -41.60658, -41.65834, -41.71327, -41.77089, -41.83188, 
        -41.89742, -41.96444, -42.03289, -42.1064, -42.18089, -42.25737, 
        -42.33593, -42.41656, -42.49862, -42.58434, -42.67345, -42.76606, 
        -42.86126, -42.95762, -43.0568, -43.15861, -43.25938, -43.35908, 
        -43.45674, -43.55245, -43.64543, -43.73801, -43.82969, -43.92078, 
        -44.0101, -44.09573, -44.17571, -44.24854, -44.31296, -44.36821, 
        -44.41435, -44.45173, -44.48042, -44.50072, -44.5128, -44.51769, 
        -44.51578, -44.50803, -44.49548, -44.47793, -44.45688, -44.43327, 
        -44.40853, -44.38422, -44.36172, -44.34186, -44.32379, -44.30568, 
        -44.28566, -44.26007, -44.22656, -44.18263, -44.12828, -44.0651, 
        -43.9954, -43.92258, -43.84959, -43.78326, -43.72651, -43.6824, 
        -43.65312, -43.63939, -43.64054, -43.65611, -43.68594, -43.72797, 
        -43.78068, -43.84399, -43.91523, -43.9919, -44.0711, -44.14968, 
        -44.22544, -44.29608, -44.35999, -44.41608, -44.46345, -44.5007, 
        -44.52729, -44.54238, -44.54534, -44.53558, -44.51366, -44.48051, 
        -44.43837, -44.39027, -44.33996, -44.29133, -44.24734, -44.20937, 
        -44.17687,
  -39.00856, -39.02607, -39.04051, -39.05206, -39.0595, -39.06514, 
        -39.0687, -39.06982, -39.06784, -39.06338, -39.05779, -39.05218, 
        -39.04747, -39.04367, -39.04212, -39.04368, -39.04929, -39.06069, 
        -39.07806, -39.1038, -39.13753, -39.1799, -39.23074, -39.2905, 
        -39.36121, -39.44308, -39.53796, -39.64928, -39.77941, -39.9292, 
        -40.10095, -40.29494, -40.50927, -40.74142, -40.985, -41.2356, 
        -41.4854, -41.72819, -41.95877, -42.17205, -42.36608, -42.53875, 
        -42.69024, -42.82113, -42.9318, -43.02375, -43.09684, -43.15126, 
        -43.18773, -43.20443, -43.20425, -43.18538, -43.14795, -43.0938, 
        -43.02132, -42.93394, -42.83402, -42.72399, -42.60674, -42.48742, 
        -42.36867, -42.25276, -42.14467, -42.04809, -41.96759, -41.90379, 
        -41.856, -41.82714, -41.81739, -41.81824, -41.83172, -41.8563, 
        -41.88867, -41.92604, -41.96616, -42.00445, -42.03836, -42.06507, 
        -42.08294, -42.09197, -42.09157, -42.08323, -42.06886, -42.04726, 
        -42.0205, -41.98647, -41.94401, -41.89053, -41.82469, -41.74551, 
        -41.65401, -41.55278, -41.44556, -41.33401, -41.22209, -41.11225, 
        -41.00653, -40.90685, -40.81414, -40.72897, -40.65023, -40.57683, 
        -40.50626, -40.43953, -40.37309, -40.30554, -40.23669, -40.16761, 
        -40.10054, -40.03491, -39.97453, -39.91739, -39.86024, -39.80666, 
        -39.76341, -39.72731, -39.6962, -39.66912, -39.64442, -39.61934, 
        -39.5962, -39.57822, -39.55905, -39.53786, -39.51495, -39.49158, 
        -39.48368, -39.47236, -39.45504, -39.43533, -39.40652, -39.38414, 
        -39.36284, -39.33618, -39.31184, -39.28835, -39.27454, -39.269, 
        -39.25452, -39.24433, -39.24771, -39.24429, -39.23885, -39.23256, 
        -39.22592, -39.2226, -39.21053, -39.19764, -39.17738, -39.15265, 
        -39.11913, -39.07924, -39.03988, -39.00537, -38.97881, -38.94512, 
        -38.90543, -38.87092, -38.82983, -38.77827, -38.7243, -38.68391, 
        -38.6409, -38.61828, -38.60169, -38.5742, -38.53905, -38.49798, 
        -38.47532, -38.45152, -38.42684, -38.4302, -38.43213, -38.47701, 
        -38.53052, -38.59553, -38.68635, -38.77818, -38.86388, -38.93222, 
        -39.02106, -39.12089, -39.24423, -39.36724, -39.49972, -39.64027, 
        -39.76877, -39.89835, -40.02814, -40.16149, -40.29449, -40.42542, 
        -40.55192, -40.66928, -40.79028, -40.91219, -41.03398, -41.15264, 
        -41.2661, -41.36749, -41.45649, -41.53247, -41.59799, -41.65584, 
        -41.70861, -41.76226, -41.81868, -41.87761, -41.93949, -42.00528, 
        -42.07288, -42.14197, -42.2139, -42.29082, -42.36897, -42.45011, 
        -42.53428, -42.62221, -42.71316, -42.80696, -42.9049, -43.00532, 
        -43.10645, -43.20743, -43.30914, -43.41032, -43.50994, -43.60645, 
        -43.69968, -43.79, -43.87811, -43.9643, -44.0494, -44.1342, -44.2176, 
        -44.2977, -44.37241, -44.44064, -44.50128, -44.55332, -44.59666, 
        -44.63095, -44.65675, -44.67465, -44.68394, -44.68557, -44.67977, 
        -44.66792, -44.65042, -44.62822, -44.602, -44.57265, -44.54134, 
        -44.50861, -44.47741, -44.44701, -44.41655, -44.38441, -44.3488, 
        -44.30651, -44.25583, -44.19498, -44.12484, -44.048, -43.96679, 
        -43.88507, -43.80674, -43.73648, -43.67747, -43.63182, -43.60119, 
        -43.58519, -43.58307, -43.59429, -43.61924, -43.65601, -43.7039, 
        -43.76338, -43.83292, -43.90889, -43.98804, -44.06787, -44.14518, 
        -44.21732, -44.28236, -44.33937, -44.38716, -44.42482, -44.45207, 
        -44.46873, -44.47434, -44.46898, -44.45194, -44.42521, -44.38884, 
        -44.34566, -44.29844, -44.2496, -44.20386, -44.16222, -44.125,
  -39.07465, -39.09378, -39.1101, -39.12374, -39.13437, -39.14228, 
        -39.14807, -39.15081, -39.15033, -39.14732, -39.14326, -39.13953, 
        -39.1361, -39.1326, -39.13108, -39.13235, -39.13732, -39.14816, 
        -39.16619, -39.19201, -39.22564, -39.26795, -39.31928, -39.3792, 
        -39.44979, -39.53119, -39.625, -39.7351, -39.86109, -40.00822, 
        -40.17619, -40.3646, -40.5723, -40.79681, -41.03365, -41.27662, 
        -41.51969, -41.75723, -41.98431, -42.19588, -42.38916, -42.56202, 
        -42.71424, -42.84695, -42.95827, -43.05096, -43.12556, -43.18138, 
        -43.21943, -43.23879, -43.24072, -43.22496, -43.19164, -43.14164, 
        -43.07438, -42.99243, -42.89816, -42.79333, -42.68135, -42.56732, 
        -42.45166, -42.34004, -42.23511, -42.14023, -42.05894, -41.99312, 
        -41.94104, -41.90582, -41.88684, -41.87941, -41.88424, -41.90038, 
        -41.9246, -41.95481, -41.9887, -42.02282, -42.05435, -42.0788, 
        -42.09622, -42.10495, -42.10392, -42.09464, -42.07883, -42.057, 
        -42.02932, -41.99558, -41.9545, -41.90353, -41.84062, -41.76536, 
        -41.6782, -41.58094, -41.47617, -41.36678, -41.25435, -41.14064, 
        -41.03026, -40.92482, -40.82555, -40.73339, -40.64811, -40.56908, 
        -40.49577, -40.42656, -40.35919, -40.29177, -40.22372, -40.15586, 
        -40.09068, -40.02874, -39.97099, -39.91548, -39.86308, -39.81257, 
        -39.77162, -39.73869, -39.70983, -39.6869, -39.66545, -39.64745, 
        -39.63108, -39.61845, -39.60523, -39.59449, -39.57813, -39.56292, 
        -39.55283, -39.54453, -39.5357, -39.52395, -39.50733, -39.48642, 
        -39.47651, -39.45437, -39.43812, -39.41702, -39.4009, -39.37734, 
        -39.35824, -39.35724, -39.36399, -39.3659, -39.36729, -39.36552, 
        -39.35841, -39.34586, -39.33111, -39.31703, -39.29588, -39.26521, 
        -39.23172, -39.19373, -39.15801, -39.11816, -39.08155, -39.04337, 
        -38.99779, -38.95572, -38.90297, -38.84563, -38.80249, -38.76427, 
        -38.73022, -38.71815, -38.70052, -38.67558, -38.6466, -38.61528, 
        -38.58149, -38.55359, -38.54208, -38.53392, -38.55554, -38.6052, 
        -38.64835, -38.68386, -38.76685, -38.84751, -38.95469, -39.03479, 
        -39.11056, -39.18872, -39.31018, -39.43505, -39.55104, -39.68018, 
        -39.81004, -39.94723, -40.09071, -40.25055, -40.40339, -40.5467, 
        -40.67915, -40.79905, -40.92371, -41.04884, -41.17321, -41.29436, 
        -41.4086, -41.51159, -41.60252, -41.68095, -41.74872, -41.81027, 
        -41.8673, -41.92424, -41.98607, -42.05072, -42.11825, -42.18777, 
        -42.2597, -42.33304, -42.40833, -42.48729, -42.5685, -42.65304, 
        -42.74177, -42.8348, -42.93215, -43.03334, -43.13749, -43.24278, 
        -43.34779, -43.45155, -43.55373, -43.65353, -43.75027, -43.84296, 
        -43.93148, -44.01649, -44.09853, -44.17834, -44.25713, -44.33551, 
        -44.41264, -44.48686, -44.55598, -44.61932, -44.67538, -44.72271, 
        -44.76097, -44.79123, -44.81312, -44.82698, -44.83152, -44.82924, 
        -44.81984, -44.80333, -44.78014, -44.75259, -44.72075, -44.68418, 
        -44.64573, -44.60543, -44.56491, -44.52353, -44.48072, -44.43504, 
        -44.3842, -44.32611, -44.25959, -44.1836, -44.10004, -44.01177, 
        -43.92169, -43.83319, -43.75042, -43.67769, -43.61683, -43.56885, 
        -43.53582, -43.51624, -43.50961, -43.51494, -43.53207, -43.56246, 
        -43.60695, -43.66133, -43.72823, -43.80372, -43.88327, -43.96497, 
        -44.04447, -44.11841, -44.18521, -44.24335, -44.29193, -44.33032, 
        -44.35882, -44.37715, -44.38548, -44.38322, -44.37146, -44.34917, 
        -44.31783, -44.27826, -44.2329, -44.18462, -44.13683, -44.09137, 
        -44.04969,
  -39.15796, -39.17861, -39.19626, -39.21059, -39.22255, -39.23223, 
        -39.23878, -39.24266, -39.24211, -39.24041, -39.23793, -39.23534, 
        -39.23251, -39.23109, -39.23027, -39.23111, -39.23568, -39.2464, 
        -39.26417, -39.29042, -39.32497, -39.36788, -39.41992, -39.47975, 
        -39.5508, -39.63235, -39.72718, -39.83559, -39.96207, -40.10725, 
        -40.27131, -40.45456, -40.65573, -40.87134, -41.0977, -41.33027, 
        -41.5639, -41.7933, -42.0132, -42.2207, -42.41096, -42.5827, 
        -42.73483, -42.86788, -42.98073, -43.07396, -43.14926, -43.2064, 
        -43.24575, -43.26734, -43.27171, -43.25972, -43.23119, -43.18676, 
        -43.12607, -43.05024, -42.96327, -42.86582, -42.76099, -42.65361, 
        -42.5451, -42.43898, -42.33839, -42.24567, -42.16483, -42.0971, 
        -42.04136, -41.99958, -41.97171, -41.95549, -41.95085, -41.95593, 
        -41.97081, -41.99236, -42.01815, -42.04678, -42.07442, -42.09779, 
        -42.11406, -42.12209, -42.12029, -42.11003, -42.09304, -42.06991, 
        -42.04199, -42.00868, -41.96887, -41.92043, -41.86137, -41.79013, 
        -41.70816, -41.61673, -41.51722, -41.4109, -41.29808, -41.18362, 
        -41.06931, -40.95809, -40.8521, -40.7533, -40.66091, -40.57584, 
        -40.49804, -40.4262, -40.35796, -40.29122, -40.22437, -40.15772, 
        -40.093, -40.03358, -39.97723, -39.92451, -39.87551, -39.82674, 
        -39.78996, -39.76126, -39.73953, -39.72129, -39.70369, -39.69012, 
        -39.6779, -39.6692, -39.66056, -39.65652, -39.64916, -39.64051, 
        -39.63122, -39.62547, -39.61433, -39.60813, -39.60467, -39.59549, 
        -39.59557, -39.58801, -39.57126, -39.54859, -39.53167, -39.51043, 
        -39.48911, -39.48016, -39.48297, -39.49336, -39.49591, -39.49576, 
        -39.49112, -39.47727, -39.46327, -39.44231, -39.41675, -39.38566, 
        -39.35166, -39.31821, -39.28242, -39.24347, -39.20086, -39.1566, 
        -39.10649, -39.06052, -39.00435, -38.95159, -38.91288, -38.8758, 
        -38.84872, -38.82969, -38.807, -38.77962, -38.74813, -38.71832, 
        -38.68966, -38.66871, -38.66309, -38.67116, -38.68716, -38.7337, 
        -38.75019, -38.79697, -38.88627, -38.96996, -39.05874, -39.143, 
        -39.21569, -39.29921, -39.3946, -39.5128, -39.65025, -39.78098, 
        -39.91731, -40.04778, -40.20657, -40.37411, -40.53466, -40.681, 
        -40.8153, -40.93777, -41.06441, -41.19086, -41.31525, -41.43576, 
        -41.54931, -41.65089, -41.74242, -41.82231, -41.89228, -41.95716, 
        -42.01878, -42.08143, -42.14847, -42.21933, -42.29268, -42.36944, 
        -42.44763, -42.52582, -42.60572, -42.6884, -42.77304, -42.86084, 
        -42.95288, -43.0493, -43.15015, -43.25435, -43.36169, -43.4693, 
        -43.57539, -43.67924, -43.78056, -43.87812, -43.97192, -44.06055, 
        -44.14453, -44.2233, -44.29978, -44.37369, -44.44643, -44.51875, 
        -44.58943, -44.65749, -44.7212, -44.77892, -44.82926, -44.87181, 
        -44.90627, -44.93189, -44.9481, -44.95638, -44.95602, -44.94836, 
        -44.93386, -44.9123, -44.88403, -44.85006, -44.81144, -44.76791, 
        -44.72121, -44.67217, -44.62156, -44.56953, -44.51513, -44.45625, 
        -44.39158, -44.31937, -44.23898, -44.15042, -44.05587, -43.95833, 
        -43.86063, -43.76589, -43.6793, -43.60466, -43.54194, -43.49224, 
        -43.4567, -43.433, -43.42036, -43.41922, -43.42942, -43.45384, 
        -43.49138, -43.54382, -43.60834, -43.68371, -43.76467, -43.84811, 
        -43.92941, -44.00528, -44.0735, -44.13279, -44.18233, -44.22156, 
        -44.25098, -44.27076, -44.2808, -44.28138, -44.27269, -44.25386, 
        -44.22511, -44.18724, -44.1419, -44.09214, -44.04128, -43.99143, 
        -43.94553,
  -39.25554, -39.2773, -39.29503, -39.30912, -39.32126, -39.33151, 
        -39.33867, -39.34286, -39.34452, -39.34414, -39.3429, -39.34173, 
        -39.33984, -39.33857, -39.33843, -39.33957, -39.34438, -39.35524, 
        -39.37214, -39.39857, -39.43355, -39.47727, -39.52989, -39.5916, 
        -39.66356, -39.7459, -39.84134, -39.95048, -40.07621, -40.21955, 
        -40.38057, -40.55872, -40.75204, -40.95727, -41.17265, -41.39324, 
        -41.61538, -41.835, -42.04782, -42.2489, -42.43519, -42.60424, 
        -42.75509, -42.88691, -42.99931, -43.09321, -43.16856, -43.22621, 
        -43.26698, -43.28962, -43.29675, -43.28838, -43.26461, -43.22681, 
        -43.17333, -43.1066, -43.02802, -42.93948, -42.84312, -42.74322, 
        -42.64265, -42.54339, -42.44806, -42.35909, -42.27971, -42.21, 
        -42.15112, -42.10324, -42.06761, -42.04215, -42.02708, -42.02258, 
        -42.02653, -42.03792, -42.05568, -42.07767, -42.09993, -42.1194, 
        -42.1335, -42.14032, -42.13817, -42.12694, -42.10892, -42.08395, 
        -42.05539, -42.02217, -41.98388, -41.93787, -41.88316, -41.81835, 
        -41.74323, -41.65913, -41.56476, -41.4625, -41.35383, -41.23874, 
        -41.12126, -41.00512, -40.89281, -40.78599, -40.6866, -40.59439, 
        -40.51132, -40.43674, -40.36716, -40.30152, -40.23643, -40.17109, 
        -40.10714, -40.04753, -39.99532, -39.94292, -39.89032, -39.83637, 
        -39.8097, -39.78917, -39.77463, -39.75922, -39.74697, -39.73714, 
        -39.72889, -39.72222, -39.71732, -39.71796, -39.71907, -39.71716, 
        -39.71305, -39.70899, -39.6943, -39.69461, -39.70158, -39.70782, 
        -39.71902, -39.71628, -39.70528, -39.69062, -39.6751, -39.65097, 
        -39.62518, -39.60954, -39.61261, -39.61716, -39.62221, -39.62279, 
        -39.61789, -39.60626, -39.58899, -39.56384, -39.53194, -39.49976, 
        -39.46786, -39.43758, -39.40354, -39.36685, -39.32373, -39.27459, 
        -39.22564, -39.17685, -39.12052, -39.07438, -39.03109, -38.99238, 
        -38.96602, -38.9452, -38.91611, -38.88736, -38.86044, -38.8368, 
        -38.81736, -38.80456, -38.806, -38.80453, -38.83343, -38.86936, 
        -38.90514, -38.94543, -39.02099, -39.09766, -39.17638, -39.26125, 
        -39.33968, -39.41344, -39.50792, -39.60509, -39.74234, -39.89198, 
        -40.04431, -40.20147, -40.36829, -40.52831, -40.68234, -40.82597, 
        -40.96042, -41.08396, -41.21042, -41.33487, -41.45599, -41.57204, 
        -41.6813, -41.7811, -41.87076, -41.95053, -42.02248, -42.09102, 
        -42.1574, -42.22625, -42.2991, -42.37664, -42.45745, -42.54151, 
        -42.62653, -42.71172, -42.79766, -42.88456, -42.97271, -43.06371, 
        -43.15786, -43.25576, -43.35687, -43.46199, -43.56916, -43.67563, 
        -43.78085, -43.8829, -43.98137, -44.07643, -44.16632, -44.25091, 
        -44.33128, -44.4066, -44.47813, -44.54688, -44.61414, -44.68066, 
        -44.74527, -44.80736, -44.86499, -44.91644, -44.96132, -44.99853, 
        -45.0267, -45.04567, -45.05622, -45.0584, -45.05256, -45.03959, 
        -45.01934, -44.99206, -44.95829, -44.91772, -44.87188, -44.82084, 
        -44.76451, -44.70709, -44.64687, -44.58489, -44.51927, -44.44888, 
        -44.37228, -44.28817, -44.19633, -44.09717, -43.99351, -43.88826, 
        -43.78472, -43.6867, -43.59661, -43.51934, -43.45472, -43.40368, 
        -43.36452, -43.33655, -43.31898, -43.31219, -43.31693, -43.33541, 
        -43.36869, -43.41787, -43.48137, -43.55598, -43.63762, -43.72174, 
        -43.80416, -43.88119, -43.95048, -44.01036, -44.06001, -44.09965, 
        -44.12951, -44.14959, -44.16018, -44.1617, -44.15398, -44.13624, 
        -44.10802, -44.06853, -44.02162, -43.96938, -43.91416, -43.86022, 
        -43.81045,
  -39.36201, -39.38334, -39.40181, -39.41693, -39.42976, -39.4399, 
        -39.44759, -39.45246, -39.45509, -39.45628, -39.45707, -39.45721, 
        -39.45707, -39.4557, -39.456, -39.45783, -39.46349, -39.47447, 
        -39.49251, -39.51886, -39.55383, -39.59762, -39.6505, -39.71295, 
        -39.78571, -39.86938, -39.96539, -40.07496, -40.19893, -40.34021, 
        -40.49767, -40.66966, -40.85542, -41.05182, -41.25556, -41.46432, 
        -41.67463, -41.8836, -42.08739, -42.28131, -42.46209, -42.62725, 
        -42.77529, -42.90417, -43.01545, -43.10844, -43.18348, -43.24141, 
        -43.28309, -43.30864, -43.31845, -43.31346, -43.29499, -43.26279, 
        -43.21714, -43.15866, -43.0889, -43.00921, -42.92215, -42.83088, 
        -42.73755, -42.64525, -42.55603, -42.47155, -42.39448, -42.32545, 
        -42.26451, -42.21227, -42.1699, -42.13596, -42.11088, -42.09509, 
        -42.08933, -42.09011, -42.0987, -42.11229, -42.12777, -42.14165, 
        -42.15259, -42.15782, -42.15479, -42.14361, -42.12484, -42.10034, 
        -42.07112, -42.03761, -41.9999, -41.95618, -41.90569, -41.84669, 
        -41.77912, -41.70231, -41.61599, -41.51952, -41.41452, -41.30037, 
        -41.18222, -41.06284, -40.94451, -40.83112, -40.72439, -40.62669, 
        -40.53815, -40.46017, -40.38968, -40.32461, -40.26207, -40.19939, 
        -40.13849, -40.08228, -40.03149, -39.97726, -39.92955, -39.88812, 
        -39.86275, -39.84387, -39.82656, -39.81291, -39.80597, -39.79874, 
        -39.79396, -39.78844, -39.78626, -39.78825, -39.79078, -39.80154, 
        -39.8039, -39.79462, -39.79015, -39.79798, -39.81348, -39.83228, 
        -39.84501, -39.84938, -39.8437, -39.83091, -39.81591, -39.79544, 
        -39.7709, -39.75572, -39.75409, -39.75352, -39.75074, -39.74767, 
        -39.73996, -39.72804, -39.70853, -39.68187, -39.64812, -39.61478, 
        -39.58206, -39.55035, -39.51539, -39.47921, -39.43628, -39.38991, 
        -39.34087, -39.29366, -39.23901, -39.19288, -39.15062, -39.11399, 
        -39.0816, -39.05844, -39.02924, -39.00044, -38.97669, -38.95891, 
        -38.94938, -38.94447, -38.94753, -38.95587, -38.97969, -39.00999, 
        -39.05068, -39.10464, -39.1657, -39.23547, -39.31009, -39.38965, 
        -39.46937, -39.55117, -39.65005, -39.74452, -39.87366, -40.01878, 
        -40.18959, -40.3529, -40.52388, -40.68441, -40.83468, -40.97619, 
        -41.11036, -41.23316, -41.35697, -41.47681, -41.59161, -41.70063, 
        -41.80212, -41.89637, -41.98201, -42.0598, -42.13224, -42.20445, 
        -42.27604, -42.35132, -42.43117, -42.51575, -42.60337, -42.69633, 
        -42.78928, -42.88126, -42.9742, -43.06614, -43.15841, -43.25289, 
        -43.34857, -43.44661, -43.54825, -43.65162, -43.7557, -43.8588, 
        -43.96045, -44.05836, -44.15395, -44.24563, -44.33199, -44.41299, 
        -44.48916, -44.56088, -44.62884, -44.69281, -44.75479, -44.81575, 
        -44.8744, -44.93039, -44.98152, -45.02695, -45.06546, -45.09513, 
        -45.11699, -45.12915, -45.13345, -45.12947, -45.11704, -45.09914, 
        -45.07297, -45.03962, -44.99992, -44.9525, -44.89989, -44.84076, 
        -44.77689, -44.71146, -44.64307, -44.57174, -44.49636, -44.41615, 
        -44.32986, -44.2365, -44.13583, -44.02851, -43.91779, -43.80632, 
        -43.69754, -43.59525, -43.50257, -43.42266, -43.35635, -43.30305, 
        -43.26184, -43.23074, -43.20932, -43.19831, -43.19902, -43.21379, 
        -43.24439, -43.29145, -43.35349, -43.42662, -43.50753, -43.59117, 
        -43.6735, -43.75013, -43.81894, -43.87795, -43.92659, -43.96535, 
        -43.99453, -44.0136, -44.0232, -44.02359, -44.01469, -43.99559, 
        -43.96523, -43.92421, -43.87378, -43.81702, -43.75758, -43.69976, 
        -43.64682,
  -39.47514, -39.49621, -39.51435, -39.53, -39.54314, -39.5539, 
        -39.56239, -39.56859, -39.57236, -39.57554, -39.57836, -39.58033, 
        -39.58211, -39.58371, -39.58514, -39.58814, -39.59433, -39.60587, 
        -39.62405, -39.65005, -39.68445, -39.72757, -39.78024, -39.842, 
        -39.91519, -39.99955, -40.09601, -40.20534, -40.32891, -40.46743, 
        -40.62024, -40.78622, -40.96395, -41.15073, -41.34385, -41.54116, 
        -41.74038, -41.93848, -42.13139, -42.31746, -42.49183, -42.65199, 
        -42.7962, -42.92311, -43.03221, -43.12363, -43.19794, -43.25567, 
        -43.29793, -43.32495, -43.33735, -43.33555, -43.32117, -43.29469, 
        -43.25452, -43.20395, -43.14275, -43.07211, -42.99364, -42.91099, 
        -42.82648, -42.74133, -42.65836, -42.57885, -42.50486, -42.43698, 
        -42.37545, -42.32075, -42.27286, -42.23198, -42.19818, -42.17303, 
        -42.15586, -42.14672, -42.14507, -42.14949, -42.15769, -42.16641, 
        -42.17329, -42.17614, -42.17229, -42.16084, -42.14253, -42.11798, 
        -42.08793, -42.05393, -42.01613, -41.97471, -41.92847, -41.87442, 
        -41.81368, -41.74515, -41.66722, -41.57863, -41.47879, -41.36984, 
        -41.2526, -41.13143, -41.00956, -40.89052, -40.77739, -40.67343, 
        -40.57936, -40.49773, -40.42603, -40.36168, -40.30168, -40.24286, 
        -40.18877, -40.13852, -40.08979, -40.0401, -40.00024, -39.96544, 
        -39.94085, -39.92742, -39.91401, -39.90251, -39.89536, -39.89169, 
        -39.88852, -39.88423, -39.87625, -39.87682, -39.88928, -39.90049, 
        -39.90336, -39.90023, -39.90874, -39.92381, -39.94263, -39.96437, 
        -39.9814, -39.99047, -39.98626, -39.97553, -39.96014, -39.94094, 
        -39.9229, -39.90827, -39.89616, -39.8872, -39.88012, -39.87211, 
        -39.86193, -39.84742, -39.82721, -39.80003, -39.76685, -39.73113, 
        -39.69572, -39.66073, -39.6233, -39.58413, -39.53976, -39.4951, 
        -39.44957, -39.40501, -39.35297, -39.30792, -39.26519, -39.22844, 
        -39.19642, -39.17303, -39.14189, -39.11399, -39.09092, -39.07711, 
        -39.07291, -39.07159, -39.07846, -39.09356, -39.11711, -39.1487, 
        -39.19565, -39.2503, -39.31223, -39.38087, -39.45493, -39.53436, 
        -39.61993, -39.71091, -39.81388, -39.92645, -40.05502, -40.19554, 
        -40.35241, -40.51472, -40.68031, -40.83596, -40.98449, -41.12502, 
        -41.2574, -41.37773, -41.49654, -41.60919, -41.71524, -41.81443, 
        -41.90519, -41.99084, -42.07042, -42.14536, -42.21871, -42.29375, 
        -42.37085, -42.45316, -42.54095, -42.6344, -42.7316, -42.8317, 
        -42.93177, -43.03232, -43.13298, -43.22979, -43.32711, -43.42375, 
        -43.5214, -43.61878, -43.71737, -43.81699, -43.91648, -44.01372, 
        -44.1095, -44.20298, -44.29393, -44.38106, -44.46388, -44.54144, 
        -44.61312, -44.68162, -44.74554, -44.80614, -44.86356, -44.91837, 
        -44.97085, -45.02026, -45.06511, -45.10386, -45.13588, -45.16037, 
        -45.17548, -45.18138, -45.17873, -45.16856, -45.1504, -45.12555, 
        -45.09491, -45.05592, -45.00934, -44.95498, -44.89451, -44.82855, 
        -44.75858, -44.68478, -44.60829, -44.52893, -44.44584, -44.35771, 
        -44.26407, -44.16409, -44.05724, -43.94471, -43.82891, -43.71192, 
        -43.59719, -43.49039, -43.39474, -43.31238, -43.24413, -43.18956, 
        -43.14673, -43.11451, -43.09154, -43.07962, -43.07831, -43.092, 
        -43.12185, -43.16843, -43.22871, -43.30089, -43.38054, -43.4627, 
        -43.54314, -43.61736, -43.68349, -43.73994, -43.786, -43.82188, 
        -43.84836, -43.86517, -43.87221, -43.86991, -43.85776, -43.83528, 
        -43.80053, -43.7546, -43.69946, -43.63759, -43.57367, -43.51218, 
        -43.45741,
  -39.59075, -39.61138, -39.62949, -39.64471, -39.65854, -39.67049, 
        -39.6808, -39.68927, -39.69638, -39.70229, -39.70774, -39.71235, 
        -39.71651, -39.72012, -39.72356, -39.7281, -39.73544, -39.74741, 
        -39.76474, -39.79024, -39.82354, -39.8658, -39.9178, -39.98004, 
        -40.05306, -40.1372, -40.23313, -40.34159, -40.46301, -40.59753, 
        -40.74559, -40.90578, -41.07556, -41.2518, -41.43511, -41.62194, 
        -41.81048, -41.99818, -42.18246, -42.36011, -42.52735, -42.68158, 
        -42.82078, -42.94389, -43.04994, -43.13914, -43.21201, -43.26938, 
        -43.31155, -43.3389, -43.35315, -43.35428, -43.34359, -43.32143, 
        -43.28857, -43.24462, -43.19113, -43.12848, -43.05833, -42.98332, 
        -42.90625, -42.82858, -42.75162, -42.67764, -42.60819, -42.54172, 
        -42.48082, -42.42494, -42.37379, -42.32751, -42.28799, -42.25485, 
        -42.22868, -42.20955, -42.19777, -42.19221, -42.19141, -42.19304, 
        -42.19493, -42.19501, -42.19011, -42.17886, -42.16002, -42.13591, 
        -42.10616, -42.07207, -42.03466, -41.99441, -41.95156, -41.90382, 
        -41.8501, -41.78969, -41.72063, -41.64049, -41.54848, -41.44503, 
        -41.33144, -41.21101, -41.08735, -40.96474, -40.84715, -40.73654, 
        -40.63797, -40.55271, -40.47871, -40.41426, -40.35683, -40.30403, 
        -40.25486, -40.20962, -40.16789, -40.1267, -40.09146, -40.06228, 
        -40.04169, -40.02853, -40.01838, -40.0113, -40.00765, -40.00614, 
        -40.00364, -40.00143, -39.99648, -39.99977, -40.00832, -40.01915, 
        -40.03203, -40.04618, -40.06076, -40.07885, -40.0994, -40.12011, 
        -40.13541, -40.14271, -40.13982, -40.12967, -40.11404, -40.0953, 
        -40.07834, -40.05958, -40.04198, -40.02574, -40.01338, -40.00082, 
        -39.9865, -39.96969, -39.94797, -39.92097, -39.88728, -39.85226, 
        -39.81493, -39.77538, -39.7337, -39.69227, -39.64786, -39.60278, 
        -39.55845, -39.51702, -39.46993, -39.42642, -39.38606, -39.34878, 
        -39.31612, -39.2897, -39.25846, -39.23106, -39.2079, -39.19409, 
        -39.1911, -39.19271, -39.20319, -39.22305, -39.25268, -39.2903, 
        -39.34286, -39.40327, -39.46889, -39.53893, -39.6148, -39.69637, 
        -39.78399, -39.87813, -39.98186, -40.09828, -40.22536, -40.36518, 
        -40.51326, -40.66641, -40.82265, -40.97309, -41.11869, -41.25666, 
        -41.38608, -41.50433, -41.6167, -41.7214, -41.81755, -41.90595, 
        -41.98728, -42.06376, -42.13687, -42.209, -42.28317, -42.3619, 
        -42.44576, -42.53647, -42.63391, -42.7371, -42.84338, -42.95155, 
        -43.05867, -43.16644, -43.27305, -43.37661, -43.47668, -43.5757, 
        -43.67265, -43.7673, -43.86163, -43.95469, -44.04718, -44.13768, 
        -44.22609, -44.31287, -44.3975, -44.47972, -44.55852, -44.63273, 
        -44.70211, -44.76718, -44.8278, -44.88472, -44.93781, -44.98711, 
        -45.03348, -45.07583, -45.11447, -45.14715, -45.1724, -45.19006, 
        -45.19855, -45.19874, -45.18989, -45.17333, -45.14982, -45.11912, 
        -45.08204, -45.03632, -44.98396, -44.92329, -44.85577, -44.78181, 
        -44.70424, -44.62257, -44.53914, -44.45302, -44.36354, -44.26986, 
        -44.17113, -44.06729, -43.95706, -43.84202, -43.7234, -43.60241, 
        -43.48434, -43.37379, -43.27483, -43.19014, -43.11966, -43.06453, 
        -43.02178, -42.98923, -42.96727, -42.95659, -42.95823, -42.97315, 
        -43.0042, -43.05103, -43.11137, -43.18101, -43.25801, -43.33713, 
        -43.41407, -43.48389, -43.54509, -43.5966, -43.63765, -43.66883, 
        -43.69086, -43.70322, -43.70613, -43.6995, -43.68294, -43.65558, 
        -43.61453, -43.56327, -43.50254, -43.43575, -43.36775, -43.30369, 
        -43.24896,
  -39.70549, -39.72591, -39.74461, -39.76131, -39.77633, -39.79035, 
        -39.80283, -39.814, -39.82418, -39.83357, -39.84211, -39.85007, 
        -39.85705, -39.86219, -39.86833, -39.87443, -39.88343, -39.89635, 
        -39.91525, -39.94, -39.97229, -40.01352, -40.06414, -40.1255, 
        -40.19744, -40.28067, -40.37521, -40.48147, -40.59897, -40.72996, 
        -40.87269, -41.02606, -41.18805, -41.35644, -41.53024, -41.70755, 
        -41.88591, -42.06381, -42.23874, -42.40765, -42.56716, -42.71471, 
        -42.84847, -42.96584, -43.06829, -43.1548, -43.22603, -43.28248, 
        -43.32471, -43.3536, -43.36933, -43.37264, -43.36501, -43.34697, 
        -43.31886, -43.28083, -43.23376, -43.17822, -43.11535, -43.04655, 
        -42.97629, -42.90525, -42.83466, -42.76689, -42.702, -42.64069, 
        -42.58209, -42.52638, -42.4744, -42.42535, -42.38029, -42.3401, 
        -42.30566, -42.27717, -42.25516, -42.23924, -42.22795, -42.22163, 
        -42.21776, -42.21461, -42.20865, -42.198, -42.18131, -42.15832, 
        -42.12978, -42.09629, -42.0594, -42.02047, -41.97935, -41.93631, 
        -41.89025, -41.83723, -41.77677, -41.70621, -41.62203, -41.52582, 
        -41.41837, -41.30144, -41.17862, -41.05545, -40.93543, -40.8226, 
        -40.72013, -40.63115, -40.55455, -40.48918, -40.43249, -40.38202, 
        -40.33748, -40.29651, -40.25969, -40.22587, -40.19624, -40.16949, 
        -40.15221, -40.14021, -40.13308, -40.12984, -40.12915, -40.13084, 
        -40.13341, -40.13605, -40.13821, -40.14465, -40.15232, -40.16709, 
        -40.18261, -40.20046, -40.21922, -40.24071, -40.26389, -40.28444, 
        -40.2994, -40.30602, -40.30354, -40.29403, -40.27795, -40.2575, 
        -40.23747, -40.21496, -40.19226, -40.17131, -40.15314, -40.13442, 
        -40.11588, -40.09547, -40.07172, -40.04378, -40.00935, -39.97318, 
        -39.93393, -39.89206, -39.84806, -39.80408, -39.75737, -39.71167, 
        -39.66702, -39.62492, -39.57952, -39.53856, -39.5006, -39.46519, 
        -39.43384, -39.40716, -39.37925, -39.35328, -39.33266, -39.31916, 
        -39.31733, -39.32119, -39.33514, -39.35981, -39.39572, -39.44006, 
        -39.49715, -39.56205, -39.63214, -39.70601, -39.78373, -39.86647, 
        -39.9536, -40.04865, -40.15231, -40.26628, -40.39036, -40.52478, 
        -40.6674, -40.81525, -40.96613, -41.11336, -41.25451, -41.3876, 
        -41.5111, -41.62287, -41.7261, -41.81919, -41.90329, -41.97905, 
        -42.04858, -42.11501, -42.18157, -42.25161, -42.32752, -42.41238, 
        -42.50486, -42.60534, -42.71264, -42.8242, -42.9391, -43.05402, 
        -43.16939, -43.28292, -43.39397, -43.50066, -43.60337, -43.70202, 
        -43.79751, -43.88938, -43.97802, -44.06366, -44.14684, -44.22815, 
        -44.30828, -44.38729, -44.46511, -44.54139, -44.61549, -44.6862, 
        -44.75245, -44.8142, -44.87117, -44.92413, -44.9728, -45.01682, 
        -45.05733, -45.09297, -45.12453, -45.15139, -45.17081, -45.18097, 
        -45.18348, -45.17772, -45.16341, -45.14109, -45.11171, -45.07521, 
        -45.03126, -44.97966, -44.9206, -44.85372, -44.77895, -44.69936, 
        -44.61563, -44.52828, -44.43882, -44.34706, -44.25292, -44.15578, 
        -44.0543, -43.94844, -43.83785, -43.7207, -43.60102, -43.47752, 
        -43.35694, -43.24278, -43.14059, -43.05229, -42.98017, -42.92338, 
        -42.88163, -42.85225, -42.83363, -42.82724, -42.83405, -42.8542, 
        -42.88905, -42.93577, -42.99556, -43.06475, -43.13873, -43.21331, 
        -43.28466, -43.34874, -43.40316, -43.44749, -43.48162, -43.50638, 
        -43.52203, -43.52868, -43.52647, -43.51479, -43.49315, -43.46017, 
        -43.41467, -43.35806, -43.29231, -43.22177, -43.15134, -43.0871, 
        -43.03331,
  -39.82113, -39.84163, -39.86087, -39.87841, -39.89473, -39.91069, 
        -39.92565, -39.94007, -39.95259, -39.96552, -39.9779, -39.98943, 
        -39.9995, -40.0092, -40.01762, -40.02673, -40.03822, -40.05254, 
        -40.07245, -40.09693, -40.12872, -40.16881, -40.21703, -40.27663, 
        -40.34706, -40.42865, -40.52116, -40.62484, -40.73982, -40.86606, 
        -41.00316, -41.14937, -41.30357, -41.46367, -41.62834, -41.79618, 
        -41.96509, -42.13356, -42.29827, -42.45847, -42.61003, -42.74998, 
        -42.87778, -42.99093, -43.08948, -43.17311, -43.24247, -43.29778, 
        -43.33952, -43.36868, -43.38538, -43.39045, -43.38512, -43.37037, 
        -43.34542, -43.3119, -43.2705, -43.2212, -43.16504, -43.10413, 
        -43.04037, -42.97594, -42.91191, -42.84966, -42.7905, -42.73351, 
        -42.67843, -42.62497, -42.57321, -42.5229, -42.47336, -42.42772, 
        -42.38582, -42.34845, -42.31625, -42.2903, -42.27031, -42.25592, 
        -42.24636, -42.2395, -42.23248, -42.22281, -42.20766, -42.18714, 
        -42.16069, -42.12911, -42.09354, -42.05607, -42.01632, -41.97693, 
        -41.93537, -41.88999, -41.83789, -41.77652, -41.70295, -41.61681, 
        -41.51708, -41.40666, -41.28842, -41.16738, -41.04767, -40.93375, 
        -40.82909, -40.7368, -40.65714, -40.58969, -40.53257, -40.48229, 
        -40.43945, -40.40201, -40.36938, -40.34015, -40.31549, -40.29405, 
        -40.27971, -40.2708, -40.26679, -40.26701, -40.26979, -40.27501, 
        -40.281, -40.28725, -40.29359, -40.30433, -40.31564, -40.32948, 
        -40.34637, -40.36549, -40.3866, -40.41047, -40.43414, -40.45493, 
        -40.47028, -40.47763, -40.47722, -40.46831, -40.45202, -40.43028, 
        -40.40785, -40.38113, -40.35417, -40.32841, -40.30411, -40.28047, 
        -40.2569, -40.23196, -40.20443, -40.17323, -40.13472, -40.09644, 
        -40.05552, -40.01228, -39.96668, -39.92128, -39.8736, -39.82625, 
        -39.7815, -39.73973, -39.69586, -39.65764, -39.6225, -39.58919, 
        -39.55929, -39.533, -39.50639, -39.48211, -39.46207, -39.44888, 
        -39.44768, -39.45299, -39.46946, -39.49705, -39.53802, -39.58833, 
        -39.65072, -39.72057, -39.79537, -39.87349, -39.95385, -40.03773, 
        -40.12532, -40.21832, -40.3184, -40.42746, -40.54585, -40.67405, 
        -40.81042, -40.95247, -41.09727, -41.23891, -41.37461, -41.50159, 
        -41.61753, -41.72034, -41.81301, -41.89436, -41.9652, -42.0271, 
        -42.08529, -42.14301, -42.20481, -42.27469, -42.35518, -42.44782, 
        -42.55102, -42.66285, -42.78074, -42.90261, -43.02579, -43.14807, 
        -43.2681, -43.38515, -43.49847, -43.60675, -43.70941, -43.80593, 
        -43.89695, -43.98301, -44.06396, -44.14058, -44.21317, -44.28363, 
        -44.35369, -44.42385, -44.49442, -44.56454, -44.63287, -44.69801, 
        -44.76109, -44.81988, -44.87329, -44.92188, -44.96592, -45.00497, 
        -45.03939, -45.06906, -45.09419, -45.11429, -45.12794, -45.13334, 
        -45.13004, -45.11843, -45.09896, -45.07124, -45.03625, -44.99365, 
        -44.94326, -44.8851, -44.81953, -44.74584, -44.66475, -44.57807, 
        -44.48804, -44.39534, -44.30084, -44.20474, -44.10725, -44.00797, 
        -43.90595, -43.80058, -43.68932, -43.57338, -43.45338, -43.32907, 
        -43.20745, -43.0905, -42.98586, -42.89676, -42.82331, -42.76604, 
        -42.72546, -42.69977, -42.68851, -42.69035, -42.70458, -42.73211, 
        -42.77233, -42.82364, -42.88459, -42.95239, -43.02319, -43.09276, 
        -43.15731, -43.21377, -43.26036, -43.29617, -43.32164, -43.33816, 
        -43.34588, -43.3458, -43.33756, -43.3204, -43.29327, -43.25493, 
        -43.20515, -43.14472, -43.07645, -43.00443, -42.93451, -42.8718, 
        -42.82107,
  -39.93671, -39.9574, -39.97676, -39.99412, -40.01214, -40.02976, 
        -40.04739, -40.0648, -40.08164, -40.09797, -40.11395, -40.12885, 
        -40.14272, -40.15543, -40.16788, -40.18053, -40.19465, -40.21128, 
        -40.2319, -40.25665, -40.28873, -40.32775, -40.37612, -40.43422, 
        -40.50317, -40.58269, -40.67264, -40.77308, -40.8839, -41.005, 
        -41.1358, -41.27488, -41.42002, -41.5718, -41.7279, -41.88662, 
        -42.04652, -42.20554, -42.3621, -42.51334, -42.65643, -42.78937, 
        -42.91044, -43.01831, -43.1126, -43.19341, -43.26041, -43.31419, 
        -43.35413, -43.3829, -43.40044, -43.40657, -43.40322, -43.39074, 
        -43.36993, -43.34094, -43.30465, -43.26111, -43.2113, -43.15705, 
        -43.09983, -43.04199, -42.98455, -42.92847, -42.87472, -42.82148, 
        -42.77061, -42.72018, -42.6697, -42.61925, -42.56917, -42.51906, 
        -42.47033, -42.42485, -42.38372, -42.34827, -42.31963, -42.29755, 
        -42.28217, -42.27222, -42.26428, -42.25515, -42.2418, -42.22424, 
        -42.20112, -42.17202, -42.1387, -42.103, -42.06618, -42.02974, 
        -41.99225, -41.95321, -41.90994, -41.85773, -41.79402, -41.71762, 
        -41.62813, -41.52623, -41.41583, -41.30007, -41.18263, -41.07011, 
        -40.96474, -40.87013, -40.78779, -40.71772, -40.65875, -40.60904, 
        -40.56733, -40.53163, -40.50111, -40.47515, -40.45392, -40.43656, 
        -40.42567, -40.42019, -40.41932, -40.42252, -40.42833, -40.43653, 
        -40.44461, -40.45393, -40.4634, -40.47617, -40.48849, -40.50296, 
        -40.52034, -40.54078, -40.56259, -40.58709, -40.6113, -40.63266, 
        -40.64885, -40.65741, -40.65806, -40.65015, -40.63416, -40.61174, 
        -40.58734, -40.55759, -40.52676, -40.49512, -40.46524, -40.43615, 
        -40.40723, -40.37735, -40.34529, -40.30929, -40.26835, -40.22754, 
        -40.18645, -40.142, -40.09492, -40.0486, -40.00055, -39.95344, 
        -39.9085, -39.86668, -39.8229, -39.78696, -39.75414, -39.7238, 
        -39.69541, -39.66945, -39.64359, -39.61983, -39.59969, -39.58601, 
        -39.58447, -39.59031, -39.60831, -39.63955, -39.68422, -39.73912, 
        -39.80622, -39.88086, -39.95994, -40.04146, -40.12365, -40.20705, 
        -40.2922, -40.38076, -40.47485, -40.5765, -40.68682, -40.80698, 
        -40.93562, -41.0704, -41.20761, -41.34329, -41.47199, -41.5916, 
        -41.69902, -41.79283, -41.87403, -41.94276, -42.00095, -42.0519, 
        -42.09999, -42.15178, -42.21193, -42.28487, -42.37282, -42.47578, 
        -42.59133, -42.71536, -42.8444, -42.97507, -43.10528, -43.23232, 
        -43.35538, -43.47384, -43.58703, -43.69378, -43.79298, -43.88548, 
        -43.96961, -44.04574, -44.11624, -44.18208, -44.24331, -44.30194, 
        -44.36087, -44.42141, -44.48375, -44.5471, -44.61004, -44.67117, 
        -44.7302, -44.78527, -44.83501, -44.87942, -44.9183, -44.95204, 
        -44.98067, -45.00439, -45.0232, -45.03673, -45.04438, -45.04414, 
        -45.03508, -45.01813, -44.99294, -44.96013, -44.92, -44.87039, 
        -44.8133, -44.74855, -44.67618, -44.59542, -44.506, -44.41333, 
        -44.31676, -44.21878, -44.12074, -44.021, -43.92162, -43.82167, 
        -43.72026, -43.61591, -43.50665, -43.39291, -43.27445, -43.15251, 
        -43.03134, -42.91607, -42.81119, -42.72139, -42.64934, -42.5944, 
        -42.55711, -42.53719, -42.53377, -42.54566, -42.57085, -42.60802, 
        -42.65597, -42.71268, -42.77571, -42.84291, -42.91018, -42.97404, 
        -43.03134, -43.0794, -43.11675, -43.14301, -43.159, -43.16616, 
        -43.1657, -43.15791, -43.14293, -43.11995, -43.08694, -43.0446, 
        -42.99219, -42.93043, -42.86246, -42.79256, -42.72571, -42.66695, 
        -42.62072,
  -40.05056, -40.07143, -40.09108, -40.11001, -40.12921, -40.14827, 
        -40.16838, -40.188, -40.20779, -40.22731, -40.24598, -40.26436, 
        -40.28149, -40.29848, -40.31503, -40.33162, -40.34952, -40.36945, 
        -40.39212, -40.41871, -40.45121, -40.49065, -40.53828, -40.59536, 
        -40.66255, -40.73975, -40.82706, -40.92297, -41.02943, -41.14501, 
        -41.26935, -41.40125, -41.53957, -41.68306, -41.83033, -41.98019, 
        -42.13093, -42.28075, -42.42798, -42.57028, -42.70528, -42.83061, 
        -42.94481, -43.04644, -43.13654, -43.21384, -43.27827, -43.33041, 
        -43.37003, -43.39819, -43.41584, -43.42286, -43.42075, -43.41021, 
        -43.39267, -43.36761, -43.33601, -43.2983, -43.25496, -43.20637, 
        -43.15615, -43.10501, -43.05398, -43.00407, -42.95544, -42.90789, 
        -42.86115, -42.81414, -42.76617, -42.71644, -42.66471, -42.612, 
        -42.55851, -42.50628, -42.45748, -42.41402, -42.37706, -42.34899, 
        -42.3287, -42.31558, -42.30627, -42.29784, -42.28783, -42.27411, 
        -42.25486, -42.2294, -42.19922, -42.16519, -42.13068, -42.09626, 
        -42.06286, -42.02906, -41.99231, -41.94844, -41.89396, -41.82808, 
        -41.74958, -41.6591, -41.55824, -41.45083, -41.34023, -41.23079, 
        -41.12727, -41.03195, -40.94731, -40.87509, -40.81369, -40.76287, 
        -40.72031, -40.68521, -40.65592, -40.63185, -40.61297, -40.59745, 
        -40.58908, -40.58623, -40.58805, -40.59371, -40.60173, -40.61229, 
        -40.62367, -40.63518, -40.64668, -40.66002, -40.67277, -40.68719, 
        -40.70401, -40.72358, -40.74474, -40.76861, -40.79258, -40.81417, 
        -40.83112, -40.83983, -40.84194, -40.83534, -40.8203, -40.79799, 
        -40.77238, -40.7406, -40.70644, -40.67167, -40.63707, -40.60265, 
        -40.56849, -40.53395, -40.49762, -40.45809, -40.41446, -40.37195, 
        -40.32952, -40.28373, -40.23608, -40.18938, -40.14178, -40.09442, 
        -40.05042, -40.00934, -39.96802, -39.93387, -39.90272, -39.87393, 
        -39.8465, -39.82152, -39.79583, -39.77166, -39.751, -39.73626, 
        -39.73317, -39.73833, -39.75653, -39.78892, -39.83544, -39.89316, 
        -39.96306, -40.04046, -40.12194, -40.20472, -40.28651, -40.36632, 
        -40.44656, -40.52816, -40.61351, -40.7054, -40.80579, -40.91606, 
        -41.03556, -41.16198, -41.29219, -41.42099, -41.54392, -41.65723, 
        -41.7559, -41.84087, -41.91047, -41.96727, -42.01361, -42.05492, 
        -42.09578, -42.14516, -42.20683, -42.28646, -42.38474, -42.49989, 
        -42.62831, -42.76484, -42.90382, -43.04207, -43.17714, -43.30656, 
        -43.43032, -43.54669, -43.65674, -43.75858, -43.85205, -43.93623, 
        -44.0107, -44.07775, -44.13616, -44.18917, -44.23801, -44.28481, 
        -44.33245, -44.38274, -44.43644, -44.49271, -44.54978, -44.60611, 
        -44.66037, -44.71104, -44.75673, -44.7966, -44.83048, -44.8583, 
        -44.8805, -44.89791, -44.91096, -44.91694, -44.91681, -44.91064, 
        -44.89644, -44.87431, -44.84338, -44.80574, -44.75989, -44.7036, 
        -44.63886, -44.5681, -44.48691, -44.39849, -44.30283, -44.20323, 
        -44.10159, -43.9986, -43.89648, -43.79534, -43.69534, -43.59658, 
        -43.49628, -43.39404, -43.28764, -43.17737, -43.06221, -42.94353, 
        -42.82694, -42.71545, -42.61429, -42.52766, -42.45872, -42.40867, 
        -42.37808, -42.36656, -42.37352, -42.39671, -42.43431, -42.4832, 
        -42.54018, -42.60333, -42.66907, -42.73589, -42.79992, -42.85777, 
        -42.9071, -42.94622, -42.97413, -42.99056, -42.99697, -42.99469, 
        -42.985, -42.96915, -42.94677, -42.91824, -42.88227, -42.83744, 
        -42.78484, -42.72469, -42.66044, -42.59545, -42.53459, -42.4822, 
        -42.4412,
  -40.16389, -40.18468, -40.20455, -40.22406, -40.24378, -40.26423, 
        -40.28548, -40.30607, -40.32787, -40.34976, -40.37129, -40.39302, 
        -40.41432, -40.43532, -40.45646, -40.47799, -40.50023, -40.524, 
        -40.54974, -40.57865, -40.61253, -40.65287, -40.69962, -40.75611, 
        -40.822, -40.89689, -40.98115, -41.07446, -41.17643, -41.28663, 
        -41.40464, -41.5295, -41.66011, -41.79543, -41.93388, -42.07462, 
        -42.21611, -42.35583, -42.49395, -42.62757, -42.75451, -42.87241, 
        -42.98013, -43.07692, -43.16219, -43.23566, -43.29728, -43.34734, 
        -43.38568, -43.41299, -43.43005, -43.43734, -43.43615, -43.42678, 
        -43.41204, -43.39121, -43.36453, -43.33279, -43.29619, -43.25575, 
        -43.21239, -43.16784, -43.12345, -43.07883, -43.03493, -42.99201, 
        -42.949, -42.9053, -42.85956, -42.81093, -42.75879, -42.70419, 
        -42.64741, -42.59095, -42.53687, -42.48779, -42.44655, -42.41408, 
        -42.39017, -42.37397, -42.36319, -42.35496, -42.34705, -42.33667, 
        -42.32159, -42.30059, -42.27319, -42.24281, -42.20871, -42.1768, 
        -42.14601, -42.11641, -42.08506, -42.04872, -42.00393, -41.9487, 
        -41.8819, -41.80324, -41.71383, -41.61601, -41.51328, -41.41028, 
        -41.31042, -41.21663, -41.1315, -41.05684, -40.99302, -40.94024, 
        -40.89659, -40.86079, -40.83148, -40.80871, -40.79087, -40.77785, 
        -40.7707, -40.76914, -40.77249, -40.77966, -40.78947, -40.80117, 
        -40.81393, -40.8267, -40.83893, -40.85163, -40.86372, -40.87689, 
        -40.89104, -40.90858, -40.92811, -40.95013, -40.97271, -40.99392, 
        -41.01118, -41.02223, -41.02571, -41.02073, -41.0069, -40.98513, 
        -40.95811, -40.92483, -40.88828, -40.85028, -40.81191, -40.77345, 
        -40.7352, -40.69694, -40.658, -40.61742, -40.57235, -40.52891, 
        -40.48527, -40.43953, -40.39242, -40.34591, -40.29935, -40.2547, 
        -40.2125, -40.17337, -40.13578, -40.10326, -40.07353, -40.04556, 
        -40.01845, -39.99253, -39.96592, -39.94045, -39.91796, -39.901, 
        -39.89398, -39.89693, -39.9134, -39.94359, -39.98957, -40.04805, 
        -40.11819, -40.19559, -40.2765, -40.35766, -40.43636, -40.51207, 
        -40.58506, -40.6573, -40.73187, -40.81229, -40.90106, -40.99995, 
        -41.10913, -41.22681, -41.34972, -41.4724, -41.58926, -41.69535, 
        -41.7877, -41.86356, -41.92361, -41.97023, -42.0072, -42.04019, 
        -42.077, -42.1263, -42.19418, -42.28344, -42.39431, -42.5228, 
        -42.66393, -42.81177, -42.96008, -43.10464, -43.24168, -43.37077, 
        -43.49105, -43.60361, -43.70699, -43.80015, -43.88445, -43.95745, 
        -44.02143, -44.07529, -44.12155, -44.16113, -44.19739, -44.23248, 
        -44.26922, -44.30973, -44.35447, -44.40356, -44.45377, -44.50502, 
        -44.55442, -44.59988, -44.6405, -44.6753, -44.70348, -44.72516, 
        -44.74072, -44.75077, -44.75603, -44.75522, -44.74798, -44.7352, 
        -44.71514, -44.68682, -44.65244, -44.60854, -44.55495, -44.49276, 
        -44.42222, -44.34185, -44.25404, -44.15822, -44.05626, -43.94989, 
        -43.84248, -43.73676, -43.63147, -43.52956, -43.43026, -43.33298, 
        -43.23507, -43.13564, -43.03329, -42.92672, -42.81582, -42.70306, 
        -42.5941, -42.49052, -42.39644, -42.31718, -42.25622, -42.21465, 
        -42.19389, -42.19326, -42.21259, -42.24974, -42.30075, -42.36223, 
        -42.4306, -42.50084, -42.5705, -42.63645, -42.69673, -42.74849, 
        -42.78978, -42.82003, -42.83862, -42.84571, -42.84262, -42.83058, 
        -42.81199, -42.78806, -42.75895, -42.72497, -42.68542, -42.64019, 
        -42.58854, -42.53242, -42.47444, -42.41726, -42.36454, -42.31903, 
        -42.28525,
  -40.27369, -40.29456, -40.31345, -40.33315, -40.35298, -40.37419, 
        -40.3961, -40.41885, -40.44226, -40.46561, -40.48963, -40.51418, 
        -40.53897, -40.56415, -40.59007, -40.61655, -40.64359, -40.67057, 
        -40.70018, -40.73254, -40.76897, -40.81082, -40.8595, -40.9158, 
        -40.98035, -41.05347, -41.13517, -41.22495, -41.32251, -41.4277, 
        -41.53979, -41.65784, -41.77983, -41.9069, -42.03656, -42.16824, 
        -42.30066, -42.43224, -42.56146, -42.68641, -42.80527, -42.9159, 
        -43.01681, -43.10749, -43.18755, -43.257, -43.31529, -43.3629, 
        -43.3986, -43.42463, -43.44103, -43.44884, -43.44869, -43.44248, 
        -43.4307, -43.41389, -43.39289, -43.36714, -43.33765, -43.30452, 
        -43.26837, -43.23041, -43.19147, -43.15204, -43.11138, -43.07206, 
        -43.03216, -42.99132, -42.94782, -42.9008, -42.85008, -42.79534, 
        -42.73792, -42.67945, -42.6232, -42.5715, -42.52736, -42.4924, 
        -42.46594, -42.44724, -42.43489, -42.42638, -42.41836, -42.41046, 
        -42.39893, -42.38203, -42.35891, -42.3308, -42.30119, -42.2714, 
        -42.24292, -42.21636, -42.18913, -42.15886, -42.12217, -42.0761, 
        -42.0201, -41.95306, -41.87506, -41.7879, -41.69369, -41.59774, 
        -41.50322, -41.41299, -41.32877, -41.25426, -41.19044, -41.13637, 
        -41.09183, -41.05565, -41.02578, -41.00254, -40.98452, -40.97163, 
        -40.96463, -40.96318, -40.96662, -40.97432, -40.98462, -40.99592, 
        -41.00925, -41.02247, -41.03498, -41.04692, -41.05805, -41.06946, 
        -41.08224, -41.0972, -41.11401, -41.13333, -41.15382, -41.17389, 
        -41.19135, -41.20347, -41.20896, -41.20635, -41.19492, -41.17509, 
        -41.14877, -41.11577, -41.0775, -41.0378, -40.99722, -40.95606, 
        -40.91511, -40.87435, -40.83339, -40.79205, -40.7483, -40.70454, 
        -40.65964, -40.61396, -40.56781, -40.52182, -40.47636, -40.43275, 
        -40.39171, -40.35382, -40.31779, -40.28592, -40.25635, -40.22823, 
        -40.2007, -40.17242, -40.1445, -40.11749, -40.09328, -40.07446, 
        -40.06458, -40.06505, -40.07898, -40.10775, -40.15107, -40.20724, 
        -40.2744, -40.34841, -40.42523, -40.50104, -40.57319, -40.64053, 
        -40.70359, -40.76428, -40.82597, -40.89303, -40.96848, -41.05481, 
        -41.15273, -41.26075, -41.37463, -41.49061, -41.60231, -41.70348, 
        -41.79064, -41.86103, -41.9152, -41.95527, -41.98679, -42.01686, 
        -42.05423, -42.10815, -42.18365, -42.28375, -42.40725, -42.54826, 
        -42.70063, -42.85705, -43.01103, -43.15845, -43.29498, -43.42029, 
        -43.53445, -43.63771, -43.7315, -43.81443, -43.88569, -43.9465, 
        -43.99654, -44.03815, -44.07137, -44.0989, -44.12318, -44.14746, 
        -44.17476, -44.20606, -44.24278, -44.28449, -44.32964, -44.37589, 
        -44.41953, -44.45937, -44.49379, -44.52229, -44.54426, -44.55867, 
        -44.5663, -44.5671, -44.56299, -44.55416, -44.53901, -44.51884, 
        -44.4921, -44.459, -44.41751, -44.36788, -44.30775, -44.23897, 
        -44.15905, -44.0713, -43.97535, -43.87108, -43.76332, -43.65173, 
        -43.53978, -43.43202, -43.3254, -43.22363, -43.12637, -43.03212, 
        -42.9382, -42.84265, -42.74592, -42.64551, -42.5447, -42.44073, 
        -42.34173, -42.24956, -42.16788, -42.10022, -42.05182, -42.024, 
        -42.01676, -42.0316, -42.06555, -42.11825, -42.18272, -42.25636, 
        -42.33411, -42.41021, -42.48254, -42.54763, -42.60355, -42.64891, 
        -42.68262, -42.70444, -42.71418, -42.71255, -42.70073, -42.68008, 
        -42.65292, -42.62094, -42.58508, -42.54479, -42.50222, -42.45605, 
        -42.40708, -42.35638, -42.30591, -42.25753, -42.21391, -42.17714, 
        -42.15029,
  -40.37732, -40.39821, -40.41762, -40.43693, -40.45698, -40.47812, 
        -40.50015, -40.52336, -40.54732, -40.57237, -40.59842, -40.62564, 
        -40.65298, -40.68221, -40.71246, -40.74362, -40.77586, -40.80865, 
        -40.84272, -40.87883, -40.91854, -40.96288, -41.01294, -41.06965, 
        -41.13385, -41.20557, -41.28492, -41.37091, -41.46489, -41.56542, 
        -41.67181, -41.78343, -41.89917, -42.01815, -42.13935, -42.26208, 
        -42.38547, -42.50792, -42.62834, -42.74476, -42.85546, -42.95855, 
        -43.05146, -43.13585, -43.21059, -43.27548, -43.33033, -43.37512, 
        -43.41001, -43.43484, -43.45082, -43.4592, -43.46045, -43.45621, 
        -43.44751, -43.43513, -43.41913, -43.39993, -43.37759, -43.35072, 
        -43.32143, -43.28948, -43.25563, -43.22061, -43.18465, -43.14817, 
        -43.11094, -43.07196, -43.03036, -42.98528, -42.93597, -42.88277, 
        -42.82647, -42.76924, -42.71338, -42.66187, -42.61631, -42.5803, 
        -42.55243, -42.53193, -42.51817, -42.50888, -42.50192, -42.49536, 
        -42.48633, -42.47273, -42.45312, -42.4287, -42.40187, -42.37471, 
        -42.34877, -42.32442, -42.30064, -42.2749, -42.24324, -42.20551, 
        -42.1589, -42.10208, -42.03468, -41.95789, -41.8743, -41.78675, 
        -41.69866, -41.61306, -41.53204, -41.45907, -41.39526, -41.34073, 
        -41.29546, -41.25849, -41.2282, -41.2037, -41.18495, -41.17034, 
        -41.1626, -41.16039, -41.1633, -41.17029, -41.18063, -41.19299, 
        -41.20655, -41.2198, -41.23176, -41.24278, -41.25248, -41.26193, 
        -41.272, -41.28354, -41.29714, -41.3134, -41.33159, -41.35011, 
        -41.3672, -41.37943, -41.38692, -41.38698, -41.37849, -41.3614, 
        -41.33704, -41.3055, -41.26894, -41.22922, -41.18782, -41.14604, 
        -41.10426, -41.06305, -41.02186, -40.98045, -40.9378, -40.89476, 
        -40.85075, -40.80591, -40.76037, -40.71525, -40.67068, -40.62682, 
        -40.58629, -40.54854, -40.51319, -40.48095, -40.45058, -40.42131, 
        -40.3921, -40.36285, -40.33315, -40.30421, -40.27782, -40.25656, 
        -40.2436, -40.24091, -40.25139, -40.27605, -40.31501, -40.36622, 
        -40.42759, -40.495, -40.56447, -40.6321, -40.69475, -40.75045, 
        -40.80149, -40.84915, -40.89717, -40.95004, -41.01175, -41.08515, 
        -41.17145, -41.26983, -41.37674, -41.48685, -41.59414, -41.69228, 
        -41.77668, -41.8445, -41.89578, -41.9334, -41.96334, -41.99385, 
        -42.03463, -42.09436, -42.17899, -42.28987, -42.42354, -42.57465, 
        -42.73499, -42.8969, -43.05211, -43.19766, -43.33018, -43.44854, 
        -43.55354, -43.64605, -43.72697, -43.79615, -43.85443, -43.90227, 
        -43.94038, -43.96939, -43.99176, -44.00879, -44.02358, -44.0388, 
        -44.05722, -44.08113, -44.11102, -44.14662, -44.18544, -44.22491, 
        -44.26267, -44.29577, -44.32322, -44.34374, -44.35629, -44.36181, 
        -44.36005, -44.35219, -44.3383, -44.31881, -44.29564, -44.26733, 
        -44.23409, -44.19434, -44.14668, -44.08967, -44.02254, -43.94555, 
        -43.85811, -43.76288, -43.65869, -43.54994, -43.43742, -43.3227, 
        -43.20824, -43.10024, -42.99395, -42.89384, -42.79945, -42.70953, 
        -42.62093, -42.5318, -42.44281, -42.3519, -42.2595, -42.16805, 
        -42.08302, -42.00602, -41.94051, -41.8901, -41.85905, -41.84824, 
        -41.85919, -41.89117, -41.94246, -42.01033, -42.08839, -42.17175, 
        -42.25631, -42.33686, -42.40983, -42.47257, -42.52351, -42.56219, 
        -42.58845, -42.60281, -42.60472, -42.59516, -42.57552, -42.54699, 
        -42.51144, -42.47141, -42.42847, -42.38372, -42.33751, -42.29082, 
        -42.24432, -42.19901, -42.15595, -42.11657, -42.08199, -42.05376, 
        -42.03378,
  -40.47526, -40.4956, -40.51428, -40.5328, -40.5526, -40.57363, 
        -40.59564, -40.61803, -40.64249, -40.66894, -40.697, -40.72666, 
        -40.75788, -40.79103, -40.82574, -40.86101, -40.89812, -40.93566, 
        -40.97426, -41.01457, -41.05785, -41.10507, -41.15626, -41.21432, 
        -41.2788, -41.34989, -41.42788, -41.51241, -41.60328, -41.69979, 
        -41.80114, -41.90678, -42.0157, -42.12733, -42.24048, -42.3545, 
        -42.46929, -42.58188, -42.69324, -42.8009, -42.90342, -42.9986, 
        -43.08524, -43.16328, -43.23247, -43.29273, -43.34398, -43.38594, 
        -43.41879, -43.44269, -43.45837, -43.4672, -43.46985, -43.46653, 
        -43.46064, -43.45229, -43.44161, -43.42839, -43.41297, -43.39418, 
        -43.37126, -43.34479, -43.31547, -43.28418, -43.25102, -43.21701, 
        -43.18177, -43.14464, -43.10484, -43.06174, -43.01378, -42.96322, 
        -42.91026, -42.85623, -42.80372, -42.75498, -42.71181, -42.67648, 
        -42.64855, -42.62699, -42.61162, -42.6008, -42.59303, -42.58651, 
        -42.57897, -42.56803, -42.55234, -42.53107, -42.50795, -42.48357, 
        -42.45949, -42.43658, -42.4149, -42.39206, -42.36595, -42.33427, 
        -42.29522, -42.24703, -42.18872, -42.1215, -42.04715, -41.96789, 
        -41.88705, -41.80721, -41.7308, -41.66024, -41.59646, -41.54229, 
        -41.49673, -41.45909, -41.42787, -41.40249, -41.38229, -41.36784, 
        -41.35889, -41.35562, -41.35756, -41.36396, -41.37408, -41.38646, 
        -41.4, -41.41319, -41.42495, -41.43506, -41.44368, -41.45103, 
        -41.45729, -41.46562, -41.47606, -41.48902, -41.50445, -41.52114, 
        -41.53778, -41.55204, -41.56153, -41.56431, -41.55904, -41.54526, 
        -41.52351, -41.49445, -41.45984, -41.4217, -41.38151, -41.34087, 
        -41.30029, -41.26039, -41.22062, -41.18004, -41.13953, -41.09835, 
        -41.05586, -41.01205, -40.96734, -40.92261, -40.87837, -40.83531, 
        -40.79435, -40.75586, -40.71981, -40.68587, -40.65354, -40.62188, 
        -40.59027, -40.5583, -40.52617, -40.49481, -40.46596, -40.44212, 
        -40.42591, -40.41978, -40.42501, -40.4448, -40.47765, -40.52205, 
        -40.57542, -40.63387, -40.69358, -40.75065, -40.80206, -40.84646, 
        -40.8847, -40.91903, -40.95341, -40.99244, -41.04063, -41.10146, 
        -41.17649, -41.26548, -41.36465, -41.46951, -41.57367, -41.66991, 
        -41.75359, -41.82127, -41.87282, -41.91116, -41.94149, -41.97514, 
        -42.0215, -42.08858, -42.18188, -42.30168, -42.4427, -42.60025, 
        -42.7643, -42.92646, -43.08018, -43.22095, -43.34632, -43.45543, 
        -43.54864, -43.62792, -43.69424, -43.74931, -43.79362, -43.82842, 
        -43.85461, -43.87357, -43.88723, -43.89629, -43.90393, -43.91264, 
        -43.92484, -43.94275, -43.96654, -43.99611, -44.02731, -44.06005, 
        -44.09092, -44.11653, -44.13578, -44.14683, -44.14931, -44.14473, 
        -44.13234, -44.11372, -44.08986, -44.06192, -44.02994, -43.99384, 
        -43.95362, -43.90708, -43.85263, -43.78769, -43.71268, -43.6273, 
        -43.53259, -43.43003, -43.32002, -43.20734, -43.09267, -42.9769, 
        -42.86214, -42.75573, -42.65084, -42.55356, -42.46442, -42.3798, 
        -42.29817, -42.21756, -42.1384, -42.05601, -41.97766, -41.89867, 
        -41.83028, -41.77211, -41.7265, -41.69663, -41.68619, -41.69684, 
        -41.72897, -41.78139, -41.8505, -41.93306, -42.02282, -42.11507, 
        -42.20409, -42.28631, -42.3577, -42.41631, -42.46152, -42.49355, 
        -42.51297, -42.5204, -42.51567, -42.49988, -42.47327, -42.43705, 
        -42.39379, -42.34511, -42.29427, -42.2427, -42.19183, -42.14335, 
        -42.09812, -42.05719, -42.02095, -41.98938, -41.96317, -41.94248, 
        -41.92896,
  -40.56448, -40.58463, -40.60195, -40.6201, -40.63926, -40.65962, 
        -40.68141, -40.70488, -40.72982, -40.75732, -40.78678, -40.81841, 
        -40.85264, -40.88927, -40.92739, -40.9672, -41.00828, -41.04889, 
        -41.09175, -41.13616, -41.18317, -41.23363, -41.28865, -41.34878, 
        -41.41457, -41.48629, -41.56342, -41.64652, -41.7348, -41.82769, 
        -41.9244, -42.0245, -42.12605, -42.23092, -42.33675, -42.44314, 
        -42.54898, -42.65417, -42.75682, -42.8558, -42.94967, -43.0369, 
        -43.11632, -43.18808, -43.25175, -43.30751, -43.35509, -43.3943, 
        -43.42444, -43.44758, -43.46323, -43.47286, -43.47726, -43.47725, 
        -43.47403, -43.46908, -43.46287, -43.45541, -43.44529, -43.43205, 
        -43.41446, -43.39241, -43.36681, -43.33829, -43.30666, -43.27476, 
        -43.24147, -43.20607, -43.16821, -43.12728, -43.08362, -43.03721, 
        -42.98848, -42.93953, -42.89176, -42.84718, -42.80731, -42.77368, 
        -42.74623, -42.72451, -42.70786, -42.69498, -42.68616, -42.6792, 
        -42.67219, -42.66288, -42.65036, -42.63376, -42.61386, -42.59246, 
        -42.57092, -42.54979, -42.52964, -42.50882, -42.48606, -42.45887, 
        -42.4249, -42.38312, -42.33277, -42.27231, -42.20571, -42.1339, 
        -42.06001, -41.98613, -41.91416, -41.8468, -41.78591, -41.73255, 
        -41.68692, -41.64853, -41.61661, -41.59035, -41.56958, -41.55426, 
        -41.54462, -41.54082, -41.54221, -41.54863, -41.55883, -41.57082, 
        -41.58503, -41.59869, -41.61086, -41.62085, -41.6288, -41.63488, 
        -41.64006, -41.64568, -41.65298, -41.66291, -41.67585, -41.69083, 
        -41.70676, -41.72156, -41.73276, -41.73837, -41.73614, -41.7256, 
        -41.70703, -41.68106, -41.64832, -41.61289, -41.57537, -41.53735, 
        -41.49959, -41.46272, -41.42613, -41.38952, -41.35196, -41.31333, 
        -41.27285, -41.23028, -41.18607, -41.14111, -41.09604, -41.05219, 
        -41.00959, -40.9692, -40.93102, -40.89461, -40.85945, -40.82457, 
        -40.78893, -40.75362, -40.71852, -40.68444, -40.65298, -40.62649, 
        -40.60719, -40.59753, -40.59942, -40.61357, -40.63962, -40.6761, 
        -40.72015, -40.76839, -40.81733, -40.86282, -40.90236, -40.9346, 
        -40.96048, -40.98246, -41.0044, -41.03098, -41.06713, -41.11654, 
        -41.18102, -41.25965, -41.35177, -41.45194, -41.5528, -41.64808, 
        -41.73217, -41.80134, -41.85497, -41.8962, -41.93156, -41.97022, 
        -42.02225, -42.09577, -42.19473, -42.31929, -42.46435, -42.62291, 
        -42.78492, -42.94308, -43.09052, -43.22306, -43.33819, -43.43536, 
        -43.51564, -43.58044, -43.63248, -43.67369, -43.70575, -43.72892, 
        -43.7465, -43.75768, -43.76529, -43.76999, -43.77349, -43.77792, 
        -43.78616, -43.79953, -43.81842, -43.8421, -43.8676, -43.89314, 
        -43.91544, -43.93229, -43.94171, -43.94193, -43.93351, -43.91714, 
        -43.89375, -43.86462, -43.83102, -43.79512, -43.75559, -43.7117, 
        -43.66333, -43.60939, -43.5471, -43.47369, -43.39016, -43.29713, 
        -43.19501, -43.08717, -42.97238, -42.85855, -42.74446, -42.63042, 
        -42.51858, -42.41563, -42.31229, -42.21834, -42.13791, -42.06475, 
        -41.99245, -41.92128, -41.85246, -41.78528, -41.72085, -41.65718, 
        -41.60766, -41.57108, -41.54717, -41.53997, -41.5538, -41.58764, 
        -41.64162, -41.7135, -41.79913, -41.89403, -41.99221, -42.08941, 
        -42.17944, -42.25924, -42.32691, -42.37984, -42.41878, -42.4444, 
        -42.45789, -42.45927, -42.4491, -42.42739, -42.39434, -42.35083, 
        -42.29903, -42.24108, -42.18013, -42.12046, -42.06345, -42.01162, 
        -41.96589, -41.92723, -41.89567, -41.87021, -41.85081, -41.83692, 
        -41.82872,
  -40.64402, -40.6646, -40.68306, -40.70102, -40.71917, -40.73892, 
        -40.76038, -40.7837, -40.80939, -40.83752, -40.86803, -40.90136, 
        -40.9369, -40.97617, -41.01775, -41.06113, -41.1055, -41.15087, 
        -41.19725, -41.24546, -41.29625, -41.35036, -41.40858, -41.4713, 
        -41.53909, -41.61173, -41.68901, -41.77002, -41.85609, -41.94568, 
        -42.03823, -42.13332, -42.23048, -42.32897, -42.42814, -42.52711, 
        -42.62526, -42.72203, -42.81639, -42.90694, -42.99252, -43.07194, 
        -43.14352, -43.20911, -43.26761, -43.31881, -43.3629, -43.39965, 
        -43.42937, -43.4521, -43.46819, -43.47869, -43.48475, -43.48689, 
        -43.48626, -43.48439, -43.48162, -43.47768, -43.47102, -43.46212, 
        -43.44851, -43.42985, -43.4068, -43.38063, -43.35216, -43.32183, 
        -43.29, -43.25623, -43.22041, -43.18242, -43.14227, -43.10046, 
        -43.05744, -43.01447, -42.97235, -42.93172, -42.8958, -42.86485, 
        -42.8391, -42.81797, -42.80112, -42.78838, -42.77856, -42.77098, 
        -42.76392, -42.75605, -42.74581, -42.73244, -42.71603, -42.69781, 
        -42.67847, -42.65937, -42.64065, -42.62054, -42.59956, -42.57499, 
        -42.54474, -42.5074, -42.46226, -42.40907, -42.34875, -42.28347, 
        -42.21516, -42.14649, -42.07882, -42.01441, -41.95537, -41.90278, 
        -41.85714, -41.81815, -41.78575, -41.75928, -41.73743, -41.7222, 
        -41.71273, -41.7092, -41.71128, -41.71848, -41.72986, -41.74432, 
        -41.76007, -41.77567, -41.78952, -41.80106, -41.80958, -41.81544, 
        -41.81973, -41.82373, -41.82886, -41.83636, -41.847, -41.86039, 
        -41.87471, -41.88987, -41.90241, -41.91008, -41.91068, -41.90331, 
        -41.8879, -41.86519, -41.83679, -41.80475, -41.77075, -41.73648, 
        -41.70256, -41.66953, -41.63683, -41.60407, -41.5699, -41.53376, 
        -41.49506, -41.45347, -41.40939, -41.36369, -41.31602, -41.27029, 
        -41.22507, -41.18185, -41.13993, -41.10012, -41.06105, -41.02214, 
        -40.98379, -40.9456, -40.90754, -40.87088, -40.83717, -40.80825, 
        -40.7865, -40.77392, -40.77172, -40.78051, -40.79969, -40.82784, 
        -40.86255, -40.9006, -40.93861, -40.97315, -41.00063, -41.02206, 
        -41.03743, -41.04914, -41.06086, -41.07751, -41.10359, -41.14329, 
        -41.19879, -41.27041, -41.35577, -41.45021, -41.54761, -41.64115, 
        -41.72503, -41.79532, -41.85145, -41.89581, -41.93579, -41.97934, 
        -42.03558, -42.11278, -42.21459, -42.33967, -42.48286, -42.63702, 
        -42.79311, -42.94211, -43.07988, -43.20138, -43.30431, -43.38804, 
        -43.45487, -43.50629, -43.54556, -43.57561, -43.59796, -43.61419, 
        -43.62544, -43.63271, -43.63723, -43.63949, -43.64133, -43.64437, 
        -43.65054, -43.66102, -43.67596, -43.69384, -43.71295, -43.73058, 
        -43.74394, -43.75058, -43.74884, -43.73761, -43.71748, -43.68976, 
        -43.65569, -43.61694, -43.57427, -43.53028, -43.48394, -43.4342, 
        -43.3792, -43.3173, -43.24619, -43.1634, -43.07124, -42.97023, 
        -42.86249, -42.75009, -42.63273, -42.52015, -42.40874, -42.29956, 
        -42.19334, -42.09348, -41.99768, -41.9166, -41.84847, -41.79083, 
        -41.73035, -41.66971, -41.61314, -41.55984, -41.51114, -41.46249, 
        -41.43274, -41.41624, -41.41489, -41.43219, -41.47017, -41.52618, 
        -41.60036, -41.68906, -41.78735, -41.89171, -41.99365, -42.09103, 
        -42.17921, -42.25441, -42.31553, -42.36197, -42.39466, -42.41463, 
        -42.42268, -42.41912, -42.40396, -42.37674, -42.33707, -42.28552, 
        -42.22405, -42.15622, -42.08593, -42.01691, -41.95226, -41.89517, 
        -41.84729, -41.80891, -41.77971, -41.75859, -41.74403, -41.73507, 
        -41.73114,
  -40.71443, -40.73623, -40.75542, -40.7735, -40.79156, -40.81088, 
        -40.8324, -40.85503, -40.88132, -40.91002, -40.94152, -40.97644, 
        -41.01469, -41.05641, -41.10043, -41.14643, -41.19385, -41.24231, 
        -41.29175, -41.3432, -41.39744, -41.45494, -41.51537, -41.58087, 
        -41.65062, -41.72462, -41.80248, -41.88373, -41.96785, -42.05429, 
        -42.14305, -42.23385, -42.32624, -42.41925, -42.51252, -42.60508, 
        -42.69608, -42.78423, -42.87041, -42.9528, -43.03049, -43.10264, 
        -43.16865, -43.22839, -43.28171, -43.3287, -43.36965, -43.40433, 
        -43.4329, -43.45549, -43.4724, -43.48411, -43.49159, -43.49468, 
        -43.49606, -43.49619, -43.49576, -43.49415, -43.4909, -43.48451, 
        -43.47344, -43.45695, -43.43557, -43.41113, -43.3844, -43.35583, 
        -43.3255, -43.29325, -43.25946, -43.22315, -43.18687, -43.14988, 
        -43.11264, -43.07593, -43.04003, -43.00606, -42.97496, -42.94753, 
        -42.92396, -42.90421, -42.88806, -42.87545, -42.86538, -42.85704, 
        -42.84999, -42.84276, -42.83436, -42.82281, -42.80984, -42.7947, 
        -42.77826, -42.76133, -42.74419, -42.72614, -42.70641, -42.68316, 
        -42.65474, -42.62008, -42.57835, -42.52932, -42.47389, -42.41336, 
        -42.34959, -42.28478, -42.22046, -42.15851, -42.09963, -42.04744, 
        -42.00157, -41.96252, -41.9303, -41.9048, -41.88535, -41.87142, 
        -41.86358, -41.86187, -41.86618, -41.87542, -41.88929, -41.90643, 
        -41.92529, -41.94372, -41.96059, -41.97436, -41.98473, -41.99083, 
        -41.99549, -41.99895, -42.00282, -42.00869, -42.01767, -42.0299, 
        -42.04433, -42.05953, -42.0728, -42.08195, -42.0846, -42.07947, 
        -42.06664, -42.04656, -42.0212, -41.99268, -41.96256, -41.93247, 
        -41.90294, -41.87442, -41.84631, -41.81658, -41.78605, -41.75252, 
        -41.71552, -41.67464, -41.63025, -41.5837, -41.53529, -41.48767, 
        -41.43985, -41.39377, -41.34937, -41.30581, -41.26298, -41.22059, 
        -41.17836, -41.13636, -41.09504, -41.05549, -41.0191, -40.98748, 
        -40.96316, -40.94772, -40.94067, -40.94451, -40.95745, -40.97804, 
        -41.00415, -41.03298, -41.06166, -41.08676, -41.10633, -41.1195, 
        -41.12707, -41.13173, -41.13625, -41.14567, -41.16397, -41.19536, 
        -41.24248, -41.306, -41.38401, -41.47189, -41.56417, -41.6543, 
        -41.73625, -41.8065, -41.86403, -41.91122, -41.9531, -42.00014, 
        -42.05872, -42.13745, -42.23787, -42.35901, -42.49575, -42.64085, 
        -42.78644, -42.92493, -43.05047, -43.15881, -43.24818, -43.31858, 
        -43.37254, -43.41129, -43.43954, -43.46157, -43.47764, -43.48986, 
        -43.49841, -43.50495, -43.50928, -43.51221, -43.51468, -43.51792, 
        -43.52341, -43.53157, -43.54305, -43.5546, -43.56731, -43.57678, 
        -43.58058, -43.57692, -43.56382, -43.54111, -43.50968, -43.47092, 
        -43.42691, -43.38031, -43.3323, -43.28264, -43.23124, -43.17609, 
        -43.11468, -43.04412, -42.96366, -42.87165, -42.77076, -42.66302, 
        -42.54962, -42.43067, -42.30433, -42.19835, -42.08674, -41.9774, 
        -41.87473, -41.79336, -41.72231, -41.65651, -41.60516, -41.55314, 
        -41.50182, -41.45267, -41.40966, -41.37203, -41.34264, -41.31527, 
        -41.30675, -41.312, -41.33405, -41.37379, -41.43505, -41.51144, 
        -41.60259, -41.70459, -41.81272, -41.92213, -42.02614, -42.11994, 
        -42.20179, -42.27012, -42.32366, -42.36336, -42.38988, -42.40488, 
        -42.40858, -42.40063, -42.38071, -42.34772, -42.30107, -42.24102, 
        -42.16959, -42.09057, -42.00873, -41.92868, -41.85514, -41.79133, 
        -41.73911, -41.69893, -41.66979, -41.64994, -41.6375, -41.6313, 
        -41.62978,
  -40.77695, -40.8004, -40.8201, -40.83869, -40.85697, -40.87652, 
        -40.89794, -40.92249, -40.94907, -40.97821, -41.01072, -41.04662, 
        -41.08634, -41.12951, -41.17543, -41.22357, -41.27237, -41.32315, 
        -41.37558, -41.42993, -41.48679, -41.54715, -41.61092, -41.6787, 
        -41.75033, -41.82547, -41.90361, -41.9844, -42.06725, -42.1514, 
        -42.23742, -42.32445, -42.41167, -42.50006, -42.58808, -42.67467, 
        -42.75917, -42.84118, -42.91995, -42.99496, -43.06538, -43.13078, 
        -43.19046, -43.24437, -43.29282, -43.33591, -43.37381, -43.40581, 
        -43.43352, -43.45614, -43.47394, -43.48685, -43.49564, -43.50164, 
        -43.50483, -43.50639, -43.50686, -43.50621, -43.50381, -43.49814, 
        -43.48796, -43.47303, -43.45327, -43.42999, -43.40361, -43.3763, 
        -43.34729, -43.31661, -43.28495, -43.25217, -43.21941, -43.18707, 
        -43.15525, -43.12437, -43.09448, -43.06627, -43.04008, -43.01638, 
        -42.99553, -42.9777, -42.96292, -42.95016, -42.94019, -42.93229, 
        -42.92554, -42.91913, -42.9123, -42.9043, -42.89442, -42.88287, 
        -42.86935, -42.85484, -42.83915, -42.82215, -42.80299, -42.7802, 
        -42.75266, -42.71943, -42.67974, -42.63255, -42.58028, -42.52287, 
        -42.46237, -42.40011, -42.33787, -42.27707, -42.21982, -42.16779, 
        -42.12215, -42.08354, -42.05235, -42.02831, -42.01114, -42.00057, 
        -41.99612, -41.99787, -42.00554, -42.01876, -42.03566, -42.05699, 
        -42.0798, -42.1024, -42.12328, -42.141, -42.15456, -42.16401, 
        -42.17007, -42.17434, -42.17846, -42.1838, -42.19191, -42.20312, 
        -42.2167, -42.23163, -42.24506, -42.25474, -42.25831, -42.25435, 
        -42.24316, -42.22421, -42.2015, -42.17599, -42.14964, -42.12351, 
        -42.09847, -42.07438, -42.0504, -42.02557, -41.99831, -41.96729, 
        -41.93202, -41.89158, -41.8468, -41.79899, -41.74979, -41.69968, 
        -41.65031, -41.60224, -41.55523, -41.50887, -41.46309, -41.41742, 
        -41.37061, -41.32507, -41.28044, -41.23775, -41.19893, -41.16488, 
        -41.1381, -41.11981, -41.11053, -41.11016, -41.11784, -41.13187, 
        -41.15078, -41.17204, -41.19316, -41.21123, -41.22448, -41.23237, 
        -41.23542, -41.23581, -41.23618, -41.24091, -41.25369, -41.27848, 
        -41.31839, -41.37307, -41.44289, -41.52277, -41.60764, -41.69129, 
        -41.76847, -41.83548, -41.89158, -41.93903, -41.98273, -42.0308, 
        -42.08959, -42.16507, -42.26069, -42.37435, -42.50116, -42.6347, 
        -42.76748, -42.89249, -43.00415, -43.09895, -43.17524, -43.23313, 
        -43.27514, -43.3047, -43.3264, -43.34232, -43.35579, -43.36569, 
        -43.3746, -43.38164, -43.38725, -43.39156, -43.39493, -43.39945, 
        -43.40461, -43.41119, -43.42036, -43.42885, -43.43504, -43.4361, 
        -43.43135, -43.4178, -43.3942, -43.36096, -43.31937, -43.27176, 
        -43.22104, -43.16914, -43.1165, -43.06369, -43.00874, -42.94872, 
        -42.88049, -42.80212, -42.71239, -42.61062, -42.501, -42.38696, 
        -42.26771, -42.13395, -41.99623, -41.88397, -41.78552, -41.70469, 
        -41.62591, -41.5801, -41.5269, -41.46761, -41.41673, -41.37281, 
        -41.33091, -41.29291, -41.26316, -41.24018, -41.22703, -41.22143, 
        -41.23576, -41.26046, -41.30746, -41.36843, -41.44817, -41.53968, 
        -41.64256, -41.75404, -41.86677, -41.97637, -42.0771, -42.1655, 
        -42.24017, -42.30042, -42.34671, -42.38008, -42.4019, -42.41283, 
        -42.4124, -42.40015, -42.37497, -42.33561, -42.28093, -42.21135, 
        -42.12914, -42.03746, -41.9438, -41.85265, -41.76941, -41.69777, 
        -41.63986, -41.59589, -41.56435, -41.54374, -41.53152, -41.52604, 
        -41.52554,
  -40.83246, -40.85799, -40.88025, -40.90014, -40.91917, -40.93913, 
        -40.9611, -40.98568, -41.01287, -41.04314, -41.07624, -41.11192, 
        -41.15256, -41.19689, -41.24393, -41.29351, -41.34507, -41.39803, 
        -41.45278, -41.50919, -41.5682, -41.63023, -41.6958, -41.76485, 
        -41.83739, -41.9132, -41.99055, -42.07088, -42.15271, -42.23523, 
        -42.31924, -42.40355, -42.48804, -42.57258, -42.65562, -42.73728, 
        -42.81618, -42.89175, -42.96386, -43.03199, -43.09591, -43.1548, 
        -43.20753, -43.25595, -43.29976, -43.33925, -43.37439, -43.40572, 
        -43.43274, -43.45562, -43.47407, -43.48814, -43.49875, -43.50612, 
        -43.51017, -43.51221, -43.51298, -43.51233, -43.50832, -43.50251, 
        -43.49258, -43.47798, -43.45921, -43.43709, -43.41258, -43.38626, 
        -43.35879, -43.32946, -43.29972, -43.26969, -43.24001, -43.21144, 
        -43.18423, -43.15841, -43.13379, -43.10953, -43.0878, -43.06779, 
        -43.04996, -43.03456, -43.02159, -43.01107, -43.0023, -42.99508, 
        -42.98923, -42.98422, -42.97923, -42.97363, -42.96661, -42.95836, 
        -42.9482, -42.9361, -42.92237, -42.90538, -42.88648, -42.86388, 
        -42.83635, -42.80365, -42.76496, -42.72055, -42.67025, -42.6148, 
        -42.55564, -42.49498, -42.43328, -42.37318, -42.31589, -42.26396, 
        -42.21893, -42.1816, -42.15253, -42.13148, -42.11724, -42.11123, 
        -42.1118, -42.11866, -42.1314, -42.14977, -42.17275, -42.19917, 
        -42.22697, -42.25455, -42.28033, -42.30266, -42.3203, -42.33302, 
        -42.34174, -42.34776, -42.35295, -42.35894, -42.3667, -42.37706, 
        -42.38904, -42.40318, -42.41631, -42.42548, -42.42886, -42.42532, 
        -42.41492, -42.39828, -42.37737, -42.35447, -42.33123, -42.30883, 
        -42.28769, -42.26761, -42.24741, -42.22607, -42.20167, -42.17258, 
        -42.13876, -42.099, -42.05416, -42.00611, -41.9555, -41.90499, 
        -41.85445, -41.80508, -41.75679, -41.70916, -41.66113, -41.61278, 
        -41.56413, -41.51559, -41.46813, -41.42295, -41.38141, -41.34563, 
        -41.31672, -41.29604, -41.2837, -41.27954, -41.28232, -41.29139, 
        -41.30432, -41.32009, -41.33571, -41.34914, -41.35773, -41.36298, 
        -41.36427, -41.36323, -41.36206, -41.36409, -41.3731, -41.39243, 
        -41.42558, -41.47331, -41.53405, -41.60413, -41.67874, -41.75279, 
        -41.82158, -41.88202, -41.93385, -41.97836, -42.02042, -42.06636, 
        -42.12204, -42.19304, -42.281, -42.38464, -42.49957, -42.61933, 
        -42.73795, -42.84762, -42.94558, -43.02725, -43.09147, -43.13881, 
        -43.17216, -43.19507, -43.2122, -43.22629, -43.239, -43.2505, 
        -43.26083, -43.26886, -43.27592, -43.28209, -43.28658, -43.29127, 
        -43.2961, -43.30216, -43.30878, -43.31345, -43.31402, -43.30906, 
        -43.29573, -43.27336, -43.241, -43.19932, -43.1505, -43.09692, 
        -43.04159, -42.98547, -42.93149, -42.87669, -42.81912, -42.75462, 
        -42.68036, -42.5943, -42.49572, -42.38583, -42.26926, -42.14922, 
        -42.02161, -41.8862, -41.74707, -41.64448, -41.57055, -41.51897, 
        -41.47375, -41.44078, -41.39656, -41.35055, -41.29788, -41.25305, 
        -41.21386, -41.19007, -41.18713, -41.18351, -41.18973, -41.20023, 
        -41.23005, -41.27508, -41.33331, -41.40876, -41.49779, -41.59914, 
        -41.71017, -41.8249, -41.93785, -42.04376, -42.13879, -42.22007, 
        -42.28736, -42.34074, -42.38038, -42.4086, -42.42653, -42.43403, 
        -42.42984, -42.41324, -42.38247, -42.33587, -42.27255, -42.19285, 
        -42.09954, -41.99693, -41.89131, -41.78927, -41.69604, -41.61596, 
        -41.55122, -41.50179, -41.46626, -41.44305, -41.42875, -41.42233, 
        -41.42127,
  -40.88445, -40.91251, -40.93668, -40.95799, -40.97833, -40.99892, 
        -41.02152, -41.04568, -41.0735, -41.10435, -41.13855, -41.17609, 
        -41.21725, -41.26191, -41.30984, -41.36031, -41.41306, -41.46764, 
        -41.52392, -41.58172, -41.6417, -41.70364, -41.76959, -41.83899, 
        -41.91193, -41.98746, -42.06543, -42.14541, -42.22665, -42.30821, 
        -42.39031, -42.47253, -42.55426, -42.63512, -42.71465, -42.7915, 
        -42.86538, -42.93436, -43.00049, -43.06252, -43.12016, -43.17328, 
        -43.22161, -43.26512, -43.3048, -43.34081, -43.37353, -43.40314, 
        -43.4294, -43.45219, -43.47141, -43.4866, -43.49712, -43.50547, 
        -43.51074, -43.51297, -43.51356, -43.5116, -43.5073, -43.50035, 
        -43.48974, -43.47528, -43.45719, -43.43549, -43.41184, -43.38662, 
        -43.36037, -43.333, -43.30493, -43.27602, -43.24916, -43.22332, 
        -43.19967, -43.17758, -43.15714, -43.13792, -43.12009, -43.10351, 
        -43.08869, -43.07548, -43.06451, -43.05567, -43.04843, -43.04282, 
        -43.03848, -43.03502, -43.032, -43.02779, -43.02375, -43.0186, 
        -43.0117, -43.00232, -42.99064, -42.976, -42.95769, -42.93519, 
        -42.90775, -42.87513, -42.8369, -42.79309, -42.74371, -42.68947, 
        -42.63093, -42.56996, -42.50842, -42.44712, -42.39015, -42.33863, 
        -42.29458, -42.25942, -42.23359, -42.21689, -42.20922, -42.20913, 
        -42.21648, -42.22995, -42.24909, -42.27368, -42.30256, -42.33442, 
        -42.3677, -42.4006, -42.43153, -42.45872, -42.48072, -42.4963, 
        -42.50821, -42.51648, -42.52348, -42.5311, -42.53922, -42.5493, 
        -42.56159, -42.57483, -42.58653, -42.59472, -42.59726, -42.59325, 
        -42.58262, -42.56664, -42.54715, -42.52607, -42.5054, -42.48596, 
        -42.46817, -42.45145, -42.43353, -42.41489, -42.3929, -42.36581, 
        -42.33315, -42.29422, -42.25061, -42.20336, -42.15419, -42.10429, 
        -42.05416, -42.00509, -41.95696, -41.90929, -41.8606, -41.81091, 
        -41.7603, -41.70984, -41.6602, -41.61276, -41.5694, -41.53144, 
        -41.50041, -41.47639, -41.46191, -41.45446, -41.45337, -41.45779, 
        -41.46644, -41.47784, -41.49007, -41.50095, -41.50912, -41.514, 
        -41.51564, -41.51485, -41.51323, -41.51406, -41.51998, -41.53479, 
        -41.56124, -41.60005, -41.65029, -41.7085, -41.77055, -41.83209, 
        -41.8893, -41.94039, -41.98454, -42.02224, -42.06043, -42.10232, 
        -42.15321, -42.21766, -42.29665, -42.38866, -42.49094, -42.5969, 
        -42.70084, -42.79704, -42.88165, -42.9513, -43.00505, -43.04412, 
        -43.07117, -43.09039, -43.10556, -43.11951, -43.13389, -43.14629, 
        -43.15773, -43.16751, -43.17552, -43.18193, -43.18711, -43.19174, 
        -43.19638, -43.20143, -43.20486, -43.20626, -43.20266, -43.19221, 
        -43.17263, -43.14317, -43.10394, -43.05632, -43.00288, -42.94627, 
        -42.88935, -42.83402, -42.78058, -42.72558, -42.66618, -42.5968, 
        -42.51701, -42.42348, -42.31705, -42.20053, -42.07935, -41.95584, 
        -41.82701, -41.69889, -41.57624, -41.49127, -41.43783, -41.39754, 
        -41.36552, -41.33927, -41.30795, -41.27332, -41.23279, -41.19561, 
        -41.17426, -41.16477, -41.17372, -41.18786, -41.20769, -41.2299, 
        -41.27328, -41.32808, -41.39559, -41.4769, -41.57388, -41.68024, 
        -41.79316, -41.90732, -42.01705, -42.11848, -42.20674, -42.28092, 
        -42.34141, -42.38863, -42.42382, -42.44825, -42.46272, -42.46706, 
        -42.45968, -42.43859, -42.40167, -42.34715, -42.2748, -42.18501, 
        -42.08052, -41.96695, -41.85002, -41.7371, -41.63409, -41.54532, 
        -41.47311, -41.41709, -41.37632, -41.34832, -41.33071, -41.32148, 
        -41.31889,
  -40.93389, -40.96435, -40.98959, -41.01271, -41.03398, -41.05594, 
        -41.07939, -41.10522, -41.13395, -41.1656, -41.2004, -41.23861, 
        -41.28027, -41.3251, -41.37338, -41.42444, -41.47705, -41.53247, 
        -41.58942, -41.64786, -41.70807, -41.77053, -41.83601, -41.90486, 
        -41.97682, -42.05165, -42.12872, -42.2081, -42.2883, -42.36958, 
        -42.45038, -42.52983, -42.60946, -42.68763, -42.7635, -42.83634, 
        -42.90559, -42.97051, -43.03111, -43.08758, -43.13976, -43.18782, 
        -43.23128, -43.27061, -43.3066, -43.33935, -43.36967, -43.39651, 
        -43.42189, -43.44465, -43.46402, -43.47993, -43.49204, -43.50101, 
        -43.50682, -43.50913, -43.50869, -43.50557, -43.49978, -43.49118, 
        -43.47982, -43.46489, -43.44668, -43.42476, -43.40179, -43.37769, 
        -43.3528, -43.32729, -43.30143, -43.27578, -43.25029, -43.22656, 
        -43.20523, -43.18539, -43.16778, -43.15156, -43.13675, -43.12318, 
        -43.11068, -43.09959, -43.0905, -43.08251, -43.07718, -43.07349, 
        -43.07112, -43.06974, -43.06891, -43.06789, -43.06672, -43.06462, 
        -43.0609, -43.05455, -43.04516, -43.03207, -43.01476, -42.9927, 
        -42.96533, -42.93309, -42.89523, -42.85081, -42.8018, -42.74752, 
        -42.68906, -42.62786, -42.56601, -42.50559, -42.44878, -42.39814, 
        -42.35619, -42.32399, -42.30238, -42.29144, -42.29048, -42.29802, 
        -42.31304, -42.33424, -42.36134, -42.39278, -42.42679, -42.46436, 
        -42.50275, -42.5406, -42.57606, -42.60764, -42.63391, -42.65412, 
        -42.6691, -42.68034, -42.68935, -42.69833, -42.70744, -42.71768, 
        -42.72951, -42.74142, -42.75187, -42.75835, -42.75959, -42.75474, 
        -42.74364, -42.72681, -42.70831, -42.6889, -42.6702, -42.65326, 
        -42.63834, -42.62436, -42.61015, -42.5939, -42.57383, -42.54853, 
        -42.51731, -42.47996, -42.43806, -42.39222, -42.34494, -42.29763, 
        -42.24981, -42.20198, -42.15577, -42.10846, -42.06035, -42.00984, 
        -41.95957, -41.90781, -41.85681, -41.80819, -41.76355, -41.72393, 
        -41.69146, -41.66646, -41.64912, -41.63865, -41.63415, -41.63478, 
        -41.63973, -41.64781, -41.65762, -41.66718, -41.67513, -41.68068, 
        -41.68324, -41.68369, -41.68267, -41.68272, -41.68587, -41.69637, 
        -41.7145, -41.74378, -41.78211, -41.8269, -41.87445, -41.92128, 
        -41.96464, -42.00344, -42.0381, -42.06965, -42.10163, -42.13816, 
        -42.1827, -42.24008, -42.30991, -42.39091, -42.48047, -42.57276, 
        -42.66276, -42.74604, -42.81822, -42.87713, -42.92221, -42.95494, 
        -42.9779, -42.99526, -43.01044, -43.02477, -43.0392, -43.05384, 
        -43.06557, -43.07587, -43.08352, -43.08919, -43.09363, -43.09785, 
        -43.10197, -43.10587, -43.10847, -43.10727, -43.10056, -43.08593, 
        -43.06198, -43.0276, -42.98406, -42.93309, -42.87797, -42.82151, 
        -42.76585, -42.71198, -42.65949, -42.60467, -42.54401, -42.47157, 
        -42.3862, -42.28662, -42.17361, -42.05245, -41.92795, -41.8041, 
        -41.67907, -41.56043, -41.4637, -41.39762, -41.34942, -41.31315, 
        -41.28472, -41.26498, -41.24348, -41.22279, -41.2016, -41.18345, 
        -41.17899, -41.18609, -41.20269, -41.22745, -41.25777, -41.29204, 
        -41.34333, -41.40644, -41.47955, -41.56631, -41.66548, -41.77256, 
        -41.8835, -41.99417, -42.09844, -42.19319, -42.27462, -42.34284, 
        -42.39803, -42.44098, -42.47289, -42.49477, -42.50673, -42.50815, 
        -42.49718, -42.47147, -42.42846, -42.36653, -42.285, -42.18573, 
        -42.07013, -41.94569, -41.81863, -41.69583, -41.5836, -41.48652, 
        -41.40611, -41.3428, -41.29597, -41.26211, -41.23932, -41.22594, 
        -41.2198,
  -40.9803, -41.01336, -41.04129, -41.06617, -41.08916, -41.11278, 
        -41.13707, -41.164, -41.19362, -41.22598, -41.26148, -41.29908, 
        -41.34105, -41.38644, -41.43499, -41.48627, -41.54005, -41.59562, 
        -41.65263, -41.7109, -41.77028, -41.8316, -41.89554, -41.96267, 
        -42.03305, -42.1064, -42.1814, -42.25928, -42.33902, -42.41932, 
        -42.49917, -42.5781, -42.65577, -42.73145, -42.80409, -42.87312, 
        -42.93817, -42.99857, -43.05414, -43.10568, -43.15295, -43.19634, 
        -43.23505, -43.27064, -43.30329, -43.33337, -43.36124, -43.38725, 
        -43.41157, -43.4337, -43.45314, -43.46907, -43.48171, -43.49082, 
        -43.49647, -43.49889, -43.49771, -43.49325, -43.48531, -43.47556, 
        -43.46262, -43.44688, -43.42867, -43.40829, -43.38598, -43.3632, 
        -43.34003, -43.31654, -43.29275, -43.26888, -43.24451, -43.22184, 
        -43.20129, -43.18283, -43.16678, -43.15157, -43.13861, -43.12711, 
        -43.11648, -43.10723, -43.09978, -43.09466, -43.0914, -43.08981, 
        -43.08971, -43.0906, -43.09193, -43.09348, -43.09504, -43.09562, 
        -43.09475, -43.09137, -43.08341, -43.07195, -43.05638, -43.03524, 
        -43.00886, -42.97731, -42.94012, -42.89722, -42.84855, -42.79458, 
        -42.7361, -42.67469, -42.61259, -42.55234, -42.49633, -42.4474, 
        -42.40772, -42.37951, -42.36317, -42.35768, -42.3643, -42.38046, 
        -42.40436, -42.43439, -42.46909, -42.5078, -42.54917, -42.5919, 
        -42.63472, -42.67658, -42.71568, -42.75049, -42.77991, -42.80323, 
        -42.82101, -42.8345, -42.84557, -42.85575, -42.86601, -42.87651, 
        -42.88658, -42.89743, -42.9061, -42.91118, -42.91119, -42.90522, 
        -42.8938, -42.87825, -42.86051, -42.84247, -42.82558, -42.81095, 
        -42.79845, -42.78703, -42.77511, -42.76096, -42.74281, -42.7194, 
        -42.69015, -42.65489, -42.61528, -42.57132, -42.52714, -42.48239, 
        -42.43779, -42.39375, -42.34974, -42.30528, -42.2592, -42.21132, 
        -42.16109, -42.11021, -42.05972, -42.01131, -41.96557, -41.92526, 
        -41.89121, -41.86442, -41.84471, -41.8313, -41.82312, -41.82014, 
        -41.82178, -41.82689, -41.83457, -41.8419, -41.84984, -41.85617, 
        -41.86012, -41.86149, -41.86079, -41.85998, -41.86115, -41.8661, 
        -41.87807, -41.89663, -41.92268, -41.95276, -41.98482, -42.01609, 
        -42.04487, -42.07056, -42.09417, -42.11749, -42.14231, -42.17239, 
        -42.21097, -42.2605, -42.32178, -42.3932, -42.47104, -42.55127, 
        -42.62782, -42.69874, -42.75969, -42.80916, -42.84708, -42.87506, 
        -42.8954, -42.91185, -42.92716, -42.94218, -42.95717, -42.97149, 
        -42.98367, -42.99306, -42.99962, -43.00402, -43.00739, -43.01023, 
        -43.01307, -43.01581, -43.0173, -43.01399, -43.00504, -42.98801, 
        -42.96119, -42.92414, -42.87876, -42.82743, -42.77299, -42.71924, 
        -42.667, -42.61559, -42.56527, -42.51081, -42.44884, -42.37351, 
        -42.28359, -42.17904, -42.06165, -41.93738, -41.81173, -41.68982, 
        -41.57397, -41.47086, -41.38924, -41.33293, -41.29272, -41.26721, 
        -41.24737, -41.24184, -41.23559, -41.22967, -41.22345, -41.22509, 
        -41.23286, -41.24812, -41.27042, -41.30031, -41.3378, -41.37959, 
        -41.43478, -41.50066, -41.5773, -41.66447, -41.76189, -41.86606, 
        -41.97327, -42.07829, -42.17588, -42.26381, -42.33996, -42.40333, 
        -42.45456, -42.49465, -42.52453, -42.5449, -42.55483, -42.5537, 
        -42.53918, -42.50862, -42.45987, -42.3911, -42.30202, -42.19399, 
        -42.07035, -41.93699, -41.80072, -41.669, -41.54799, -41.44217, 
        -41.35348, -41.28227, -41.22745, -41.18693, -41.15879, -41.14, 
        -41.12805,
  -41.02632, -41.06033, -41.09049, -41.11727, -41.14252, -41.1675, 
        -41.19252, -41.22044, -41.25104, -41.28412, -41.32008, -41.35928, 
        -41.40189, -41.4477, -41.49655, -41.54792, -41.60146, -41.65683, 
        -41.71329, -41.77051, -41.82866, -41.88727, -41.94915, -42.01404, 
        -42.08208, -42.15314, -42.22717, -42.30366, -42.3819, -42.46102, 
        -42.5397, -42.61703, -42.6925, -42.76582, -42.83509, -42.90057, 
        -42.96048, -43.01666, -43.06801, -43.11517, -43.15833, -43.19793, 
        -43.23403, -43.2666, -43.29615, -43.32378, -43.34958, -43.37379, 
        -43.39651, -43.41776, -43.43653, -43.4527, -43.46403, -43.47327, 
        -43.47911, -43.48116, -43.4794, -43.47391, -43.46561, -43.45451, 
        -43.4409, -43.4247, -43.40622, -43.38634, -43.36497, -43.34365, 
        -43.32214, -43.30061, -43.27872, -43.25507, -43.23209, -43.20991, 
        -43.18913, -43.17096, -43.15518, -43.14164, -43.12982, -43.11928, 
        -43.11005, -43.10254, -43.09671, -43.09322, -43.092, -43.09245, 
        -43.09449, -43.09747, -43.10004, -43.10426, -43.10834, -43.11169, 
        -43.1135, -43.11246, -43.10765, -43.09875, -43.08492, -43.06554, 
        -43.04105, -43.01112, -42.97521, -42.93343, -42.8856, -42.83237, 
        -42.77431, -42.7135, -42.65219, -42.59176, -42.53731, -42.49066, 
        -42.45406, -42.43029, -42.41975, -42.4223, -42.43724, -42.46253, 
        -42.49569, -42.53452, -42.57719, -42.62263, -42.66963, -42.71682, 
        -42.76312, -42.8073, -42.84838, -42.88517, -42.91666, -42.94091, 
        -42.96061, -42.97598, -42.98866, -43.00006, -43.01096, -43.02168, 
        -43.03215, -43.0416, -43.04909, -43.05306, -43.05216, -43.04564, 
        -43.0342, -43.0192, -43.00263, -42.98611, -42.9712, -42.95868, 
        -42.94831, -42.93904, -42.92809, -42.91604, -42.90011, -42.87852, 
        -42.85101, -42.81816, -42.78103, -42.74151, -42.70091, -42.66027, 
        -42.61932, -42.57968, -42.53978, -42.49825, -42.45512, -42.4095, 
        -42.36184, -42.3129, -42.26391, -42.21646, -42.17145, -42.13092, 
        -42.09631, -42.06726, -42.04515, -42.0285, -42.0172, -42.01024, 
        -42.00825, -42.01056, -42.01556, -42.0227, -42.03011, -42.03671, 
        -42.04116, -42.04328, -42.04299, -42.04082, -42.03873, -42.03879, 
        -42.04279, -42.05128, -42.0638, -42.07971, -42.09596, -42.11155, 
        -42.1258, -42.1389, -42.15164, -42.16479, -42.18231, -42.20592, 
        -42.23861, -42.28167, -42.33512, -42.39774, -42.46583, -42.53528, 
        -42.60196, -42.66199, -42.71324, -42.75436, -42.78606, -42.80985, 
        -42.82829, -42.84371, -42.85825, -42.87276, -42.8867, -42.89919, 
        -42.90984, -42.91726, -42.92197, -42.92461, -42.92633, -42.92754, 
        -42.93039, -42.93213, -42.93, -42.92531, -42.91523, -42.89681, 
        -42.8686, -42.83118, -42.78633, -42.73676, -42.6858, -42.63642, 
        -42.58847, -42.54211, -42.49425, -42.4406, -42.37716, -42.29939, 
        -42.20658, -42.09892, -41.97954, -41.8544, -41.72969, -41.61096, 
        -41.50385, -41.41339, -41.34032, -41.29339, -41.2627, -41.24701, 
        -41.2423, -41.24723, -41.25259, -41.25924, -41.26799, -41.28043, 
        -41.30119, -41.32328, -41.35295, -41.38903, -41.43144, -41.4775, 
        -41.5349, -41.60054, -41.67606, -41.76051, -41.8536, -41.95326, 
        -42.05602, -42.1555, -42.24789, -42.33122, -42.40303, -42.46323, 
        -42.51207, -42.5504, -42.57902, -42.59799, -42.60649, -42.60304, 
        -42.58496, -42.55038, -42.49662, -42.42207, -42.32687, -42.21207, 
        -42.08154, -41.94081, -41.79702, -41.65731, -41.52792, -41.41362, 
        -41.31618, -41.23616, -41.17266, -41.12424, -41.08877, -41.06367, 
        -41.0463,
  -41.06997, -41.10486, -41.13494, -41.16385, -41.19138, -41.21838, 
        -41.24614, -41.27562, -41.30734, -41.3413, -41.37804, -41.41798, 
        -41.46117, -41.50748, -41.55681, -41.6081, -41.66021, -41.71487, 
        -41.77027, -41.82618, -41.88292, -41.94046, -41.99979, -42.06218, 
        -42.12746, -42.19576, -42.26697, -42.34132, -42.41764, -42.49487, 
        -42.57196, -42.6465, -42.71952, -42.78989, -42.85572, -42.9173, 
        -42.97443, -43.02688, -43.07474, -43.11858, -43.15867, -43.1951, 
        -43.22824, -43.25808, -43.28536, -43.31041, -43.33384, -43.35485, 
        -43.37593, -43.39557, -43.41362, -43.42889, -43.44161, -43.45062, 
        -43.45632, -43.45812, -43.45616, -43.45007, -43.44074, -43.42857, 
        -43.41408, -43.39764, -43.37952, -43.35911, -43.33916, -43.31903, 
        -43.2995, -43.27974, -43.25946, -43.23822, -43.2158, -43.19356, 
        -43.17241, -43.15355, -43.13745, -43.12349, -43.11158, -43.10155, 
        -43.09332, -43.08699, -43.08176, -43.0799, -43.08046, -43.083, 
        -43.08674, -43.09167, -43.09729, -43.10379, -43.11034, -43.11634, 
        -43.12062, -43.12182, -43.11946, -43.11271, -43.10134, -43.08471, 
        -43.06268, -43.03509, -43.00034, -42.96049, -42.91427, -42.86255, 
        -42.80623, -42.74693, -42.68728, -42.62963, -42.57756, -42.53396, 
        -42.50183, -42.48275, -42.47825, -42.48809, -42.51144, -42.54546, 
        -42.58738, -42.63446, -42.68441, -42.7357, -42.7861, -42.83648, 
        -42.8846, -42.9299, -42.97149, -43.00861, -43.0406, -43.06678, 
        -43.08752, -43.10399, -43.11787, -43.13026, -43.14163, -43.15226, 
        -43.16201, -43.17036, -43.17679, -43.18012, -43.17903, -43.1727, 
        -43.16127, -43.14766, -43.13249, -43.11784, -43.10499, -43.09449, 
        -43.08599, -43.07857, -43.07055, -43.06017, -43.04598, -43.02658, 
        -43.00089, -42.97022, -42.93624, -42.9005, -42.86369, -42.8269, 
        -42.79049, -42.75456, -42.7183, -42.68098, -42.64135, -42.59817, 
        -42.55402, -42.50834, -42.46223, -42.41697, -42.37388, -42.33479, 
        -42.3003, -42.27149, -42.24781, -42.22832, -42.21302, -42.20266, 
        -42.19685, -42.19562, -42.19796, -42.20308, -42.20921, -42.21514, 
        -42.21947, -42.22124, -42.21994, -42.21667, -42.21115, -42.20618, 
        -42.2019, -42.20058, -42.20093, -42.20303, -42.20481, -42.20632, 
        -42.20728, -42.20837, -42.211, -42.21674, -42.22722, -42.24484, 
        -42.27168, -42.30875, -42.35567, -42.41057, -42.47015, -42.53031, 
        -42.58722, -42.63764, -42.68024, -42.7142, -42.74034, -42.76037, 
        -42.77631, -42.78976, -42.80244, -42.81337, -42.82486, -42.83496, 
        -42.84309, -42.84807, -42.85065, -42.85154, -42.85205, -42.85263, 
        -42.85417, -42.8544, -42.85257, -42.84644, -42.83469, -42.81583, 
        -42.78769, -42.75142, -42.70879, -42.66322, -42.61739, -42.57288, 
        -42.52972, -42.48712, -42.44157, -42.38847, -42.32431, -42.24501, 
        -42.15091, -42.04234, -41.92339, -41.79972, -41.67759, -41.56326, 
        -41.46148, -41.37889, -41.31368, -41.27286, -41.2514, -41.24559, 
        -41.25133, -41.26632, -41.28326, -41.30235, -41.32392, -41.34798, 
        -41.37891, -41.41012, -41.44596, -41.48587, -41.5314, -41.5794, 
        -41.63647, -41.69955, -41.7719, -41.85225, -41.94147, -42.03624, 
        -42.13359, -42.22805, -42.31586, -42.39539, -42.46423, -42.52211, 
        -42.56957, -42.60739, -42.63516, -42.65255, -42.65929, -42.65348, 
        -42.63257, -42.59425, -42.53665, -42.45796, -42.35825, -42.23802, 
        -42.10303, -41.95721, -41.80748, -41.66104, -41.52388, -41.40098, 
        -41.2944, -41.20479, -41.13161, -41.07437, -41.03037, -40.99774, 
        -40.97368,
  -41.1088, -41.14439, -41.17704, -41.2076, -41.23694, -41.26623, 
        -41.29625, -41.32743, -41.36058, -41.39573, -41.43363, -41.47332, 
        -41.51708, -41.56429, -41.61374, -41.66478, -41.71772, -41.77129, 
        -41.82571, -41.88012, -41.93481, -41.99033, -42.04723, -42.10664, 
        -42.16856, -42.23384, -42.30116, -42.37239, -42.44608, -42.52129, 
        -42.59616, -42.66936, -42.73943, -42.80603, -42.86814, -42.92596, 
        -42.97941, -43.02837, -43.07397, -43.11549, -43.15317, -43.18614, 
        -43.21687, -43.24461, -43.26955, -43.29206, -43.3132, -43.33296, 
        -43.35178, -43.36965, -43.38599, -43.40073, -43.41241, -43.42144, 
        -43.42739, -43.42911, -43.42693, -43.41945, -43.40949, -43.39701, 
        -43.38213, -43.36575, -43.34811, -43.32978, -43.3112, -43.29235, 
        -43.27447, -43.25639, -43.2373, -43.21698, -43.19512, -43.17276, 
        -43.15107, -43.13136, -43.11303, -43.09809, -43.08564, -43.0756, 
        -43.06799, -43.06266, -43.0599, -43.0595, -43.06165, -43.06592, 
        -43.07132, -43.07776, -43.08501, -43.09335, -43.10221, -43.11069, 
        -43.11728, -43.12077, -43.11976, -43.11577, -43.10734, -43.0938, 
        -43.07471, -43.05008, -43.01916, -42.98203, -42.93871, -42.88975, 
        -42.83623, -42.77986, -42.72337, -42.66913, -42.62045, -42.58091, 
        -42.55293, -42.53875, -42.54032, -42.55669, -42.58753, -42.62976, 
        -42.67968, -42.73381, -42.78963, -42.84534, -42.89972, -42.95176, 
        -43.00035, -43.04507, -43.08576, -43.1221, -43.15355, -43.17939, 
        -43.20054, -43.2177, -43.23212, -43.24515, -43.25661, -43.26594, 
        -43.27501, -43.28259, -43.28852, -43.2916, -43.29094, -43.28576, 
        -43.27692, -43.26537, -43.25248, -43.23997, -43.22919, -43.22061, 
        -43.21391, -43.20803, -43.20137, -43.19252, -43.1799, -43.16195, 
        -43.13831, -43.10996, -43.07893, -43.04563, -43.01303, -42.98039, 
        -42.94793, -42.91563, -42.88305, -42.8491, -42.81308, -42.77495, 
        -42.73512, -42.6936, -42.65144, -42.60997, -42.57011, -42.53314, 
        -42.50009, -42.47139, -42.44607, -42.42432, -42.40636, -42.39217, 
        -42.3827, -42.37777, -42.37672, -42.37793, -42.38188, -42.3863, 
        -42.38976, -42.39076, -42.38873, -42.3834, -42.37533, -42.36572, 
        -42.35548, -42.34515, -42.33505, -42.32503, -42.31462, -42.30402, 
        -42.29386, -42.28503, -42.27852, -42.27657, -42.28054, -42.2923, 
        -42.31371, -42.3452, -42.38606, -42.43398, -42.48575, -42.53744, 
        -42.58485, -42.62683, -42.66156, -42.6888, -42.70966, -42.72556, 
        -42.73817, -42.74866, -42.75814, -42.76683, -42.77442, -42.78108, 
        -42.78606, -42.78892, -42.79006, -42.7897, -42.78917, -42.78916, 
        -42.78942, -42.78886, -42.78559, -42.77871, -42.76633, -42.74686, 
        -42.71953, -42.68522, -42.6465, -42.60571, -42.56503, -42.5258, 
        -42.48628, -42.4466, -42.40279, -42.35057, -42.28603, -42.20695, 
        -42.11311, -42.00615, -41.88968, -41.77003, -41.65158, -41.54285, 
        -41.44802, -41.37213, -41.31456, -41.27997, -41.26562, -41.26806, 
        -41.28229, -41.30531, -41.33185, -41.36085, -41.39288, -41.42636, 
        -41.46479, -41.50212, -41.54188, -41.58457, -41.63122, -41.67904, 
        -41.73344, -41.79567, -41.86301, -41.93955, -42.02367, -42.11367, 
        -42.20622, -42.2965, -42.38025, -42.4572, -42.52396, -42.58045, 
        -42.62707, -42.66376, -42.6906, -42.70675, -42.71169, -42.70366, 
        -42.68, -42.63886, -42.57832, -42.49706, -42.39495, -42.27341, 
        -42.13612, -41.98755, -41.83424, -41.68268, -41.5387, -41.40711, 
        -41.29155, -41.19124, -41.1078, -41.04015, -40.98667, -40.94474, 
        -40.91304,
  -41.14437, -41.18065, -41.21433, -41.24653, -41.27808, -41.30976, 
        -41.34097, -41.37434, -41.40907, -41.44574, -41.48484, -41.52649, 
        -41.571, -41.61824, -41.66774, -41.71892, -41.77102, -41.82383, 
        -41.87688, -41.9298, -41.98256, -42.03483, -42.08927, -42.14567, 
        -42.20469, -42.26641, -42.33097, -42.39924, -42.4702, -42.54236, 
        -42.61448, -42.68471, -42.75155, -42.81415, -42.87231, -42.92635, 
        -42.97567, -43.02245, -43.0658, -43.10543, -43.14122, -43.1734, 
        -43.20203, -43.22778, -43.25063, -43.27107, -43.28972, -43.30725, 
        -43.32389, -43.33964, -43.35419, -43.36737, -43.37761, -43.38623, 
        -43.39167, -43.39314, -43.39066, -43.38419, -43.37413, -43.3615, 
        -43.34692, -43.33095, -43.31445, -43.29724, -43.27988, -43.26267, 
        -43.24593, -43.22909, -43.21127, -43.19043, -43.16926, -43.14702, 
        -43.12493, -43.10417, -43.08552, -43.0695, -43.05623, -43.04604, 
        -43.03873, -43.03426, -43.03276, -43.03391, -43.03735, -43.04304, 
        -43.04972, -43.05736, -43.06506, -43.07493, -43.08569, -43.09603, 
        -43.10476, -43.11065, -43.1133, -43.11219, -43.10676, -43.09666, 
        -43.08092, -43.05944, -43.03223, -42.99895, -42.95962, -42.91492, 
        -42.86594, -42.81436, -42.76239, -42.71165, -42.66738, -42.63254, 
        -42.60938, -42.60064, -42.60786, -42.63134, -42.66887, -42.71775, 
        -42.77376, -42.83323, -42.89326, -42.95185, -43.00767, -43.05995, 
        -43.10763, -43.15092, -43.18988, -43.22448, -43.25322, -43.27855, 
        -43.29926, -43.31665, -43.33158, -43.34485, -43.35623, -43.36598, 
        -43.37457, -43.38156, -43.38713, -43.39051, -43.39056, -43.38729, 
        -43.38064, -43.37161, -43.3614, -43.3513, -43.34268, -43.33596, 
        -43.33081, -43.32497, -43.31932, -43.31145, -43.29964, -43.28284, 
        -43.26099, -43.23488, -43.20663, -43.17776, -43.14899, -43.12037, 
        -43.09159, -43.06301, -43.03381, -43.00336, -42.97082, -42.93679, 
        -42.90139, -42.86428, -42.8269, -42.78967, -42.75381, -42.72009, 
        -42.68909, -42.66007, -42.63448, -42.61135, -42.59086, -42.57372, 
        -42.56069, -42.55192, -42.54741, -42.54623, -42.54743, -42.54976, 
        -42.55163, -42.5516, -42.54857, -42.54198, -42.5317, -42.51813, 
        -42.50215, -42.48458, -42.46592, -42.44636, -42.4262, -42.40605, 
        -42.38679, -42.36988, -42.35479, -42.34562, -42.34404, -42.35044, 
        -42.36651, -42.3922, -42.42706, -42.46815, -42.51264, -42.55672, 
        -42.5972, -42.63165, -42.65924, -42.68005, -42.69549, -42.70677, 
        -42.71517, -42.72199, -42.72768, -42.73231, -42.73568, -42.73842, 
        -42.74053, -42.74156, -42.74156, -42.74081, -42.74, -42.73975, 
        -42.73932, -42.73676, -42.73278, -42.72525, -42.71248, -42.69292, 
        -42.66685, -42.63526, -42.60026, -42.56423, -42.52846, -42.4936, 
        -42.4586, -42.42142, -42.37921, -42.32759, -42.26352, -42.18564, 
        -42.0939, -41.99063, -41.87923, -41.76501, -41.65287, -41.55085, 
        -41.46386, -41.395, -41.34456, -41.31677, -41.30841, -41.31701, 
        -41.33724, -41.36578, -41.39861, -41.43582, -41.47403, -41.5142, 
        -41.55558, -41.59681, -41.63861, -41.6823, -41.72783, -41.77584, 
        -41.82798, -41.88625, -41.95087, -42.02341, -42.1031, -42.18847, 
        -42.27628, -42.36263, -42.44458, -42.51894, -42.58363, -42.63886, 
        -42.68447, -42.72067, -42.74642, -42.76137, -42.76496, -42.75467, 
        -42.72876, -42.68539, -42.6229, -42.54018, -42.43741, -42.31581, 
        -42.17855, -42.03002, -41.87548, -41.72086, -41.57159, -41.43253, 
        -41.3073, -41.1971, -41.1019, -41.02295, -40.95773, -40.90583, 
        -40.86476,
  -41.17487, -41.21115, -41.24608, -41.28002, -41.3136, -41.3476, 
        -41.38225, -41.41785, -41.45443, -41.4926, -41.53268, -41.57503, 
        -41.62005, -41.66759, -41.71704, -41.76783, -41.8182, -41.8701, 
        -41.9218, -41.97313, -42.02402, -42.07527, -42.1273, -42.18081, 
        -42.23674, -42.29516, -42.35643, -42.42114, -42.48854, -42.5573, 
        -42.62603, -42.69187, -42.75538, -42.81449, -42.86925, -42.92012, 
        -42.96738, -43.01173, -43.05316, -43.0913, -43.12538, -43.15581, 
        -43.1827, -43.20648, -43.22745, -43.24596, -43.26154, -43.27689, 
        -43.29123, -43.3049, -43.31751, -43.32905, -43.33899, -43.3467, 
        -43.35136, -43.35219, -43.34957, -43.34317, -43.33327, -43.32107, 
        -43.30743, -43.29249, -43.277, -43.26008, -43.24397, -43.22831, 
        -43.21227, -43.19631, -43.17905, -43.16012, -43.1398, -43.11796, 
        -43.09572, -43.07442, -43.05499, -43.03807, -43.02438, -43.0139, 
        -43.00696, -43.00337, -43.00174, -43.00406, -43.00897, -43.01563, 
        -43.02342, -43.03222, -43.04195, -43.05316, -43.06527, -43.07722, 
        -43.0878, -43.09616, -43.10151, -43.10333, -43.10081, -43.09373, 
        -43.08142, -43.06365, -43.03962, -43.01118, -42.97728, -42.93843, 
        -42.89566, -42.85021, -42.80438, -42.76047, -42.72181, -42.69173, 
        -42.67367, -42.67018, -42.68244, -42.71076, -42.75339, -42.80678, 
        -42.86691, -42.92985, -42.99216, -43.05098, -43.10685, -43.15818, 
        -43.20441, -43.24544, -43.28191, -43.31431, -43.34258, -43.3668, 
        -43.38728, -43.40472, -43.41977, -43.43298, -43.44415, -43.45347, 
        -43.46133, -43.46812, -43.47363, -43.47736, -43.47861, -43.47706, 
        -43.47179, -43.46568, -43.45822, -43.45071, -43.44418, -43.43904, 
        -43.43494, -43.43093, -43.42576, -43.41817, -43.40678, -43.39092, 
        -43.37072, -43.34709, -43.32158, -43.29594, -43.27079, -43.24558, 
        -43.2201, -43.19474, -43.16862, -43.14149, -43.11282, -43.08163, 
        -43.05025, -43.01801, -42.98524, -42.95263, -42.92081, -42.89066, 
        -42.86234, -42.83583, -42.81072, -42.78697, -42.76502, -42.74576, 
        -42.72979, -42.71778, -42.70982, -42.70539, -42.70358, -42.70364, 
        -42.70372, -42.70224, -42.69817, -42.69006, -42.67808, -42.66061, 
        -42.64062, -42.6179, -42.5931, -42.56694, -42.53971, -42.51279, 
        -42.48713, -42.46373, -42.44379, -42.42906, -42.42141, -42.42236, 
        -42.43297, -42.45317, -42.48166, -42.51599, -42.55326, -42.58996, 
        -42.62309, -42.65048, -42.67134, -42.68608, -42.69605, -42.70246, 
        -42.70636, -42.70849, -42.70993, -42.70892, -42.70862, -42.70802, 
        -42.70763, -42.70712, -42.70686, -42.70631, -42.70614, -42.70597, 
        -42.70524, -42.7032, -42.69871, -42.69077, -42.67755, -42.65832, 
        -42.63331, -42.60412, -42.57249, -42.54035, -42.50872, -42.47744, 
        -42.44524, -42.40983, -42.36862, -42.31791, -42.25549, -42.17968, 
        -42.09157, -41.99324, -41.88816, -41.78145, -41.67742, -41.58242, 
        -41.50201, -41.4397, -41.39611, -41.37375, -41.36961, -41.38064, 
        -41.40468, -41.43663, -41.47389, -41.51552, -41.55922, -41.60404, 
        -41.64966, -41.69381, -41.73729, -41.78054, -41.82512, -41.87139, 
        -41.92267, -41.97849, -42.04051, -42.1094, -42.18464, -42.26532, 
        -42.34852, -42.43103, -42.50924, -42.5808, -42.64369, -42.6976, 
        -42.74195, -42.77681, -42.80137, -42.81532, -42.81731, -42.80521, 
        -42.77729, -42.73201, -42.6683, -42.5854, -42.48237, -42.3624, 
        -42.22721, -42.08056, -41.92697, -41.77146, -41.61891, -41.47384, 
        -41.33975, -41.21892, -41.11243, -41.02083, -40.94341, -40.87941, 
        -40.82757,
  -41.19893, -41.23717, -41.27339, -41.30912, -41.3451, -41.38166, 
        -41.41888, -41.45672, -41.49515, -41.53451, -41.57533, -41.61721, 
        -41.6625, -41.71004, -41.7592, -41.80933, -41.85987, -41.91044, 
        -41.96101, -42.01084, -42.06005, -42.1095, -42.15966, -42.2107, 
        -42.26357, -42.31892, -42.37615, -42.43743, -42.50128, -42.56654, 
        -42.63147, -42.69464, -42.75454, -42.81046, -42.86223, -42.91003, 
        -42.9548, -42.99665, -43.03585, -43.07204, -43.10435, -43.13187, 
        -43.15707, -43.179, -43.19861, -43.21529, -43.23025, -43.24373, 
        -43.25603, -43.26758, -43.27812, -43.2876, -43.29586, -43.30212, 
        -43.30584, -43.30605, -43.30304, -43.2957, -43.28651, -43.27528, 
        -43.26288, -43.24936, -43.23508, -43.22041, -43.20541, -43.19013, 
        -43.17442, -43.15865, -43.14195, -43.12405, -43.10444, -43.08387, 
        -43.06231, -43.04128, -43.02078, -43.00388, -42.99019, -42.97999, 
        -42.97349, -42.97072, -42.97106, -42.97441, -42.97987, -42.98732, 
        -42.99594, -43.00586, -43.01687, -43.02903, -43.04208, -43.05547, 
        -43.06788, -43.0784, -43.08554, -43.08999, -43.0906, -43.08619, 
        -43.07699, -43.06297, -43.04457, -43.02182, -42.99446, -42.96279, 
        -42.92749, -42.88984, -42.8516, -42.81452, -42.7818, -42.75704, 
        -42.7438, -42.745, -42.76138, -42.79192, -42.8374, -42.89308, 
        -42.9552, -43.01938, -43.08231, -43.14197, -43.19696, -43.24672, 
        -43.29076, -43.32948, -43.36341, -43.39346, -43.42029, -43.44355, 
        -43.46389, -43.48153, -43.4968, -43.50985, -43.52074, -43.5286, 
        -43.53607, -43.54241, -43.54786, -43.55212, -43.55451, -43.55473, 
        -43.55296, -43.54964, -43.54498, -43.53984, -43.53514, -43.53124, 
        -43.52785, -43.52411, -43.51885, -43.51121, -43.50006, -43.48501, 
        -43.46634, -43.44503, -43.42245, -43.39886, -43.3767, -43.35472, 
        -43.33234, -43.30941, -43.28587, -43.26162, -43.23637, -43.20977, 
        -43.18254, -43.15463, -43.12642, -43.09845, -43.07096, -43.0445, 
        -43.01926, -42.9951, -42.97128, -42.94813, -42.92576, -42.90527, 
        -42.88733, -42.87288, -42.86195, -42.85348, -42.84906, -42.84655, 
        -42.84466, -42.84187, -42.83662, -42.82764, -42.81445, -42.79655, 
        -42.77423, -42.74869, -42.72041, -42.69012, -42.65898, -42.62819, 
        -42.59848, -42.57061, -42.54601, -42.52645, -42.51323, -42.5084, 
        -42.51319, -42.52717, -42.54881, -42.57609, -42.60598, -42.63433, 
        -42.66035, -42.68108, -42.69555, -42.70417, -42.70847, -42.70979, 
        -42.70909, -42.7072, -42.70404, -42.69991, -42.69568, -42.69225, 
        -42.69039, -42.68944, -42.68938, -42.69038, -42.69135, -42.69188, 
        -42.69128, -42.68914, -42.68449, -42.67583, -42.66239, -42.643, 
        -42.61861, -42.59128, -42.56236, -42.53336, -42.50456, -42.47585, 
        -42.44422, -42.41002, -42.36953, -42.31992, -42.25955, -42.18705, 
        -42.10409, -42.01242, -41.91521, -41.81714, -41.72316, -41.63791, 
        -41.56552, -41.51014, -41.4718, -41.45333, -41.45206, -41.46508, 
        -41.48998, -41.52325, -41.56303, -41.60796, -41.65427, -41.70075, 
        -41.74823, -41.7938, -41.83772, -41.88062, -41.92406, -41.96899, 
        -42.01808, -42.07217, -42.13182, -42.19755, -42.26918, -42.34532, 
        -42.42407, -42.50115, -42.57557, -42.64362, -42.70403, -42.75575, 
        -42.79831, -42.83139, -42.85432, -42.867, -42.86704, -42.85299, 
        -42.823, -42.77613, -42.71178, -42.6295, -42.52935, -42.41262, 
        -42.28119, -42.13836, -41.98785, -41.83337, -41.67937, -41.52961, 
        -41.38776, -41.25676, -41.13844, -41.03387, -40.94324, -40.86619, 
        -40.80252,
  -41.21912, -41.25853, -41.29655, -41.334, -41.37213, -41.4109, 
        -41.44924, -41.48899, -41.52883, -41.56923, -41.61084, -41.65427, 
        -41.70003, -41.74753, -41.79631, -41.84563, -41.89531, -41.94488, 
        -41.99341, -42.04198, -42.09024, -42.13719, -42.1848, -42.23368, 
        -42.28428, -42.33682, -42.3921, -42.45027, -42.51053, -42.57205, 
        -42.63317, -42.69282, -42.74933, -42.80235, -42.85136, -42.89674, 
        -42.93775, -42.9768, -43.01327, -43.047, -43.07733, -43.10393, 
        -43.12735, -43.14766, -43.16573, -43.181, -43.1948, -43.20662, 
        -43.21721, -43.22673, -43.2352, -43.24242, -43.24782, -43.25254, 
        -43.25484, -43.2543, -43.25087, -43.24456, -43.23627, -43.22606, 
        -43.21469, -43.20238, -43.18928, -43.17552, -43.16115, -43.14632, 
        -43.1312, -43.11547, -43.09839, -43.08112, -43.06279, -43.04342, 
        -43.02346, -43.00371, -42.98526, -42.96912, -42.95623, -42.94685, 
        -42.94134, -42.93957, -42.94099, -42.94514, -42.95147, -42.95967, 
        -42.96924, -42.97999, -42.99073, -43.0037, -43.01751, -43.03197, 
        -43.04585, -43.05855, -43.06891, -43.07593, -43.0788, -43.0772, 
        -43.07109, -43.06117, -43.04768, -43.03101, -43.01075, -42.98697, 
        -42.96011, -42.93104, -42.89976, -42.87028, -42.84414, -42.82515, 
        -42.81682, -42.82195, -42.84092, -42.87424, -42.92059, -42.97663, 
        -43.03851, -43.10209, -43.16416, -43.22254, -43.27597, -43.32388, 
        -43.36586, -43.40217, -43.43397, -43.46235, -43.48682, -43.50959, 
        -43.52985, -43.54767, -43.56324, -43.5764, -43.58715, -43.59574, 
        -43.60283, -43.60903, -43.6146, -43.61941, -43.623, -43.62514, 
        -43.62558, -43.62459, -43.62223, -43.61914, -43.61581, -43.61253, 
        -43.60919, -43.60404, -43.59832, -43.59029, -43.57914, -43.56516, 
        -43.54832, -43.52933, -43.50953, -43.48977, -43.47041, -43.4513, 
        -43.43138, -43.41099, -43.3898, -43.36814, -43.34564, -43.3227, 
        -43.29905, -43.27522, -43.25125, -43.22739, -43.20398, -43.1813, 
        -43.15829, -43.13688, -43.11494, -43.09306, -43.07121, -43.05054, 
        -43.03152, -43.01565, -43.00295, -42.99376, -42.98717, -42.98222, 
        -42.97824, -42.97369, -42.96696, -42.95701, -42.94312, -42.92466, 
        -42.90176, -42.87517, -42.84552, -42.81397, -42.78131, -42.74884, 
        -42.71707, -42.68668, -42.65792, -42.63417, -42.61633, -42.60609, 
        -42.60456, -42.61164, -42.62595, -42.64557, -42.66804, -42.69, 
        -42.70915, -42.72338, -42.7319, -42.73524, -42.73446, -42.731, 
        -42.72604, -42.71997, -42.71319, -42.7058, -42.69865, -42.69309, 
        -42.6899, -42.6888, -42.69001, -42.6923, -42.69469, -42.69615, 
        -42.69617, -42.69299, -42.68777, -42.67858, -42.66443, -42.64531, 
        -42.62154, -42.59496, -42.56713, -42.5399, -42.51339, -42.48617, 
        -42.45671, -42.42356, -42.38419, -42.33631, -42.27847, -42.21004, 
        -42.13255, -42.0482, -41.95972, -41.87154, -41.78723, -41.71165, 
        -41.64814, -41.59917, -41.56621, -41.55033, -41.55039, -41.56438, 
        -41.58945, -41.62269, -41.66328, -41.70824, -41.75572, -41.80289, 
        -41.85095, -41.89672, -41.94092, -41.98337, -42.02556, -42.06953, 
        -42.11687, -42.16909, -42.22614, -42.28847, -42.35619, -42.42802, 
        -42.50135, -42.57467, -42.64455, -42.70864, -42.76558, -42.81454, 
        -42.85472, -42.88548, -42.90644, -42.91718, -42.91511, -42.89852, 
        -42.86662, -42.81862, -42.75413, -42.67271, -42.57529, -42.46242, 
        -42.33579, -42.19802, -42.05173, -41.90011, -41.7464, -41.59352, 
        -41.44561, -41.30528, -41.17598, -41.05913, -40.9551, -40.86491, 
        -40.78859,
  -41.2351, -41.27497, -41.31454, -41.35393, -41.39392, -41.43447, 
        -41.47543, -41.51661, -41.55762, -41.59893, -41.64135, -41.68522, 
        -41.73101, -41.77856, -41.8268, -41.87586, -41.9235, -41.97168, 
        -42.01907, -42.06641, -42.11311, -42.15926, -42.20535, -42.25256, 
        -42.3008, -42.35098, -42.40374, -42.45876, -42.5156, -42.57327, 
        -42.63086, -42.6859, -42.73958, -42.78989, -42.83623, -42.8787, 
        -42.91782, -42.95414, -42.98795, -43.01897, -43.04696, -43.07132, 
        -43.09283, -43.11174, -43.12775, -43.14205, -43.15366, -43.16434, 
        -43.17341, -43.18109, -43.18737, -43.19256, -43.19698, -43.19997, 
        -43.2007, -43.19923, -43.19516, -43.18933, -43.18174, -43.17249, 
        -43.16211, -43.15067, -43.13833, -43.12416, -43.11045, -43.09602, 
        -43.0812, -43.06564, -43.05014, -43.03415, -43.01729, -42.99968, 
        -42.9818, -42.96403, -42.94756, -42.93306, -42.92159, -42.91388, 
        -42.90963, -42.90895, -42.91055, -42.91586, -42.92335, -42.93243, 
        -42.9431, -42.95467, -42.96709, -42.98045, -42.99488, -43.01004, 
        -43.02533, -43.0396, -43.05185, -43.06065, -43.06571, -43.0666, 
        -43.06382, -43.05798, -43.04871, -43.03811, -43.02504, -43.00914, 
        -42.99077, -42.97043, -42.94832, -42.92677, -42.90785, -42.89474, 
        -42.89072, -42.89874, -42.92003, -42.9534, -42.99848, -43.05288, 
        -43.11298, -43.17476, -43.23489, -43.29027, -43.34172, -43.38751, 
        -43.42742, -43.4621, -43.49236, -43.51937, -43.54414, -43.56674, 
        -43.58719, -43.60546, -43.62138, -43.63481, -43.64561, -43.65421, 
        -43.66127, -43.66752, -43.67355, -43.67906, -43.6838, -43.68752, 
        -43.68874, -43.6897, -43.68925, -43.68751, -43.68493, -43.68172, 
        -43.6778, -43.67284, -43.66628, -43.65781, -43.64705, -43.63428, 
        -43.61929, -43.60283, -43.58561, -43.56873, -43.55199, -43.53524, 
        -43.51769, -43.49971, -43.4808, -43.46146, -43.44058, -43.42045, 
        -43.40034, -43.3798, -43.3597, -43.33975, -43.32027, -43.3013, 
        -43.28267, -43.26394, -43.24461, -43.22458, -43.20406, -43.1838, 
        -43.16521, -43.14866, -43.13535, -43.12445, -43.11668, -43.11028, 
        -43.10434, -43.09769, -43.08951, -43.07877, -43.06448, -43.04502, 
        -43.02245, -42.99647, -42.96713, -42.93647, -42.90415, -42.87188, 
        -42.83978, -42.80839, -42.77864, -42.752, -42.7299, -42.7146, 
        -42.70678, -42.70669, -42.71312, -42.72497, -42.73941, -42.75399, 
        -42.76632, -42.77447, -42.77766, -42.77617, -42.77139, -42.76402, 
        -42.75556, -42.74634, -42.7355, -42.72552, -42.71661, -42.70976, 
        -42.70564, -42.70503, -42.70707, -42.71035, -42.7142, -42.71612, 
        -42.71685, -42.71455, -42.70903, -42.69908, -42.68415, -42.66417, 
        -42.6402, -42.61364, -42.58667, -42.56041, -42.53478, -42.50861, 
        -42.48051, -42.44854, -42.4106, -42.36507, -42.31029, -42.24648, 
        -42.17514, -42.09842, -42.01888, -41.94069, -41.86696, -41.8003, 
        -41.74522, -41.70316, -41.67503, -41.66137, -41.66217, -41.67612, 
        -41.70007, -41.73238, -41.77209, -41.81655, -41.86359, -41.91173, 
        -41.95944, -42.00491, -42.04871, -42.09032, -42.13128, -42.17414, 
        -42.21985, -42.27049, -42.32467, -42.38383, -42.44769, -42.51412, 
        -42.58219, -42.64987, -42.7146, -42.77411, -42.82704, -42.87265, 
        -42.90959, -42.93725, -42.95589, -42.96359, -42.95921, -42.9406, 
        -42.90674, -42.85783, -42.79329, -42.71331, -42.61748, -42.50858, 
        -42.38677, -42.25435, -42.11293, -41.96483, -41.81247, -41.65875, 
        -41.50598, -41.35888, -41.22064, -41.0919, -40.97555, -40.87251, 
        -40.78374,
  -41.24626, -41.28898, -41.33036, -41.37142, -41.41295, -41.45485, 
        -41.49714, -41.53916, -41.58094, -41.62289, -41.66559, -41.70874, 
        -41.75447, -41.80175, -41.84973, -41.89776, -41.94556, -41.99269, 
        -42.03912, -42.08496, -42.1304, -42.17533, -42.22025, -42.26553, 
        -42.31196, -42.36019, -42.40961, -42.46177, -42.51545, -42.56963, 
        -42.62392, -42.67676, -42.72729, -42.77495, -42.81861, -42.85838, 
        -42.89479, -42.92803, -42.95881, -42.98679, -43.01209, -43.03317, 
        -43.05255, -43.06956, -43.08414, -43.09728, -43.1086, -43.11852, 
        -43.12639, -43.13261, -43.13733, -43.14066, -43.1429, -43.14383, 
        -43.14327, -43.14046, -43.13615, -43.12938, -43.12225, -43.11369, 
        -43.10394, -43.09296, -43.08126, -43.06866, -43.05542, -43.04126, 
        -43.02686, -43.01208, -42.99714, -42.98249, -42.96751, -42.95218, 
        -42.93685, -42.92194, -42.90688, -42.89492, -42.88552, -42.87958, 
        -42.87698, -42.87782, -42.88191, -42.88874, -42.89753, -42.9079, 
        -42.91955, -42.93203, -42.94507, -42.95898, -42.97381, -42.98975, 
        -43.00598, -43.0214, -43.03398, -43.04451, -43.05135, -43.05461, 
        -43.05498, -43.05328, -43.05001, -43.0453, -43.03894, -43.03072, 
        -43.02047, -43.00827, -42.99459, -42.9808, -42.96901, -42.9616, 
        -42.96174, -42.97209, -42.99359, -43.02544, -43.06837, -43.11983, 
        -43.17682, -43.2355, -43.29277, -43.34669, -43.39584, -43.43959, 
        -43.47806, -43.51129, -43.54081, -43.56727, -43.59163, -43.61438, 
        -43.63536, -43.65416, -43.67057, -43.68439, -43.69557, -43.70343, 
        -43.71079, -43.71744, -43.72394, -43.73022, -43.73602, -43.74099, 
        -43.74479, -43.74735, -43.74828, -43.74721, -43.74487, -43.74129, 
        -43.7367, -43.73053, -43.72301, -43.71413, -43.70389, -43.69238, 
        -43.67955, -43.66551, -43.65015, -43.63576, -43.62162, -43.6073, 
        -43.59225, -43.57654, -43.56002, -43.54295, -43.5257, -43.50792, 
        -43.49035, -43.47321, -43.45644, -43.44013, -43.42406, -43.40853, 
        -43.3931, -43.37729, -43.36054, -43.34267, -43.32384, -43.3051, 
        -43.28743, -43.27153, -43.25702, -43.24596, -43.23697, -43.22939, 
        -43.22182, -43.2135, -43.20385, -43.19203, -43.17751, -43.1594, 
        -43.13787, -43.11338, -43.08589, -43.05703, -43.02667, -42.99563, 
        -42.96432, -42.93314, -42.9027, -42.87396, -42.84885, -42.82887, 
        -42.81523, -42.80801, -42.80682, -42.81042, -42.81721, -42.82356, 
        -42.82907, -42.83167, -42.83014, -42.82479, -42.81664, -42.80646, 
        -42.79543, -42.78388, -42.77219, -42.76086, -42.75078, -42.74331, 
        -42.73938, -42.73866, -42.74107, -42.74513, -42.74955, -42.75249, 
        -42.75331, -42.75122, -42.74465, -42.73345, -42.7174, -42.69629, 
        -42.67158, -42.64479, -42.61765, -42.59146, -42.56618, -42.53991, 
        -42.51284, -42.48237, -42.44673, -42.40391, -42.35302, -42.2942, 
        -42.2293, -42.16024, -42.0896, -42.02109, -41.95744, -41.90137, 
        -41.8547, -41.81915, -41.79573, -41.78471, -41.78571, -41.79891, 
        -41.82159, -41.85264, -41.89107, -41.93452, -41.98055, -42.02767, 
        -42.07453, -42.11921, -42.16151, -42.20191, -42.24178, -42.2823, 
        -42.32582, -42.37344, -42.42529, -42.48049, -42.53925, -42.60044, 
        -42.6619, -42.72379, -42.78284, -42.83727, -42.88557, -42.9268, 
        -42.95992, -42.98457, -42.99997, -43.00502, -42.99786, -42.97708, 
        -42.94179, -42.8919, -42.82731, -42.74833, -42.65585, -42.55051, 
        -42.43354, -42.30568, -42.16902, -42.02481, -41.87501, -41.72141, 
        -41.56698, -41.41534, -41.26972, -41.13203, -41.00507, -40.89051, 
        -40.78985,
  -41.25523, -41.29985, -41.34321, -41.38605, -41.42902, -41.47209, 
        -41.514, -41.55645, -41.59865, -41.64091, -41.68369, -41.72771, 
        -41.77338, -41.81998, -41.86746, -41.91479, -41.96168, -42.00788, 
        -42.05334, -42.09826, -42.1415, -42.18544, -42.22921, -42.27296, 
        -42.31754, -42.3639, -42.41188, -42.46146, -42.51228, -42.56338, 
        -42.61421, -42.66397, -42.71172, -42.75658, -42.79783, -42.83467, 
        -42.86726, -42.89756, -42.92532, -42.94998, -42.97232, -42.99198, 
        -43.00915, -43.0242, -43.03734, -43.0493, -43.05961, -43.06853, 
        -43.07562, -43.08089, -43.08426, -43.08596, -43.08506, -43.0841, 
        -43.08176, -43.0779, -43.07303, -43.06697, -43.06022, -43.05207, 
        -43.04254, -43.0317, -43.02073, -43.00856, -42.99565, -42.98223, 
        -42.96854, -42.95491, -42.94021, -42.92714, -42.9141, -42.90137, 
        -42.88876, -42.87708, -42.86596, -42.8567, -42.84971, -42.84565, 
        -42.84501, -42.84776, -42.85339, -42.86183, -42.87249, -42.88439, 
        -42.89748, -42.91121, -42.92386, -42.93838, -42.95401, -42.97029, 
        -42.98714, -43.00364, -43.01809, -43.0296, -43.03798, -43.04346, 
        -43.04683, -43.04905, -43.0506, -43.05114, -43.05082, -43.04926, 
        -43.04632, -43.04154, -43.03461, -43.02845, -43.02342, -43.0217, 
        -43.0258, -43.03775, -43.05931, -43.0904, -43.13059, -43.17849, 
        -43.23156, -43.28656, -43.3405, -43.39149, -43.43833, -43.48036, 
        -43.51732, -43.55012, -43.57892, -43.60545, -43.62904, -43.65213, 
        -43.67354, -43.69284, -43.7099, -43.72425, -43.73583, -43.74522, 
        -43.75338, -43.76074, -43.76799, -43.77503, -43.78164, -43.78762, 
        -43.79261, -43.79612, -43.7979, -43.7975, -43.79501, -43.79086, 
        -43.78534, -43.77711, -43.7688, -43.75979, -43.75014, -43.74002, 
        -43.72948, -43.71834, -43.70658, -43.69486, -43.68321, -43.67127, 
        -43.65867, -43.64534, -43.63116, -43.61615, -43.60079, -43.58565, 
        -43.57061, -43.55615, -43.54254, -43.52926, -43.51643, -43.50397, 
        -43.49058, -43.47743, -43.46327, -43.44754, -43.43085, -43.41389, 
        -43.39786, -43.38314, -43.3704, -43.35947, -43.35004, -43.34159, 
        -43.33274, -43.32292, -43.31198, -43.2992, -43.28444, -43.26689, 
        -43.24656, -43.22381, -43.19868, -43.17183, -43.14418, -43.11536, 
        -43.08555, -43.0544, -43.02371, -42.99388, -42.96675, -42.94316, 
        -42.92442, -42.91114, -42.90284, -42.89889, -42.89812, -42.89846, 
        -42.89804, -42.89519, -42.88992, -42.88172, -42.87119, -42.85918, 
        -42.84666, -42.83372, -42.82093, -42.80918, -42.79932, -42.79155, 
        -42.78765, -42.7868, -42.78909, -42.79314, -42.79734, -42.80037, 
        -42.80006, -42.79712, -42.78952, -42.77691, -42.75952, -42.73729, 
        -42.71162, -42.68405, -42.65633, -42.62981, -42.60474, -42.58024, 
        -42.55447, -42.52604, -42.49285, -42.45324, -42.40659, -42.35331, 
        -42.29483, -42.23322, -42.1713, -42.11177, -42.0572, -42.01014, 
        -41.97198, -41.94294, -41.92355, -41.91496, -41.91691, -41.92872, 
        -41.94883, -41.97894, -42.01462, -42.05556, -42.09969, -42.14401, 
        -42.1889, -42.23211, -42.27332, -42.31226, -42.35065, -42.38929, 
        -42.43012, -42.47467, -42.52298, -42.57404, -42.62788, -42.68344, 
        -42.73994, -42.79585, -42.84886, -42.89783, -42.94125, -42.97762, 
        -43.00676, -43.02834, -43.0406, -43.04269, -43.03296, -43.01025, 
        -42.97376, -42.92307, -42.85845, -42.78011, -42.68916, -42.58618, 
        -42.47235, -42.34832, -42.21549, -42.07504, -41.92848, -41.77676, 
        -41.62281, -41.46931, -41.31977, -41.17576, -41.0409, -40.91684, 
        -40.80565,
  -41.26114, -41.30671, -41.35205, -41.39678, -41.44113, -41.48512, 
        -41.52857, -41.57147, -41.614, -41.65635, -41.69925, -41.74297, 
        -41.78788, -41.83392, -41.88054, -41.92611, -41.97231, -42.01751, 
        -42.0619, -42.10583, -42.14888, -42.19184, -42.23462, -42.27711, 
        -42.32022, -42.36447, -42.4102, -42.45734, -42.50512, -42.55318, 
        -42.59996, -42.6468, -42.69175, -42.73384, -42.77203, -42.80647, 
        -42.83722, -42.86479, -42.8895, -42.91187, -42.93095, -42.94798, 
        -42.96273, -42.97579, -42.9875, -42.99789, -43.00623, -43.01429, 
        -43.02065, -43.02523, -43.02761, -43.02786, -43.02663, -43.02365, 
        -43.01979, -43.01493, -43.00895, -43.00247, -42.99512, -42.98713, 
        -42.97789, -42.9674, -42.95563, -42.94402, -42.93202, -42.91964, 
        -42.90715, -42.89487, -42.88314, -42.8721, -42.8616, -42.85149, 
        -42.84185, -42.83269, -42.8247, -42.81804, -42.81336, -42.81164, 
        -42.81295, -42.81767, -42.82415, -42.83443, -42.84688, -42.86053, 
        -42.87486, -42.88974, -42.90467, -42.92025, -42.93673, -42.95359, 
        -42.97113, -42.98785, -43.00269, -43.01512, -43.02486, -43.03234, 
        -43.0386, -43.04408, -43.04865, -43.05378, -43.05853, -43.06278, 
        -43.0661, -43.06775, -43.06889, -43.06981, -43.07106, -43.07453, 
        -43.08236, -43.09603, -43.11717, -43.14653, -43.18386, -43.22786, 
        -43.27662, -43.32754, -43.37785, -43.42481, -43.46923, -43.50951, 
        -43.54569, -43.57807, -43.60726, -43.63386, -43.65891, -43.6825, 
        -43.70427, -43.72406, -43.7415, -43.75638, -43.76855, -43.77888, 
        -43.78778, -43.79601, -43.80399, -43.81172, -43.81906, -43.82576, 
        -43.8305, -43.83481, -43.83706, -43.83688, -43.83442, -43.8297, 
        -43.82342, -43.81542, -43.8067, -43.79781, -43.78916, -43.78075, 
        -43.77241, -43.76377, -43.75489, -43.74594, -43.73691, -43.72725, 
        -43.71699, -43.70584, -43.69373, -43.68076, -43.66654, -43.65346, 
        -43.64092, -43.629, -43.61783, -43.60737, -43.59725, -43.5877, 
        -43.57796, -43.56744, -43.55548, -43.54196, -43.52745, -43.51284, 
        -43.49881, -43.48576, -43.47406, -43.46366, -43.45424, -43.44519, 
        -43.43559, -43.42486, -43.41289, -43.39944, -43.38343, -43.36626, 
        -43.34678, -43.32533, -43.30233, -43.27844, -43.25299, -43.22672, 
        -43.19905, -43.16985, -43.13998, -43.10989, -43.08119, -43.0551, 
        -43.03255, -43.01416, -42.99997, -42.9896, -42.98215, -42.97629, 
        -42.97052, -42.96372, -42.95508, -42.9446, -42.93245, -42.91959, 
        -42.90601, -42.89287, -42.87912, -42.86757, -42.85818, -42.85061, 
        -42.84636, -42.8451, -42.84635, -42.84921, -42.85229, -42.85498, 
        -42.85448, -42.8505, -42.84179, -42.82791, -42.80899, -42.78551, 
        -42.75906, -42.73076, -42.70279, -42.67617, -42.65131, -42.62753, 
        -42.60331, -42.57688, -42.54635, -42.51031, -42.46811, -42.42022, 
        -42.36801, -42.31372, -42.25983, -42.20905, -42.16221, -42.12307, 
        -42.09196, -42.06939, -42.05464, -42.0481, -42.05011, -42.06079, 
        -42.07989, -42.10689, -42.13995, -42.17802, -42.21927, -42.26176, 
        -42.3044, -42.34542, -42.38446, -42.42197, -42.45784, -42.49387, 
        -42.53226, -42.57314, -42.61684, -42.66349, -42.71196, -42.76213, 
        -42.81267, -42.86285, -42.91003, -42.95361, -42.99137, -43.02315, 
        -43.04845, -43.06661, -43.07598, -43.07553, -43.06379, -43.03946, 
        -43.00182, -42.95037, -42.88527, -42.80618, -42.7158, -42.61383, 
        -42.5016, -42.37994, -42.24986, -42.11236, -41.9689, -41.82063, 
        -41.66907, -41.51667, -41.36602, -41.21945, -41.07965, -40.94921, 
        -40.82994,
  -41.26333, -41.31146, -41.35864, -41.4052, -41.45085, -41.49583, 
        -41.53993, -41.58345, -41.62638, -41.66897, -41.71181, -41.75421, 
        -41.79843, -41.84346, -41.88927, -41.93497, -41.98001, -42.02447, 
        -42.0676, -42.11067, -42.15292, -42.1948, -42.23616, -42.27746, 
        -42.31922, -42.36076, -42.40434, -42.44872, -42.49355, -42.53862, 
        -42.58343, -42.62743, -42.66937, -42.7085, -42.74422, -42.77628, 
        -42.80479, -42.83005, -42.85221, -42.87125, -42.88791, -42.90104, 
        -42.91374, -42.92467, -42.93465, -42.94349, -42.95173, -42.95889, 
        -42.96465, -42.96856, -42.97018, -42.96958, -42.96714, -42.96281, 
        -42.95732, -42.95117, -42.94424, -42.93578, -42.92792, -42.9195, 
        -42.91006, -42.8997, -42.88932, -42.87879, -42.86808, -42.85715, 
        -42.8467, -42.83667, -42.82754, -42.81876, -42.81063, -42.80323, 
        -42.79649, -42.79005, -42.78343, -42.77929, -42.77684, -42.77703, 
        -42.78038, -42.78672, -42.79632, -42.80844, -42.82248, -42.83754, 
        -42.85329, -42.86938, -42.88612, -42.90304, -42.9203, -42.93816, 
        -42.95612, -42.97178, -42.98691, -43.00012, -43.01102, -43.02037, 
        -43.02912, -43.03762, -43.04637, -43.05537, -43.06438, -43.07314, 
        -43.08154, -43.08921, -43.09617, -43.10316, -43.11013, -43.11828, 
        -43.1296, -43.14505, -43.16477, -43.1925, -43.22715, -43.26766, 
        -43.31226, -43.35896, -43.40555, -43.45048, -43.49275, -43.53139, 
        -43.56675, -43.59901, -43.62857, -43.65594, -43.68155, -43.70525, 
        -43.72726, -43.74732, -43.76513, -43.78045, -43.79241, -43.80339, 
        -43.81324, -43.82243, -43.83123, -43.83963, -43.84754, -43.85486, 
        -43.86117, -43.866, -43.86858, -43.86851, -43.86602, -43.86119, 
        -43.85438, -43.84641, -43.83765, -43.82934, -43.82176, -43.81499, 
        -43.80887, -43.80279, -43.79575, -43.78956, -43.78308, -43.77575, 
        -43.76762, -43.75837, -43.7481, -43.73707, -43.72583, -43.71474, 
        -43.70425, -43.69457, -43.68568, -43.67753, -43.67015, -43.66291, 
        -43.65559, -43.64718, -43.6373, -43.62585, -43.61376, -43.60154, 
        -43.58982, -43.57861, -43.56734, -43.55789, -43.5487, -43.53923, 
        -43.52928, -43.51805, -43.5056, -43.49156, -43.47634, -43.45921, 
        -43.44012, -43.41996, -43.39889, -43.37716, -43.35452, -43.3303, 
        -43.30449, -43.2766, -43.24731, -43.21743, -43.18804, -43.16044, 
        -43.13537, -43.11354, -43.0951, -43.07986, -43.06611, -43.0552, 
        -43.04506, -43.03447, -43.02326, -43.01093, -42.99786, -42.98436, 
        -42.97068, -42.95749, -42.9453, -42.93451, -42.92572, -42.91867, 
        -42.91385, -42.91164, -42.91141, -42.91219, -42.91361, -42.91478, 
        -42.91341, -42.90764, -42.8975, -42.88214, -42.86232, -42.83805, 
        -42.81091, -42.78278, -42.755, -42.72858, -42.70417, -42.68026, 
        -42.6574, -42.63293, -42.60502, -42.57225, -42.53426, -42.49147, 
        -42.44519, -42.39795, -42.35148, -42.30831, -42.2702, -42.23849, 
        -42.21383, -42.1962, -42.18535, -42.18092, -42.18373, -42.19382, 
        -42.21096, -42.2346, -42.26439, -42.29916, -42.33752, -42.37701, 
        -42.41657, -42.45503, -42.49168, -42.52649, -42.55996, -42.5935, 
        -42.62821, -42.66494, -42.70397, -42.74543, -42.78904, -42.83375, 
        -42.87787, -42.92184, -42.96367, -43.00171, -43.03458, -43.06204, 
        -43.08364, -43.09848, -43.10492, -43.10234, -43.089, -43.0636, 
        -43.0252, -42.97313, -42.90749, -42.82882, -42.7379, -42.63556, 
        -42.52292, -42.40176, -42.27274, -42.13765, -41.99752, -41.85316, 
        -41.70588, -41.55708, -41.40878, -41.26298, -41.12212, -40.98873, 
        -40.86435,
  -41.26429, -41.31324, -41.36179, -41.4099, -41.45687, -41.50283, 
        -41.54692, -41.59124, -41.63453, -41.67708, -41.71985, -41.76305, 
        -41.80644, -41.85059, -41.8952, -41.93959, -41.98347, -42.02661, 
        -42.06877, -42.11124, -42.151, -42.19247, -42.23275, -42.27353, 
        -42.31403, -42.35509, -42.39653, -42.43836, -42.48051, -42.52254, 
        -42.56418, -42.60501, -42.64414, -42.68073, -42.71386, -42.74365, 
        -42.7689, -42.79179, -42.81121, -42.82751, -42.84153, -42.85307, 
        -42.86306, -42.87188, -42.88047, -42.88806, -42.89524, -42.90182, 
        -42.90728, -42.91059, -42.91183, -42.90964, -42.90627, -42.90092, 
        -42.89405, -42.88676, -42.87891, -42.87056, -42.86169, -42.85276, 
        -42.84283, -42.83321, -42.8236, -42.81409, -42.80487, -42.79648, 
        -42.78854, -42.78119, -42.77338, -42.76764, -42.7622, -42.75772, 
        -42.75358, -42.74977, -42.74656, -42.74464, -42.74413, -42.74611, 
        -42.75077, -42.75892, -42.7701, -42.78339, -42.79863, -42.81497, 
        -42.83194, -42.84828, -42.86608, -42.88448, -42.90276, -42.9217, 
        -42.93941, -42.95666, -42.97198, -42.98563, -42.99775, -43.00897, 
        -43.01972, -43.03086, -43.0425, -43.05463, -43.06727, -43.08023, 
        -43.09318, -43.10587, -43.1171, -43.12891, -43.1408, -43.15322, 
        -43.16774, -43.18465, -43.20554, -43.23169, -43.26389, -43.30107, 
        -43.34188, -43.38469, -43.42802, -43.47012, -43.50995, -43.54726, 
        -43.58178, -43.61362, -43.64315, -43.66962, -43.69542, -43.71937, 
        -43.74164, -43.76181, -43.77979, -43.79553, -43.80915, -43.82097, 
        -43.83163, -43.84162, -43.85124, -43.86034, -43.86886, -43.87674, 
        -43.88353, -43.88868, -43.89151, -43.89171, -43.88936, -43.88475, 
        -43.87836, -43.8697, -43.86153, -43.85406, -43.84777, -43.84296, 
        -43.839, -43.83524, -43.83184, -43.82826, -43.82412, -43.81905, 
        -43.81265, -43.80507, -43.79649, -43.78699, -43.77766, -43.76836, 
        -43.75972, -43.75168, -43.74538, -43.73933, -43.73414, -43.72893, 
        -43.72268, -43.71609, -43.7081, -43.69864, -43.68864, -43.67873, 
        -43.66922, -43.66001, -43.65129, -43.64278, -43.63426, -43.62527, 
        -43.61485, -43.60312, -43.59035, -43.57621, -43.56111, -43.54433, 
        -43.52553, -43.5064, -43.48684, -43.4668, -43.44611, -43.42393, 
        -43.39927, -43.37169, -43.34313, -43.31382, -43.28442, -43.25606, 
        -43.2298, -43.20601, -43.18509, -43.16673, -43.15062, -43.13605, 
        -43.12238, -43.10901, -43.09525, -43.08142, -43.06738, -43.05346, 
        -43.03981, -43.02728, -43.01589, -43.00605, -42.99771, -42.99081, 
        -42.98561, -42.98229, -42.98016, -42.97906, -42.9784, -42.97755, 
        -42.97308, -42.96593, -42.95426, -42.93755, -42.917, -42.8927, 
        -42.86578, -42.8381, -42.81123, -42.78571, -42.76207, -42.74, 
        -42.71855, -42.69556, -42.66985, -42.63995, -42.60555, -42.56733, 
        -42.52693, -42.48585, -42.446, -42.40937, -42.37806, -42.35253, 
        -42.33321, -42.31994, -42.31213, -42.30976, -42.31336, -42.32291, 
        -42.33813, -42.35901, -42.38544, -42.41634, -42.44977, -42.4857, 
        -42.52137, -42.55679, -42.59048, -42.62254, -42.65311, -42.68385, 
        -42.71505, -42.74761, -42.78215, -42.8187, -42.85717, -42.89671, 
        -42.93661, -42.97519, -43.01155, -43.0443, -43.07261, -43.09608, 
        -43.11423, -43.12613, -43.12999, -43.12542, -43.11079, -43.08422, 
        -43.0449, -42.99202, -42.92577, -42.84658, -42.75444, -42.65021, 
        -42.53624, -42.41396, -42.28505, -42.15121, -42.01419, -41.87431, 
        -41.73221, -41.58884, -41.44553, -41.30398, -41.16549, -41.03266, 
        -40.90658,
  -41.26267, -41.31142, -41.36069, -41.40965, -41.45741, -41.50453, 
        -41.55047, -41.59535, -41.6391, -41.68209, -41.72478, -41.76775, 
        -41.81086, -41.85428, -41.89766, -41.93985, -41.98249, -42.02419, 
        -42.06546, -42.10681, -42.14725, -42.18756, -42.2276, -42.26736, 
        -42.30696, -42.34676, -42.38671, -42.4263, -42.4658, -42.50494, 
        -42.54255, -42.58009, -42.61613, -42.6498, -42.68061, -42.70813, 
        -42.73231, -42.75287, -42.76984, -42.78352, -42.79456, -42.80345, 
        -42.81072, -42.81774, -42.82507, -42.8319, -42.83734, -42.84313, 
        -42.84806, -42.85129, -42.85221, -42.85071, -42.84685, -42.84106, 
        -42.8336, -42.82492, -42.81587, -42.80634, -42.79647, -42.78678, 
        -42.77726, -42.76812, -42.75859, -42.75079, -42.74382, -42.73817, 
        -42.73285, -42.72842, -42.72489, -42.72208, -42.71965, -42.71758, 
        -42.71601, -42.71495, -42.71406, -42.71375, -42.71489, -42.71815, 
        -42.72424, -42.73242, -42.7446, -42.75917, -42.77524, -42.79232, 
        -42.81013, -42.82847, -42.8474, -42.86663, -42.88617, -42.90514, 
        -42.92352, -42.94088, -42.95648, -42.97062, -42.98402, -42.99674, 
        -43.00972, -43.02306, -43.03592, -43.05084, -43.06657, -43.08303, 
        -43.09974, -43.11645, -43.13278, -43.14918, -43.16535, -43.18178, 
        -43.19881, -43.21759, -43.23898, -43.26408, -43.29394, -43.3282, 
        -43.36602, -43.40555, -43.44543, -43.48405, -43.52192, -43.55778, 
        -43.59117, -43.62215, -43.65091, -43.67815, -43.70376, -43.72771, 
        -43.74965, -43.76979, -43.78793, -43.8041, -43.81821, -43.83075, 
        -43.84219, -43.85297, -43.8632, -43.87307, -43.88243, -43.88999, 
        -43.89733, -43.90288, -43.90609, -43.90673, -43.90498, -43.90103, 
        -43.89547, -43.88873, -43.88178, -43.87553, -43.87072, -43.86748, 
        -43.86551, -43.86409, -43.86298, -43.86153, -43.85937, -43.85597, 
        -43.85102, -43.84492, -43.83763, -43.82984, -43.82082, -43.8129, 
        -43.80593, -43.80002, -43.79549, -43.79137, -43.78778, -43.78441, 
        -43.78091, -43.7763, -43.77, -43.76244, -43.75437, -43.74671, 
        -43.73933, -43.73225, -43.72532, -43.71798, -43.70983, -43.70107, 
        -43.69072, -43.67901, -43.66637, -43.65239, -43.63662, -43.6199, 
        -43.60238, -43.58385, -43.56548, -43.54694, -43.52747, -43.50628, 
        -43.48278, -43.45702, -43.42945, -43.40084, -43.37189, -43.34363, 
        -43.31719, -43.29297, -43.27111, -43.25147, -43.23338, -43.21655, 
        -43.20036, -43.18449, -43.16882, -43.15361, -43.13868, -43.12453, 
        -43.11115, -43.09912, -43.08738, -43.07799, -43.07012, -43.06334, 
        -43.05735, -43.05265, -43.04873, -43.0456, -43.04296, -43.03948, 
        -43.03376, -43.02473, -43.01165, -42.99451, -42.97367, -42.94998, 
        -42.92427, -42.89814, -42.87274, -42.84868, -42.82613, -42.80501, 
        -42.78425, -42.76262, -42.73844, -42.71099, -42.67982, -42.64552, 
        -42.60976, -42.57396, -42.5397, -42.50907, -42.48229, -42.46188, 
        -42.44681, -42.43679, -42.43137, -42.43063, -42.43457, -42.44333, 
        -42.45673, -42.47491, -42.49768, -42.52467, -42.55481, -42.58657, 
        -42.61879, -42.65048, -42.68101, -42.71016, -42.73806, -42.76588, 
        -42.79385, -42.82258, -42.85298, -42.88482, -42.91843, -42.95306, 
        -42.98767, -43.02133, -43.05248, -43.08068, -43.10516, -43.1252, 
        -43.14021, -43.14916, -43.15093, -43.14485, -43.12882, -43.10107, 
        -43.06116, -43.00766, -42.93955, -42.8587, -42.76487, -42.65846, 
        -42.54163, -42.41698, -42.28667, -42.15324, -42.01845, -41.88252, 
        -41.74637, -41.61001, -41.47387, -41.33912, -41.20648, -41.07729, 
        -40.95262,
  -41.25756, -41.30757, -41.35702, -41.40618, -41.45448, -41.5021, 
        -41.54866, -41.59391, -41.63817, -41.68151, -41.72356, -41.7666, 
        -41.80957, -41.85238, -41.89465, -41.93651, -41.97781, -42.01873, 
        -42.05921, -42.09948, -42.13979, -42.17968, -42.21924, -42.2586, 
        -42.29776, -42.33576, -42.37439, -42.41225, -42.44928, -42.48558, 
        -42.52119, -42.55566, -42.58875, -42.61983, -42.64818, -42.67322, 
        -42.69495, -42.71289, -42.72706, -42.73766, -42.74565, -42.75082, 
        -42.75618, -42.76148, -42.76693, -42.77268, -42.77867, -42.78449, 
        -42.78936, -42.79248, -42.79346, -42.79176, -42.78792, -42.78175, 
        -42.7738, -42.76424, -42.75412, -42.74265, -42.73243, -42.72275, 
        -42.71376, -42.70568, -42.69883, -42.69296, -42.68826, -42.68509, 
        -42.68272, -42.6814, -42.68094, -42.681, -42.68146, -42.68224, 
        -42.68333, -42.68435, -42.68466, -42.68614, -42.68871, -42.69315, 
        -42.70018, -42.7104, -42.72332, -42.73847, -42.7548, -42.77224, 
        -42.79047, -42.80948, -42.82878, -42.84848, -42.86808, -42.88734, 
        -42.90574, -42.92233, -42.93852, -42.95369, -42.96814, -42.98242, 
        -42.99722, -43.01244, -43.02871, -43.04617, -43.06489, -43.08436, 
        -43.10415, -43.1244, -43.14449, -43.16446, -43.18415, -43.20376, 
        -43.22343, -43.24389, -43.26496, -43.28949, -43.31756, -43.34952, 
        -43.3848, -43.42175, -43.45892, -43.4961, -43.53223, -43.56635, 
        -43.59803, -43.62759, -43.65514, -43.68127, -43.70607, -43.7294, 
        -43.75097, -43.77102, -43.78912, -43.80543, -43.81905, -43.83226, 
        -43.84442, -43.85581, -43.86684, -43.87753, -43.88759, -43.89698, 
        -43.90495, -43.91109, -43.91489, -43.91624, -43.91539, -43.91257, 
        -43.90834, -43.90321, -43.89786, -43.89318, -43.89008, -43.88864, 
        -43.88834, -43.88871, -43.88829, -43.88856, -43.88786, -43.88565, 
        -43.8819, -43.87707, -43.8711, -43.86457, -43.8577, -43.8515, 
        -43.84608, -43.84174, -43.83829, -43.83584, -43.83409, -43.8325, 
        -43.83043, -43.8273, -43.82268, -43.81665, -43.81046, -43.80449, 
        -43.79867, -43.79332, -43.78677, -43.78073, -43.77343, -43.76496, 
        -43.75502, -43.74361, -43.73125, -43.7179, -43.70356, -43.68817, 
        -43.67111, -43.65385, -43.63582, -43.6182, -43.59944, -43.57847, 
        -43.55635, -43.53158, -43.505, -43.47715, -43.44933, -43.42205, 
        -43.39623, -43.3728, -43.35138, -43.33161, -43.31203, -43.29387, 
        -43.27603, -43.25835, -43.2412, -43.22496, -43.20942, -43.19499, 
        -43.18172, -43.17001, -43.15972, -43.15047, -43.14257, -43.13531, 
        -43.12868, -43.1227, -43.11731, -43.11243, -43.10746, -43.10155, 
        -43.09369, -43.08296, -43.06882, -43.0515, -43.03129, -43.00873, 
        -42.98473, -42.96064, -42.9369, -42.91442, -42.89185, -42.87167, 
        -42.85155, -42.83064, -42.80787, -42.7824, -42.75402, -42.72328, 
        -42.69133, -42.65989, -42.63045, -42.60468, -42.58333, -42.56688, 
        -42.55496, -42.54705, -42.5434, -42.54399, -42.54841, -42.55651, 
        -42.56822, -42.5836, -42.60305, -42.62608, -42.65188, -42.67953, 
        -42.70797, -42.73589, -42.76309, -42.78873, -42.8139, -42.83878, 
        -42.86375, -42.88917, -42.91566, -42.94324, -42.97229, -43.00117, 
        -43.03103, -43.05976, -43.08625, -43.11028, -43.13145, -43.14839, 
        -43.16039, -43.16721, -43.16711, -43.15963, -43.14225, -43.1137, 
        -43.07277, -43.01849, -42.95028, -42.86777, -42.77133, -42.66227, 
        -42.54227, -42.41428, -42.28184, -42.14781, -42.01432, -41.88226, 
        -41.75208, -41.62311, -41.49533, -41.36884, -41.24402, -41.12111, 
        -41.00031,
  -41.25076, -41.30003, -41.34922, -41.39812, -41.44642, -41.49426, 
        -41.54018, -41.58601, -41.63067, -41.67471, -41.7183, -41.76147, 
        -41.80444, -41.84679, -41.88837, -41.92924, -41.96949, -42.00949, 
        -42.04932, -42.08928, -42.12845, -42.1684, -42.20803, -42.24727, 
        -42.28605, -42.32439, -42.36173, -42.39801, -42.43299, -42.46692, 
        -42.49975, -42.53153, -42.56175, -42.58998, -42.6158, -42.63743, 
        -42.65646, -42.67148, -42.68273, -42.6902, -42.69502, -42.69847, 
        -42.70153, -42.70488, -42.70908, -42.71407, -42.71981, -42.72565, 
        -42.73069, -42.7341, -42.73547, -42.73298, -42.72894, -42.72243, 
        -42.7141, -42.70416, -42.69323, -42.68258, -42.67245, -42.66317, 
        -42.65519, -42.64868, -42.64389, -42.64034, -42.63802, -42.63709, 
        -42.63763, -42.639, -42.64032, -42.64323, -42.64655, -42.64993, 
        -42.65337, -42.65677, -42.66008, -42.66338, -42.66732, -42.67289, 
        -42.68079, -42.69167, -42.70497, -42.72038, -42.73701, -42.75426, 
        -42.7723, -42.79027, -42.8096, -42.82912, -42.84854, -42.8676, 
        -42.88599, -42.90367, -42.92076, -42.93682, -42.95248, -42.96827, 
        -42.98463, -43.00181, -43.02008, -43.03986, -43.06107, -43.08323, 
        -43.10606, -43.12917, -43.15138, -43.17438, -43.19696, -43.21907, 
        -43.24093, -43.26295, -43.2859, -43.3105, -43.33755, -43.36768, 
        -43.40059, -43.43527, -43.47047, -43.50537, -43.53932, -43.57181, 
        -43.6017, -43.62967, -43.6556, -43.6792, -43.70266, -43.72482, 
        -43.74537, -43.76485, -43.7827, -43.79916, -43.81419, -43.82805, 
        -43.84096, -43.85318, -43.86502, -43.87645, -43.88731, -43.89745, 
        -43.90609, -43.91299, -43.91764, -43.91998, -43.92029, -43.91906, 
        -43.91544, -43.91218, -43.90862, -43.90601, -43.90454, -43.90471, 
        -43.906, -43.90769, -43.90944, -43.91082, -43.91121, -43.91002, 
        -43.90723, -43.90329, -43.89843, -43.89318, -43.88782, -43.88285, 
        -43.87875, -43.87576, -43.87384, -43.87276, -43.87227, -43.87104, 
        -43.87035, -43.86852, -43.86522, -43.86067, -43.85583, -43.85127, 
        -43.84695, -43.8427, -43.83838, -43.83345, -43.82715, -43.81939, 
        -43.80995, -43.79905, -43.78708, -43.77441, -43.7611, -43.74675, 
        -43.73117, -43.71437, -43.69726, -43.67997, -43.66169, -43.64168, 
        -43.61985, -43.59499, -43.56955, -43.54301, -43.51648, -43.49071, 
        -43.46649, -43.44423, -43.42399, -43.40492, -43.38654, -43.36807, 
        -43.34956, -43.33093, -43.31297, -43.29583, -43.27975, -43.26517, 
        -43.25191, -43.2402, -43.22998, -43.22071, -43.21225, -43.20415, 
        -43.19688, -43.18971, -43.1827, -43.17612, -43.16909, -43.16108, 
        -43.15015, -43.1381, -43.12344, -43.10656, -43.08744, -43.06661, 
        -43.04459, -43.0224, -43.00056, -42.97942, -42.95897, -42.93918, 
        -42.91973, -42.89943, -42.87787, -42.85409, -42.82821, -42.80047, 
        -42.77204, -42.74432, -42.71886, -42.69695, -42.679, -42.66515, 
        -42.65546, -42.64947, -42.64713, -42.64833, -42.65276, -42.66018, 
        -42.66994, -42.68282, -42.69915, -42.71856, -42.73955, -42.76352, 
        -42.78793, -42.81226, -42.8356, -42.85856, -42.88081, -42.90264, 
        -42.9245, -42.94666, -42.9696, -42.99334, -43.01829, -43.04395, 
        -43.06923, -43.09343, -43.1159, -43.13638, -43.15403, -43.16801, 
        -43.17768, -43.18229, -43.18081, -43.17175, -43.15317, -43.12364, 
        -43.08176, -43.02644, -42.95689, -42.87278, -42.77401, -42.66168, 
        -42.53793, -42.40641, -42.27134, -42.13582, -42.00291, -41.87383, 
        -41.7487, -41.62688, -41.50764, -41.3902, -41.27413, -41.15885, 
        -41.04387,
  -41.24048, -41.28745, -41.33569, -41.38397, -41.43185, -41.47968, 
        -41.52692, -41.57314, -41.61872, -41.66353, -41.70811, -41.75187, 
        -41.79495, -41.83708, -41.87791, -41.91683, -41.95628, -41.99585, 
        -42.03557, -42.07564, -42.11606, -42.15629, -42.19616, -42.23526, 
        -42.27375, -42.31113, -42.34744, -42.38235, -42.41578, -42.44781, 
        -42.47738, -42.50646, -42.53402, -42.55956, -42.5827, -42.60261, 
        -42.61874, -42.63075, -42.63877, -42.64327, -42.64493, -42.64566, 
        -42.64649, -42.6484, -42.65157, -42.65612, -42.6606, -42.66651, 
        -42.67176, -42.67576, -42.67713, -42.67601, -42.67197, -42.66547, 
        -42.65701, -42.64715, -42.63626, -42.62577, -42.61638, -42.60822, 
        -42.60195, -42.59724, -42.59354, -42.59224, -42.59221, -42.59319, 
        -42.59582, -42.59973, -42.60454, -42.61029, -42.61627, -42.6223, 
        -42.62804, -42.63352, -42.63875, -42.64394, -42.64939, -42.65626, 
        -42.66483, -42.67523, -42.68887, -42.70418, -42.72042, -42.73727, 
        -42.75474, -42.77282, -42.79162, -42.81063, -42.82966, -42.84829, 
        -42.86653, -42.88452, -42.90221, -42.91954, -42.9365, -42.95364, 
        -42.97144, -42.98936, -43.00937, -43.03102, -43.05443, -43.07916, 
        -43.1045, -43.13031, -43.15591, -43.18142, -43.20614, -43.23022, 
        -43.25391, -43.2774, -43.30122, -43.32616, -43.35272, -43.38144, 
        -43.41236, -43.44497, -43.4782, -43.51009, -43.54196, -43.5722, 
        -43.60028, -43.62635, -43.65024, -43.67303, -43.69483, -43.7154, 
        -43.73496, -43.7534, -43.77089, -43.78756, -43.80298, -43.81738, 
        -43.83102, -43.84406, -43.85669, -43.86893, -43.88058, -43.89048, 
        -43.9, -43.90773, -43.91333, -43.91681, -43.91853, -43.91875, 
        -43.91808, -43.91679, -43.91549, -43.91492, -43.91525, -43.91685, 
        -43.91923, -43.92204, -43.92468, -43.92684, -43.92782, -43.92733, 
        -43.9254, -43.92255, -43.91883, -43.9137, -43.90952, -43.90576, 
        -43.9029, -43.90125, -43.90069, -43.90096, -43.90166, -43.90261, 
        -43.90275, -43.90237, -43.90052, -43.89705, -43.89333, -43.8897, 
        -43.88639, -43.88317, -43.87984, -43.8758, -43.87037, -43.86355, 
        -43.85482, -43.84439, -43.83311, -43.82116, -43.80802, -43.79519, 
        -43.7811, -43.76585, -43.7497, -43.73274, -43.71468, -43.69512, 
        -43.67376, -43.65067, -43.62637, -43.60134, -43.57634, -43.5522, 
        -43.52983, -43.50931, -43.49044, -43.4725, -43.45471, -43.43673, 
        -43.41798, -43.39924, -43.38073, -43.36303, -43.34676, -43.33203, 
        -43.31874, -43.30573, -43.29489, -43.28497, -43.27596, -43.26716, 
        -43.25859, -43.25044, -43.2425, -43.23457, -43.22589, -43.2159, 
        -43.20448, -43.19118, -43.17651, -43.16042, -43.14268, -43.1236, 
        -43.10389, -43.08379, -43.06368, -43.04371, -43.02402, -43.00486, 
        -42.98567, -42.9662, -42.9457, -42.92355, -42.89964, -42.87462, 
        -42.84916, -42.82473, -42.80285, -42.78399, -42.76787, -42.75627, 
        -42.74803, -42.74311, -42.74169, -42.74315, -42.74725, -42.7535, 
        -42.76178, -42.77224, -42.78548, -42.80133, -42.81968, -42.83985, 
        -42.86076, -42.88158, -42.90163, -42.92125, -42.94037, -42.95941, 
        -42.97863, -42.99789, -43.01769, -43.03802, -43.05924, -43.08072, 
        -43.1022, -43.12259, -43.14167, -43.15887, -43.17348, -43.18472, 
        -43.19187, -43.19438, -43.19093, -43.18025, -43.16039, -43.12951, 
        -43.08667, -43.03046, -42.95858, -42.87275, -42.77187, -42.65672, 
        -42.52961, -42.39455, -42.25613, -42.11852, -41.98512, -41.8577, 
        -41.73656, -41.62083, -41.50917, -41.40035, -41.29305, -41.18599, 
        -41.078,
  -41.22461, -41.2711, -41.31821, -41.36563, -41.4132, -41.46079, 
        -41.50833, -41.5553, -41.60163, -41.64741, -41.69163, -41.73629, 
        -41.7796, -41.82161, -41.86214, -41.9017, -41.94072, -41.97992, 
        -42.01981, -42.06024, -42.10101, -42.14141, -42.18135, -42.22068, 
        -42.25901, -42.29501, -42.33048, -42.36418, -42.39617, -42.42659, 
        -42.45513, -42.48191, -42.507, -42.53009, -42.55051, -42.56789, 
        -42.5812, -42.59019, -42.59538, -42.5969, -42.59581, -42.59303, 
        -42.59184, -42.59212, -42.59445, -42.59864, -42.60399, -42.60983, 
        -42.61549, -42.61945, -42.62116, -42.62038, -42.61676, -42.61043, 
        -42.60218, -42.59264, -42.58249, -42.57155, -42.56322, -42.55681, 
        -42.55256, -42.5501, -42.54923, -42.55015, -42.55198, -42.55495, 
        -42.5594, -42.56513, -42.5722, -42.58028, -42.58877, -42.59705, 
        -42.60498, -42.61122, -42.61835, -42.62515, -42.63225, -42.64013, 
        -42.64974, -42.66174, -42.67555, -42.69069, -42.70654, -42.72277, 
        -42.7392, -42.7562, -42.77385, -42.79196, -42.81064, -42.82888, 
        -42.84698, -42.86425, -42.88239, -42.90076, -42.91903, -42.93731, 
        -42.95655, -42.97682, -42.9987, -43.02184, -43.04702, -43.07354, 
        -43.10112, -43.12896, -43.15668, -43.18405, -43.21048, -43.23624, 
        -43.26139, -43.2861, -43.30984, -43.33504, -43.36136, -43.38906, 
        -43.41837, -43.44883, -43.48005, -43.51118, -43.54095, -43.56907, 
        -43.59516, -43.6191, -43.64137, -43.66222, -43.68197, -43.70091, 
        -43.71908, -43.7365, -43.75352, -43.76996, -43.78468, -43.79973, 
        -43.81406, -43.82788, -43.84133, -43.85432, -43.86664, -43.87817, 
        -43.88834, -43.89681, -43.90339, -43.90814, -43.91141, -43.9135, 
        -43.91489, -43.91563, -43.9165, -43.91777, -43.91988, -43.92273, 
        -43.92603, -43.92949, -43.93182, -43.93443, -43.93612, -43.93634, 
        -43.93525, -43.93327, -43.93088, -43.92789, -43.92478, -43.92212, 
        -43.92085, -43.92043, -43.9211, -43.9225, -43.92401, -43.9257, 
        -43.92687, -43.92753, -43.92656, -43.92403, -43.92133, -43.91842, 
        -43.91594, -43.91278, -43.91018, -43.907, -43.90255, -43.89669, 
        -43.88876, -43.87913, -43.86861, -43.85765, -43.84658, -43.83507, 
        -43.8225, -43.80855, -43.79348, -43.77726, -43.75963, -43.74065, 
        -43.71993, -43.6979, -43.67493, -43.65128, -43.62797, -43.60569, 
        -43.58507, -43.56616, -43.54869, -43.53164, -43.51387, -43.49632, 
        -43.47816, -43.4596, -43.44107, -43.42339, -43.40718, -43.39262, 
        -43.37942, -43.3673, -43.35588, -43.34522, -43.33508, -43.32527, 
        -43.31551, -43.30614, -43.29706, -43.28778, -43.27776, -43.26643, 
        -43.25408, -43.24026, -43.22575, -43.21057, -43.19423, -43.17703, 
        -43.15902, -43.14051, -43.1218, -43.10281, -43.0829, -43.06431, 
        -43.04592, -43.02758, -43.0084, -42.98821, -42.96653, -42.94379, 
        -42.92118, -42.89981, -42.88072, -42.86451, -42.85123, -42.84115, 
        -42.83401, -42.83012, -42.82895, -42.83031, -42.83392, -42.83892, 
        -42.84565, -42.85395, -42.86437, -42.87724, -42.89222, -42.90874, 
        -42.92634, -42.94369, -42.9607, -42.97734, -42.99348, -43.0097, 
        -43.02615, -43.04244, -43.05919, -43.07671, -43.0943, -43.11113, 
        -43.12908, -43.14633, -43.16244, -43.17675, -43.18834, -43.19687, 
        -43.20151, -43.20167, -43.19603, -43.18342, -43.16196, -43.12996, 
        -43.08611, -43.02912, -42.95751, -42.87032, -42.76778, -42.65025, 
        -42.52048, -42.38223, -42.24044, -42.10007, -41.96514, -41.83787, 
        -41.71912, -41.60768, -41.50222, -41.40067, -41.30129, -41.20221, 
        -41.10152,
  -41.20354, -41.24892, -41.29508, -41.34184, -41.3892, -41.43586, 
        -41.48363, -41.5313, -41.57838, -41.62498, -41.6711, -41.71632, 
        -41.76011, -41.80234, -41.84277, -41.88232, -41.92122, -41.96069, 
        -42.00069, -42.04131, -42.08134, -42.12206, -42.16234, -42.20192, 
        -42.24016, -42.2768, -42.31153, -42.34423, -42.37506, -42.40382, 
        -42.43071, -42.45546, -42.4782, -42.49904, -42.51702, -42.53079, 
        -42.54156, -42.54813, -42.55059, -42.54985, -42.54665, -42.54288, 
        -42.53995, -42.5392, -42.54054, -42.54426, -42.54932, -42.55505, 
        -42.56048, -42.56473, -42.56683, -42.56546, -42.56237, -42.5565, 
        -42.54871, -42.5398, -42.5308, -42.52239, -42.51538, -42.51079, 
        -42.5082, -42.50786, -42.50885, -42.51163, -42.51544, -42.52023, 
        -42.52641, -42.534, -42.54214, -42.5519, -42.56194, -42.57224, 
        -42.58179, -42.59075, -42.59935, -42.60769, -42.61609, -42.6254, 
        -42.63602, -42.64815, -42.66214, -42.67725, -42.69286, -42.70838, 
        -42.72385, -42.73831, -42.75491, -42.7723, -42.78977, -42.80788, 
        -42.82591, -42.84438, -42.86292, -42.88214, -42.90166, -42.92118, 
        -42.94131, -42.96293, -42.98605, -43.0108, -43.03709, -43.06532, 
        -43.09451, -43.12406, -43.15239, -43.18115, -43.20903, -43.236, 
        -43.26228, -43.28801, -43.31327, -43.33853, -43.3644, -43.39117, 
        -43.41885, -43.44726, -43.47652, -43.5056, -43.53362, -43.5597, 
        -43.58395, -43.60635, -43.62685, -43.645, -43.66305, -43.68011, 
        -43.69672, -43.71307, -43.72934, -43.74549, -43.76133, -43.77659, 
        -43.79144, -43.80607, -43.82004, -43.83353, -43.84657, -43.85863, 
        -43.86928, -43.87833, -43.88581, -43.89199, -43.89698, -43.90102, 
        -43.90339, -43.90636, -43.90932, -43.91246, -43.91599, -43.91982, 
        -43.92386, -43.92789, -43.93188, -43.93512, -43.93721, -43.93838, 
        -43.93831, -43.93748, -43.93593, -43.93424, -43.93261, -43.93117, 
        -43.93094, -43.9314, -43.93303, -43.93547, -43.938, -43.93925, 
        -43.94121, -43.94224, -43.94186, -43.9404, -43.93859, -43.93654, 
        -43.93501, -43.93375, -43.93205, -43.92968, -43.92604, -43.92074, 
        -43.91352, -43.90516, -43.89576, -43.88578, -43.87603, -43.8656, 
        -43.85443, -43.84179, -43.82784, -43.81242, -43.79552, -43.77711, 
        -43.75683, -43.73571, -43.71396, -43.69187, -43.67016, -43.6495, 
        -43.63043, -43.61282, -43.59631, -43.58026, -43.56421, -43.54741, 
        -43.52994, -43.51184, -43.49386, -43.47671, -43.46098, -43.44666, 
        -43.43368, -43.42151, -43.41001, -43.39859, -43.38747, -43.37637, 
        -43.36557, -43.35499, -43.34461, -43.33424, -43.32314, -43.31002, 
        -43.29686, -43.28297, -43.26885, -43.25444, -43.23924, -43.22335, 
        -43.20668, -43.18946, -43.17151, -43.15346, -43.13525, -43.11786, 
        -43.10072, -43.08377, -43.06652, -43.04843, -43.0289, -43.00856, 
        -42.98856, -42.97018, -42.95332, -42.93926, -42.92748, -42.91862, 
        -42.91259, -42.90929, -42.90826, -42.90949, -42.91206, -42.91607, 
        -42.92123, -42.92757, -42.93567, -42.9454, -42.95623, -42.96963, 
        -42.98384, -42.99816, -43.01233, -43.02592, -43.03928, -43.05275, 
        -43.06631, -43.08002, -43.094, -43.10828, -43.12276, -43.13736, 
        -43.15217, -43.1668, -43.18035, -43.19198, -43.20112, -43.20697, 
        -43.20889, -43.20617, -43.19787, -43.18302, -43.16005, -43.12697, 
        -43.08237, -43.02491, -42.95284, -42.86526, -42.76188, -42.64303, 
        -42.51112, -42.37004, -42.22501, -42.08147, -41.944, -41.81552, 
        -41.69715, -41.58817, -41.48664, -41.3905, -41.29772, -41.20579, 
        -41.11137,
  -41.1768, -41.22024, -41.26585, -41.31238, -41.35944, -41.40708, 
        -41.45513, -41.50304, -41.55071, -41.59803, -41.64476, -41.69039, 
        -41.73475, -41.77724, -41.81808, -41.85685, -41.89625, -41.93584, 
        -41.97615, -42.01697, -42.0579, -42.09903, -42.13948, -42.17927, 
        -42.21758, -42.25397, -42.28809, -42.32003, -42.34966, -42.3771, 
        -42.40137, -42.42435, -42.44516, -42.46377, -42.47964, -42.49228, 
        -42.50076, -42.50506, -42.50566, -42.50332, -42.49888, -42.49387, 
        -42.48975, -42.48779, -42.48857, -42.49168, -42.49556, -42.50098, 
        -42.5064, -42.5107, -42.51305, -42.5132, -42.51041, -42.50523, 
        -42.49858, -42.49089, -42.48321, -42.47671, -42.47145, -42.46867, 
        -42.46812, -42.46929, -42.47113, -42.47516, -42.48055, -42.48701, 
        -42.49474, -42.50384, -42.5143, -42.52546, -42.53696, -42.5483, 
        -42.55892, -42.56908, -42.57901, -42.58878, -42.59868, -42.60913, 
        -42.62069, -42.63238, -42.64629, -42.66124, -42.67666, -42.69157, 
        -42.70615, -42.72078, -42.7361, -42.75217, -42.76912, -42.78671, 
        -42.80428, -42.82274, -42.84235, -42.86208, -42.88235, -42.90342, 
        -42.92469, -42.9461, -42.97004, -42.99583, -43.02335, -43.05248, 
        -43.08288, -43.11376, -43.14439, -43.1745, -43.20347, -43.23145, 
        -43.25827, -43.28437, -43.30978, -43.33488, -43.36012, -43.38577, 
        -43.41193, -43.43848, -43.46434, -43.49149, -43.51759, -43.54205, 
        -43.56464, -43.58545, -43.60465, -43.62224, -43.63867, -43.65422, 
        -43.66935, -43.6846, -43.70011, -43.71585, -43.73155, -43.74713, 
        -43.76228, -43.77707, -43.79149, -43.80563, -43.8188, -43.83001, 
        -43.84101, -43.85065, -43.8591, -43.86656, -43.87313, -43.87919, 
        -43.88464, -43.88977, -43.89485, -43.89966, -43.90459, -43.90934, 
        -43.91394, -43.9186, -43.92318, -43.92716, -43.93022, -43.93269, 
        -43.9338, -43.93419, -43.93394, -43.93254, -43.93184, -43.93158, 
        -43.93237, -43.93392, -43.93663, -43.93905, -43.94217, -43.9451, 
        -43.94736, -43.94867, -43.94898, -43.94831, -43.94709, -43.94618, 
        -43.94566, -43.94524, -43.94438, -43.9426, -43.93947, -43.93469, 
        -43.92847, -43.92081, -43.91258, -43.9036, -43.89379, -43.88445, 
        -43.8745, -43.86322, -43.85034, -43.83595, -43.82037, -43.80314, 
        -43.78482, -43.76514, -43.74418, -43.72384, -43.7038, -43.68478, 
        -43.66703, -43.65032, -43.63449, -43.61906, -43.6035, -43.58747, 
        -43.57063, -43.55328, -43.5362, -43.51993, -43.50492, -43.49126, 
        -43.47874, -43.46609, -43.45446, -43.44267, -43.43066, -43.41862, 
        -43.40649, -43.39473, -43.38321, -43.37188, -43.35995, -43.34714, 
        -43.33372, -43.32019, -43.30638, -43.29239, -43.27802, -43.26277, 
        -43.24701, -43.23047, -43.21308, -43.19581, -43.17907, -43.16267, 
        -43.14717, -43.13226, -43.11729, -43.10147, -43.0847, -43.06685, 
        -43.04953, -43.03331, -43.01871, -43.00519, -42.99483, -42.98698, 
        -42.98188, -42.97915, -42.97824, -42.97899, -42.9808, -42.98382, 
        -42.9877, -42.99209, -42.99788, -43.00519, -43.01402, -43.02438, 
        -43.03551, -43.0471, -43.05861, -43.06947, -43.0802, -43.09102, 
        -43.10182, -43.11304, -43.12452, -43.1357, -43.14713, -43.15895, 
        -43.17114, -43.18309, -43.19418, -43.20366, -43.21058, -43.21395, 
        -43.21303, -43.20727, -43.19638, -43.17903, -43.15382, -43.11959, 
        -43.07438, -43.0158, -42.94396, -42.85674, -42.75327, -42.63416, 
        -42.5014, -42.35839, -42.21051, -42.06374, -41.92278, -41.79181, 
        -41.67209, -41.56326, -41.46352, -41.37084, -41.28255, -41.19622, 
        -41.10942,
  -41.14253, -41.18671, -41.23222, -41.2789, -41.32616, -41.37369, 
        -41.42167, -41.46957, -41.51749, -41.56506, -41.61119, -41.65719, 
        -41.70195, -41.74517, -41.78678, -41.82705, -41.86685, -41.90676, 
        -41.94704, -41.98794, -42.02893, -42.07001, -42.11058, -42.15031, 
        -42.18852, -42.22364, -42.2572, -42.28841, -42.31721, -42.34354, 
        -42.36765, -42.38921, -42.40819, -42.42493, -42.439, -42.44957, 
        -42.4563, -42.45924, -42.45876, -42.45549, -42.44938, -42.44381, 
        -42.43924, -42.43672, -42.43677, -42.43967, -42.44412, -42.44965, 
        -42.45495, -42.45923, -42.46185, -42.46207, -42.46004, -42.45588, 
        -42.44995, -42.44398, -42.43701, -42.4325, -42.42951, -42.4283, 
        -42.42922, -42.432, -42.43601, -42.44126, -42.44784, -42.45587, 
        -42.46522, -42.47552, -42.48691, -42.49894, -42.51106, -42.52288, 
        -42.53416, -42.54428, -42.55499, -42.56608, -42.57718, -42.58885, 
        -42.60117, -42.61454, -42.6287, -42.64342, -42.65865, -42.67324, 
        -42.68732, -42.70119, -42.71556, -42.73066, -42.74691, -42.76386, 
        -42.78143, -42.79894, -42.81831, -42.83859, -42.85968, -42.88183, 
        -42.90444, -42.92757, -42.95215, -42.9783, -43.00636, -43.0362, 
        -43.06739, -43.09914, -43.13089, -43.16196, -43.19185, -43.22025, 
        -43.2473, -43.27316, -43.29726, -43.32177, -43.34594, -43.37011, 
        -43.39466, -43.41945, -43.44432, -43.46924, -43.49368, -43.51677, 
        -43.53818, -43.55752, -43.57546, -43.59204, -43.60715, -43.62142, 
        -43.63554, -43.64961, -43.66442, -43.67975, -43.69402, -43.70948, 
        -43.72471, -43.73944, -43.75401, -43.76802, -43.78125, -43.79353, 
        -43.80478, -43.81486, -43.82414, -43.83286, -43.84108, -43.84887, 
        -43.85637, -43.86357, -43.8705, -43.87717, -43.88345, -43.88906, 
        -43.89474, -43.89897, -43.90424, -43.90922, -43.91365, -43.91731, 
        -43.91995, -43.92165, -43.9226, -43.92311, -43.92371, -43.92462, 
        -43.92636, -43.92891, -43.93187, -43.93509, -43.93827, -43.94121, 
        -43.94357, -43.94533, -43.94612, -43.94591, -43.94573, -43.94593, 
        -43.94658, -43.94602, -43.94591, -43.94458, -43.94189, -43.93755, 
        -43.93177, -43.92522, -43.91775, -43.90988, -43.90205, -43.89373, 
        -43.88465, -43.87461, -43.86297, -43.84972, -43.83517, -43.81926, 
        -43.8021, -43.78364, -43.76468, -43.74537, -43.72694, -43.70918, 
        -43.69266, -43.67663, -43.6611, -43.64499, -43.62988, -43.61449, 
        -43.59844, -43.58192, -43.56584, -43.55074, -43.5368, -43.52402, 
        -43.51216, -43.50083, -43.48948, -43.47799, -43.46521, -43.45238, 
        -43.43924, -43.42644, -43.41415, -43.40173, -43.38913, -43.3759, 
        -43.36247, -43.34905, -43.33548, -43.32168, -43.30733, -43.2924, 
        -43.27703, -43.26093, -43.24443, -43.22845, -43.21174, -43.19719, 
        -43.18382, -43.17101, -43.15845, -43.14522, -43.13102, -43.11623, 
        -43.10165, -43.08782, -43.07495, -43.06371, -43.05441, -43.04749, 
        -43.04307, -43.04072, -43.03989, -43.0401, -43.04122, -43.04341, 
        -43.04596, -43.04887, -43.05273, -43.05762, -43.06405, -43.07169, 
        -43.08032, -43.08947, -43.09835, -43.10709, -43.11531, -43.12363, 
        -43.13229, -43.14091, -43.14947, -43.15797, -43.16675, -43.17514, 
        -43.18476, -43.19442, -43.20345, -43.21087, -43.21553, -43.21624, 
        -43.21251, -43.20401, -43.19025, -43.17053, -43.14342, -43.10783, 
        -43.06211, -43.00467, -42.93338, -42.84698, -42.74458, -42.62621, 
        -42.49355, -42.34968, -42.19979, -42.04932, -41.90488, -41.77032, 
        -41.64776, -41.53709, -41.43724, -41.34594, -41.26055, -41.17847, 
        -41.09656,
  -41.10292, -41.14755, -41.19321, -41.24012, -41.28773, -41.33412, 
        -41.3817, -41.42926, -41.47697, -41.52447, -41.57162, -41.61793, 
        -41.66333, -41.70731, -41.74965, -41.79073, -41.83095, -41.87096, 
        -41.91113, -41.95184, -41.99189, -42.03279, -42.07329, -42.11283, 
        -42.1507, -42.18639, -42.21951, -42.25018, -42.27819, -42.30383, 
        -42.32707, -42.34753, -42.3653, -42.38041, -42.39273, -42.40068, 
        -42.40633, -42.40835, -42.40741, -42.40389, -42.39889, -42.39369, 
        -42.38939, -42.38687, -42.38665, -42.38898, -42.39323, -42.39865, 
        -42.40404, -42.40842, -42.4109, -42.41045, -42.40891, -42.40561, 
        -42.40121, -42.39674, -42.3931, -42.3908, -42.39004, -42.39072, 
        -42.39283, -42.39669, -42.40154, -42.40795, -42.41543, -42.42476, 
        -42.43545, -42.44704, -42.45801, -42.47026, -42.4823, -42.49401, 
        -42.50542, -42.5167, -42.52808, -42.54016, -42.55246, -42.56527, 
        -42.5784, -42.59243, -42.6071, -42.62206, -42.63692, -42.65145, 
        -42.66535, -42.67807, -42.69167, -42.70604, -42.72141, -42.7378, 
        -42.75496, -42.77322, -42.79265, -42.81347, -42.83505, -42.85791, 
        -42.88138, -42.90552, -42.93031, -42.95645, -42.98444, -43.01429, 
        -43.04561, -43.07693, -43.10926, -43.14095, -43.17138, -43.20005, 
        -43.22694, -43.25227, -43.27635, -43.29974, -43.32252, -43.34515, 
        -43.36786, -43.39096, -43.4141, -43.43733, -43.46013, -43.48216, 
        -43.50236, -43.52092, -43.53763, -43.55217, -43.5665, -43.58007, 
        -43.5932, -43.60662, -43.62062, -43.63514, -43.65004, -43.66522, 
        -43.67994, -43.69457, -43.70874, -43.7224, -43.73539, -43.74763, 
        -43.75899, -43.7697, -43.77968, -43.78939, -43.79911, -43.80878, 
        -43.81722, -43.82631, -43.83497, -43.84308, -43.85068, -43.8577, 
        -43.86419, -43.87062, -43.87677, -43.8829, -43.88855, -43.89341, 
        -43.89751, -43.90049, -43.90277, -43.90457, -43.90644, -43.90862, 
        -43.91117, -43.9143, -43.91784, -43.92143, -43.92461, -43.92647, 
        -43.92863, -43.9305, -43.93179, -43.93268, -43.93363, -43.93505, 
        -43.93668, -43.93818, -43.93874, -43.93782, -43.93532, -43.93135, 
        -43.92626, -43.92033, -43.91385, -43.90709, -43.90021, -43.89281, 
        -43.88467, -43.87525, -43.86441, -43.85221, -43.8389, -43.82415, 
        -43.80724, -43.79029, -43.77258, -43.75478, -43.73746, -43.72091, 
        -43.70514, -43.68982, -43.67464, -43.65976, -43.64494, -43.62987, 
        -43.61452, -43.59927, -43.58453, -43.57051, -43.55769, -43.54597, 
        -43.53479, -43.52403, -43.5132, -43.50163, -43.48899, -43.47568, 
        -43.46198, -43.44848, -43.43531, -43.42209, -43.40887, -43.39454, 
        -43.38124, -43.36781, -43.35407, -43.33995, -43.32537, -43.31047, 
        -43.29523, -43.27968, -43.26424, -43.24945, -43.23559, -43.22326, 
        -43.21215, -43.20192, -43.19171, -43.18087, -43.16956, -43.15785, 
        -43.14578, -43.13393, -43.12271, -43.11278, -43.10452, -43.09826, 
        -43.0942, -43.09214, -43.09093, -43.09086, -43.09143, -43.09278, 
        -43.09408, -43.09587, -43.09801, -43.1002, -43.10454, -43.10995, 
        -43.11662, -43.12374, -43.1308, -43.13734, -43.14369, -43.14997, 
        -43.15625, -43.1623, -43.16823, -43.17427, -43.18074, -43.18755, 
        -43.19497, -43.20263, -43.20981, -43.21519, -43.21747, -43.21567, 
        -43.20935, -43.19811, -43.18179, -43.16003, -43.13147, -43.09474, 
        -43.04831, -42.99123, -42.92067, -42.83543, -42.73447, -42.61749, 
        -42.48574, -42.34174, -42.19033, -42.03768, -41.88936, -41.75071, 
        -41.62422, -41.51054, -41.40883, -41.31727, -41.2331, -41.15343, 
        -41.07425,
  -41.05631, -41.10042, -41.14673, -41.19396, -41.24156, -41.28887, 
        -41.33629, -41.38353, -41.43078, -41.47801, -41.525, -41.57156, 
        -41.61742, -41.66203, -41.70522, -41.74578, -41.78635, -41.82638, 
        -41.8666, -41.90714, -41.94812, -41.98886, -42.02896, -42.06813, 
        -42.10537, -42.14046, -42.17302, -42.20323, -42.2309, -42.25606, 
        -42.27749, -42.29728, -42.31406, -42.32803, -42.339, -42.34688, 
        -42.35164, -42.35358, -42.35257, -42.34954, -42.34534, -42.34099, 
        -42.33736, -42.33544, -42.33544, -42.33749, -42.34047, -42.3457, 
        -42.35105, -42.35557, -42.35809, -42.35896, -42.35815, -42.35596, 
        -42.35321, -42.35081, -42.34942, -42.34937, -42.35086, -42.35339, 
        -42.35686, -42.3614, -42.3661, -42.37324, -42.38186, -42.39212, 
        -42.40368, -42.41591, -42.42818, -42.44021, -42.45189, -42.46317, 
        -42.47412, -42.4853, -42.49731, -42.50989, -42.52313, -42.53679, 
        -42.55104, -42.56467, -42.57969, -42.59496, -42.60987, -42.62427, 
        -42.63823, -42.65174, -42.66513, -42.67907, -42.6936, -42.70935, 
        -42.72625, -42.74427, -42.76375, -42.78464, -42.80678, -42.82988, 
        -42.85413, -42.87746, -42.90232, -42.92807, -42.95555, -42.98477, 
        -43.01577, -43.04783, -43.08028, -43.11214, -43.14273, -43.17144, 
        -43.19797, -43.22243, -43.24536, -43.2672, -43.28851, -43.30937, 
        -43.3303, -43.35163, -43.37238, -43.39425, -43.41565, -43.43642, 
        -43.45592, -43.47382, -43.48989, -43.50455, -43.51839, -43.53134, 
        -43.54405, -43.55671, -43.56992, -43.58384, -43.59807, -43.61246, 
        -43.62674, -43.64063, -43.65436, -43.66734, -43.68013, -43.69133, 
        -43.70291, -43.71409, -43.72498, -43.73587, -43.74695, -43.75811, 
        -43.76911, -43.77968, -43.78979, -43.79933, -43.8083, -43.81658, 
        -43.82436, -43.83187, -43.83932, -43.84647, -43.85325, -43.85963, 
        -43.86483, -43.86934, -43.87293, -43.87513, -43.8784, -43.88174, 
        -43.88531, -43.88885, -43.89296, -43.89688, -43.90014, -43.9028, 
        -43.90527, -43.90765, -43.90934, -43.91139, -43.9134, -43.91579, 
        -43.91851, -43.92071, -43.92196, -43.9216, -43.91963, -43.91611, 
        -43.91146, -43.90604, -43.9004, -43.89359, -43.88774, -43.8808, 
        -43.87329, -43.86473, -43.85464, -43.84347, -43.83099, -43.81732, 
        -43.8026, -43.7868, -43.77033, -43.75351, -43.73742, -43.72201, 
        -43.70698, -43.69201, -43.67725, -43.66262, -43.64825, -43.63372, 
        -43.61934, -43.60516, -43.59174, -43.57901, -43.56737, -43.55628, 
        -43.54571, -43.5345, -43.52414, -43.51267, -43.50018, -43.48687, 
        -43.47307, -43.45926, -43.44531, -43.43162, -43.418, -43.40468, 
        -43.39125, -43.37757, -43.36371, -43.34912, -43.33429, -43.31919, 
        -43.30434, -43.28972, -43.27559, -43.26255, -43.25091, -43.24094, 
        -43.23246, -43.22449, -43.21661, -43.20826, -43.19971, -43.1905, 
        -43.18057, -43.1706, -43.16094, -43.15112, -43.14365, -43.13815, 
        -43.13431, -43.13187, -43.13038, -43.1298, -43.12993, -43.13026, 
        -43.13073, -43.13144, -43.13223, -43.13404, -43.1368, -43.14094, 
        -43.14594, -43.15147, -43.15689, -43.16218, -43.167, -43.17149, 
        -43.17543, -43.17916, -43.18284, -43.18663, -43.19068, -43.19522, 
        -43.20065, -43.20644, -43.21162, -43.21488, -43.21503, -43.21076, 
        -43.2021, -43.18891, -43.17069, -43.1474, -43.11716, -43.07936, 
        -43.03268, -42.97432, -42.90453, -42.82054, -42.72114, -42.60603, 
        -42.47575, -42.33259, -42.18081, -42.02588, -41.87456, -41.73187, 
        -41.60127, -41.48384, -41.37927, -41.28604, -41.20149, -41.12266, 
        -41.04656,
  -41.00103, -41.04707, -41.09406, -41.14159, -41.1891, -41.23647, 
        -41.28338, -41.33035, -41.37712, -41.424, -41.46992, -41.51663, 
        -41.56278, -41.60788, -41.65161, -41.69361, -41.73444, -41.77485, 
        -41.81507, -41.85572, -41.89641, -41.9368, -41.97633, -42.01456, 
        -42.05088, -42.08416, -42.11626, -42.14605, -42.17353, -42.19859, 
        -42.22086, -42.24022, -42.2564, -42.26944, -42.27963, -42.28678, 
        -42.29138, -42.2933, -42.29293, -42.29082, -42.28677, -42.28368, 
        -42.28131, -42.28034, -42.28065, -42.28283, -42.28669, -42.29162, 
        -42.29685, -42.30138, -42.30425, -42.30558, -42.30561, -42.30472, 
        -42.30397, -42.30366, -42.30369, -42.30603, -42.30951, -42.31378, 
        -42.3186, -42.32384, -42.33025, -42.33803, -42.34748, -42.35843, 
        -42.37038, -42.38292, -42.39523, -42.40669, -42.41755, -42.42809, 
        -42.4385, -42.44831, -42.46036, -42.4734, -42.4874, -42.50184, 
        -42.51664, -42.53208, -42.54759, -42.56322, -42.57839, -42.59274, 
        -42.60664, -42.62025, -42.63367, -42.64714, -42.66113, -42.67619, 
        -42.69284, -42.70992, -42.7294, -42.75033, -42.77256, -42.79575, 
        -42.81986, -42.84431, -42.86898, -42.89423, -42.92046, -42.94863, 
        -42.97879, -43.00998, -43.04173, -43.07335, -43.10383, -43.13239, 
        -43.15839, -43.18186, -43.20238, -43.22256, -43.24209, -43.26147, 
        -43.28118, -43.30117, -43.32152, -43.34229, -43.36271, -43.38254, 
        -43.4012, -43.41848, -43.43422, -43.44857, -43.46183, -43.47452, 
        -43.4867, -43.49884, -43.51143, -43.52443, -43.53687, -43.55043, 
        -43.56379, -43.577, -43.58995, -43.60246, -43.61482, -43.6271, 
        -43.63901, -43.65069, -43.66246, -43.67442, -43.68672, -43.69901, 
        -43.71128, -43.72322, -43.73447, -43.74523, -43.75546, -43.76516, 
        -43.7743, -43.78204, -43.7908, -43.79923, -43.80712, -43.8146, 
        -43.82122, -43.82693, -43.83197, -43.83651, -43.84092, -43.84541, 
        -43.84983, -43.85439, -43.8587, -43.86267, -43.86649, -43.86953, 
        -43.87229, -43.87488, -43.87748, -43.8804, -43.88362, -43.88705, 
        -43.89069, -43.89281, -43.89478, -43.89508, -43.89372, -43.89085, 
        -43.88709, -43.88243, -43.87765, -43.87276, -43.86706, -43.86094, 
        -43.85383, -43.84581, -43.83632, -43.82585, -43.81422, -43.80169, 
        -43.78782, -43.77283, -43.75736, -43.74181, -43.7266, -43.71196, 
        -43.69746, -43.68304, -43.66874, -43.65364, -43.63974, -43.62592, 
        -43.61256, -43.59981, -43.58756, -43.57616, -43.56512, -43.55478, 
        -43.54485, -43.53503, -43.52471, -43.51342, -43.50139, -43.48821, 
        -43.47451, -43.46056, -43.4464, -43.43207, -43.41825, -43.4049, 
        -43.39132, -43.37743, -43.36331, -43.34848, -43.33341, -43.31857, 
        -43.30433, -43.29093, -43.2785, -43.26758, -43.2575, -43.24998, 
        -43.24384, -43.23822, -43.23268, -43.22684, -43.2205, -43.21324, 
        -43.20544, -43.19738, -43.18903, -43.18123, -43.1745, -43.16925, 
        -43.16537, -43.16245, -43.16053, -43.15949, -43.15876, -43.15833, 
        -43.15775, -43.15748, -43.15744, -43.15821, -43.16014, -43.16327, 
        -43.16728, -43.17164, -43.17603, -43.18024, -43.18386, -43.18667, 
        -43.18888, -43.19065, -43.19231, -43.19389, -43.19453, -43.19699, 
        -43.20061, -43.20451, -43.20765, -43.20886, -43.20681, -43.20085, 
        -43.19056, -43.17577, -43.15636, -43.13171, -43.10079, -43.06198, 
        -43.01466, -42.95704, -42.88759, -42.80437, -42.7065, -42.59326, 
        -42.46466, -42.32281, -42.17125, -42.01532, -41.86162, -41.71553, 
        -41.58098, -41.45951, -41.35156, -41.25563, -41.1696, -41.09035, 
        -41.01482,
  -40.93847, -40.98518, -41.03275, -41.08058, -41.12811, -41.17435, 
        -41.22102, -41.26757, -41.31412, -41.36095, -41.40798, -41.45492, 
        -41.50131, -41.54663, -41.59043, -41.63295, -41.67414, -41.71476, 
        -41.75536, -41.7961, -41.83551, -41.87548, -41.91402, -41.95101, 
        -41.98621, -42.01958, -42.05117, -42.08083, -42.10847, -42.13362, 
        -42.15588, -42.17504, -42.19094, -42.20368, -42.21349, -42.21941, 
        -42.224, -42.22647, -42.22704, -42.22604, -42.22435, -42.22267, 
        -42.22187, -42.22195, -42.22314, -42.22557, -42.22945, -42.23418, 
        -42.2393, -42.24379, -42.24731, -42.24844, -42.24949, -42.2502, 
        -42.25124, -42.25327, -42.2564, -42.26092, -42.26631, -42.27227, 
        -42.27822, -42.28418, -42.29126, -42.29961, -42.30977, -42.32124, 
        -42.33329, -42.34454, -42.35643, -42.36723, -42.37719, -42.38724, 
        -42.39699, -42.40755, -42.4194, -42.43246, -42.44651, -42.4615, 
        -42.47698, -42.49295, -42.50922, -42.52528, -42.54059, -42.5552, 
        -42.56894, -42.58153, -42.59499, -42.60843, -42.62195, -42.6368, 
        -42.65313, -42.67124, -42.69064, -42.71136, -42.73339, -42.75631, 
        -42.77994, -42.80413, -42.82827, -42.85284, -42.87805, -42.90499, 
        -42.9333, -42.96219, -42.99278, -43.02357, -43.05342, -43.08172, 
        -43.10708, -43.12952, -43.14963, -43.16828, -43.18625, -43.20451, 
        -43.22315, -43.24244, -43.26192, -43.28167, -43.30138, -43.32036, 
        -43.33828, -43.35487, -43.37023, -43.38334, -43.39646, -43.40862, 
        -43.42044, -43.43207, -43.44388, -43.45599, -43.4685, -43.481, 
        -43.49358, -43.5059, -43.51822, -43.53008, -43.54235, -43.55453, 
        -43.56698, -43.57928, -43.59189, -43.6048, -43.61815, -43.63156, 
        -43.64379, -43.65661, -43.66879, -43.68057, -43.69177, -43.70263, 
        -43.71318, -43.72359, -43.73359, -43.74308, -43.75229, -43.76065, 
        -43.76809, -43.77502, -43.78127, -43.78714, -43.79284, -43.79841, 
        -43.80402, -43.80918, -43.81414, -43.81864, -43.82279, -43.82555, 
        -43.82874, -43.83183, -43.83535, -43.83934, -43.84367, -43.84821, 
        -43.85281, -43.85678, -43.85973, -43.86097, -43.86069, -43.85894, 
        -43.85577, -43.85216, -43.84818, -43.84367, -43.83851, -43.83282, 
        -43.82633, -43.81889, -43.8102, -43.80032, -43.78961, -43.77768, 
        -43.76349, -43.74915, -43.73447, -43.71986, -43.70576, -43.69157, 
        -43.67756, -43.66365, -43.64994, -43.63626, -43.62298, -43.61008, 
        -43.59803, -43.58663, -43.57578, -43.56511, -43.55493, -43.54508, 
        -43.53539, -43.52568, -43.51521, -43.50407, -43.49217, -43.47939, 
        -43.46604, -43.45199, -43.43743, -43.42304, -43.40913, -43.39439, 
        -43.38089, -43.36694, -43.35261, -43.33801, -43.32332, -43.30914, 
        -43.2961, -43.28419, -43.27399, -43.2655, -43.25884, -43.2536, 
        -43.24964, -43.24607, -43.24257, -43.23899, -43.2346, -43.22927, 
        -43.22321, -43.21656, -43.20947, -43.20266, -43.19649, -43.19122, 
        -43.18702, -43.18378, -43.18151, -43.17984, -43.17819, -43.17671, 
        -43.17537, -43.17419, -43.17331, -43.1725, -43.17399, -43.17645, 
        -43.17966, -43.18321, -43.18694, -43.19022, -43.1927, -43.19441, 
        -43.19526, -43.19576, -43.19556, -43.19489, -43.19442, -43.19489, 
        -43.1964, -43.19831, -43.19935, -43.19863, -43.19501, -43.18793, 
        -43.17673, -43.1613, -43.14123, -43.11589, -43.08408, -43.04444, 
        -42.99646, -42.93839, -42.86871, -42.78605, -42.68921, -42.57742, 
        -42.4506, -42.31046, -42.15978, -42.00381, -41.84869, -41.70019, 
        -41.56213, -41.43699, -41.32553, -41.22667, -41.13823, -41.05661, 
        -40.98078,
  -40.866, -40.91238, -40.96071, -41.00904, -41.05686, -41.10406, 
        -41.15087, -41.1974, -41.24383, -41.29049, -41.33746, -41.38436, 
        -41.43076, -41.47608, -41.52032, -41.56211, -41.60394, -41.64527, 
        -41.68633, -41.72718, -41.76746, -41.80646, -41.84393, -41.87964, 
        -41.91369, -41.94624, -41.97726, -42.0066, -42.0342, -42.05964, 
        -42.08124, -42.10057, -42.11667, -42.12948, -42.13929, -42.14655, 
        -42.15143, -42.15454, -42.15607, -42.15628, -42.15593, -42.15602, 
        -42.15657, -42.15799, -42.16037, -42.1636, -42.16673, -42.17161, 
        -42.17665, -42.18127, -42.1853, -42.18848, -42.19091, -42.19326, 
        -42.19614, -42.20018, -42.20556, -42.21208, -42.21915, -42.22629, 
        -42.23343, -42.24017, -42.24657, -42.25539, -42.26587, -42.27714, 
        -42.28916, -42.3007, -42.31171, -42.32199, -42.3315, -42.34086, 
        -42.35042, -42.36072, -42.37244, -42.38511, -42.39927, -42.41443, 
        -42.43036, -42.44596, -42.46273, -42.47912, -42.49467, -42.50942, 
        -42.52324, -42.53646, -42.54971, -42.56296, -42.57677, -42.59156, 
        -42.60772, -42.62569, -42.64524, -42.66573, -42.68708, -42.70942, 
        -42.7322, -42.75445, -42.77806, -42.80181, -42.82622, -42.85207, 
        -42.87897, -42.90723, -42.93645, -42.96605, -42.99509, -43.02244, 
        -43.04712, -43.06861, -43.08754, -43.10496, -43.12191, -43.13932, 
        -43.15726, -43.17582, -43.19382, -43.21284, -43.23169, -43.25006, 
        -43.26719, -43.28311, -43.2978, -43.31157, -43.3244, -43.33628, 
        -43.34761, -43.35892, -43.37021, -43.38168, -43.39323, -43.40501, 
        -43.41629, -43.42783, -43.43934, -43.45106, -43.46292, -43.47459, 
        -43.48721, -43.50007, -43.51334, -43.52715, -43.54128, -43.55553, 
        -43.56946, -43.58291, -43.5959, -43.60842, -43.62075, -43.63248, 
        -43.64433, -43.65619, -43.66768, -43.67839, -43.68856, -43.6979, 
        -43.70616, -43.71387, -43.72104, -43.72695, -43.73375, -43.74037, 
        -43.74681, -43.75278, -43.75864, -43.76394, -43.76913, -43.77374, 
        -43.77818, -43.78253, -43.78727, -43.79224, -43.79742, -43.80263, 
        -43.80782, -43.81235, -43.81612, -43.81832, -43.81908, -43.81839, 
        -43.81615, -43.81365, -43.81059, -43.80562, -43.80087, -43.7956, 
        -43.7897, -43.78297, -43.7753, -43.76624, -43.75628, -43.74517, 
        -43.73265, -43.71909, -43.70542, -43.69151, -43.67793, -43.66437, 
        -43.65083, -43.63744, -43.62418, -43.61116, -43.59884, -43.58713, 
        -43.57642, -43.56615, -43.55641, -43.54675, -43.53713, -43.52755, 
        -43.51771, -43.50671, -43.49607, -43.48481, -43.47301, -43.46067, 
        -43.44743, -43.43357, -43.41933, -43.40528, -43.3913, -43.37758, 
        -43.3639, -43.34993, -43.33597, -43.32163, -43.30774, -43.29482, 
        -43.28297, -43.27325, -43.26536, -43.25898, -43.25484, -43.25168, 
        -43.24943, -43.24768, -43.24619, -43.24424, -43.24156, -43.23793, 
        -43.2334, -43.22811, -43.22229, -43.21532, -43.2094, -43.2039, 
        -43.19924, -43.19571, -43.19307, -43.19065, -43.18845, -43.18628, 
        -43.1842, -43.18245, -43.18102, -43.18064, -43.18134, -43.18306, 
        -43.18573, -43.18882, -43.1917, -43.1941, -43.19605, -43.19716, 
        -43.19738, -43.19661, -43.19477, -43.19225, -43.18998, -43.1884, 
        -43.18751, -43.18716, -43.18641, -43.18415, -43.1794, -43.17182, 
        -43.16051, -43.14488, -43.12433, -43.09835, -43.06561, -43.02528, 
        -42.97627, -42.91649, -42.84675, -42.76446, -42.66857, -42.55807, 
        -42.43287, -42.29451, -42.1453, -41.98987, -41.83423, -41.68407, 
        -41.54345, -41.41514, -41.30034, -41.19845, -41.10733, -41.02489, 
        -40.94764,
  -40.78221, -40.83046, -40.87929, -40.92798, -40.97665, -41.02406, 
        -41.0709, -41.11787, -41.1644, -41.2112, -41.25696, -41.30392, 
        -41.35003, -41.39558, -41.44002, -41.48349, -41.52612, -41.56821, 
        -41.60985, -41.65069, -41.69053, -41.72858, -41.76506, -41.79967, 
        -41.83254, -41.86319, -41.89346, -41.92258, -41.95004, -41.97556, 
        -41.99833, -42.01822, -42.03459, -42.04797, -42.05812, -42.06596, 
        -42.07167, -42.07557, -42.07793, -42.07943, -42.07967, -42.08128, 
        -42.08356, -42.08651, -42.0903, -42.09483, -42.09977, -42.10504, 
        -42.1104, -42.11526, -42.11968, -42.12384, -42.12786, -42.13182, 
        -42.1366, -42.14229, -42.14841, -42.15667, -42.16516, -42.17358, 
        -42.18118, -42.1887, -42.19668, -42.20564, -42.21601, -42.22742, 
        -42.23867, -42.24969, -42.26018, -42.26973, -42.27882, -42.28791, 
        -42.29757, -42.30666, -42.3179, -42.33036, -42.34409, -42.35924, 
        -42.37536, -42.39242, -42.40975, -42.42644, -42.44242, -42.4571, 
        -42.47087, -42.48397, -42.49682, -42.50999, -42.52404, -42.53925, 
        -42.55555, -42.57244, -42.59186, -42.61207, -42.63274, -42.65409, 
        -42.676, -42.69825, -42.721, -42.74425, -42.76806, -42.79285, 
        -42.81853, -42.84523, -42.87293, -42.90118, -42.92923, -42.95546, 
        -42.97903, -42.99978, -43.01674, -43.03321, -43.04927, -43.06602, 
        -43.08366, -43.10193, -43.12044, -43.13897, -43.15707, -43.17447, 
        -43.19094, -43.20604, -43.22001, -43.23297, -43.24553, -43.25706, 
        -43.26821, -43.27889, -43.28971, -43.30064, -43.31046, -43.32121, 
        -43.33158, -43.34227, -43.35329, -43.36493, -43.37696, -43.38963, 
        -43.40262, -43.41614, -43.4299, -43.44433, -43.45916, -43.47394, 
        -43.48844, -43.50248, -43.51593, -43.52885, -43.54173, -43.55481, 
        -43.56787, -43.57978, -43.59229, -43.60437, -43.61562, -43.62565, 
        -43.6346, -43.64287, -43.65063, -43.65828, -43.66578, -43.67323, 
        -43.68037, -43.68744, -43.69432, -43.70113, -43.70755, -43.71368, 
        -43.71969, -43.72559, -43.7314, -43.73734, -43.74339, -43.74915, 
        -43.75491, -43.75911, -43.76347, -43.76654, -43.76826, -43.76858, 
        -43.76764, -43.76586, -43.76353, -43.76049, -43.75666, -43.75218, 
        -43.74712, -43.74132, -43.73444, -43.72668, -43.71758, -43.70719, 
        -43.69565, -43.68337, -43.67048, -43.65718, -43.64392, -43.63081, 
        -43.61774, -43.60488, -43.59215, -43.57892, -43.56755, -43.55708, 
        -43.54766, -43.53862, -43.52985, -43.52063, -43.51139, -43.50191, 
        -43.49182, -43.48126, -43.47039, -43.45903, -43.44732, -43.43495, 
        -43.42218, -43.40899, -43.39551, -43.38179, -43.36792, -43.3543, 
        -43.34069, -43.32711, -43.31339, -43.30009, -43.28733, -43.27571, 
        -43.26597, -43.25813, -43.25262, -43.248, -43.24539, -43.24373, 
        -43.24305, -43.24265, -43.24243, -43.24174, -43.24037, -43.23823, 
        -43.23524, -43.23138, -43.22686, -43.22162, -43.21581, -43.21012, 
        -43.20533, -43.20142, -43.19824, -43.19543, -43.19288, -43.19041, 
        -43.188, -43.18575, -43.18399, -43.18266, -43.18266, -43.18378, 
        -43.1857, -43.18805, -43.19009, -43.19186, -43.19315, -43.19389, 
        -43.19345, -43.19165, -43.1888, -43.18513, -43.18021, -43.17664, 
        -43.17355, -43.17112, -43.16859, -43.165, -43.15988, -43.15216, 
        -43.14112, -43.12563, -43.10509, -43.07848, -43.04491, -43.00359, 
        -42.95369, -42.89434, -42.82431, -42.74224, -42.64719, -42.53782, 
        -42.41428, -42.27737, -42.12993, -41.9756, -41.82016, -41.66895, 
        -41.52652, -41.39563, -41.27795, -41.17311, -41.07953, -40.99495, 
        -40.91635,
  -40.68935, -40.73812, -40.7879, -40.83735, -40.88633, -40.93385, 
        -40.98113, -41.02805, -41.07484, -41.12175, -41.16859, -41.21503, 
        -41.26124, -41.30685, -41.35169, -41.39574, -41.43927, -41.48216, 
        -41.52436, -41.56531, -41.60351, -41.64078, -41.6763, -41.70982, 
        -41.74172, -41.77244, -41.80211, -41.83066, -41.85789, -41.88322, 
        -41.90637, -41.9266, -41.94365, -41.95763, -41.96865, -41.97635, 
        -41.98285, -41.98753, -41.99109, -41.99379, -41.99654, -41.99989, 
        -42.0038, -42.0087, -42.01448, -42.02053, -42.02666, -42.03272, 
        -42.0384, -42.04391, -42.04897, -42.05314, -42.05853, -42.06411, 
        -42.07027, -42.07743, -42.08577, -42.09526, -42.10526, -42.11443, 
        -42.12276, -42.13051, -42.13871, -42.14796, -42.15815, -42.16904, 
        -42.18002, -42.1895, -42.19927, -42.20832, -42.21695, -42.2259, 
        -42.2355, -42.24577, -42.25681, -42.26906, -42.28256, -42.29759, 
        -42.31401, -42.33135, -42.34899, -42.36611, -42.38202, -42.39672, 
        -42.41038, -42.42215, -42.435, -42.44814, -42.46254, -42.47816, 
        -42.49483, -42.51279, -42.53196, -42.55192, -42.57202, -42.59256, 
        -42.61321, -42.63481, -42.65685, -42.6797, -42.70304, -42.7272, 
        -42.75192, -42.77654, -42.80295, -42.82972, -42.85664, -42.88217, 
        -42.90444, -42.92416, -42.94142, -42.95675, -42.97238, -42.98862, 
        -43.00576, -43.02375, -43.04198, -43.05997, -43.07729, -43.09369, 
        -43.10921, -43.12341, -43.13654, -43.14764, -43.15928, -43.17048, 
        -43.18139, -43.19189, -43.20216, -43.21253, -43.22266, -43.23262, 
        -43.24247, -43.25263, -43.26324, -43.27472, -43.28693, -43.29986, 
        -43.31329, -43.32721, -43.3416, -43.3565, -43.37176, -43.38696, 
        -43.40082, -43.41524, -43.42903, -43.44247, -43.45576, -43.46943, 
        -43.48327, -43.49718, -43.51083, -43.52395, -43.53597, -43.54667, 
        -43.5562, -43.56464, -43.57263, -43.58069, -43.58873, -43.59663, 
        -43.60468, -43.61303, -43.62111, -43.62938, -43.63767, -43.64473, 
        -43.65269, -43.66031, -43.66773, -43.67467, -43.68155, -43.68803, 
        -43.6941, -43.6996, -43.70444, -43.70826, -43.7108, -43.71207, 
        -43.71208, -43.71129, -43.70999, -43.70803, -43.70536, -43.70217, 
        -43.69819, -43.69336, -43.68773, -43.6812, -43.67323, -43.6638, 
        -43.65258, -43.64139, -43.62932, -43.61687, -43.60423, -43.59145, 
        -43.57867, -43.56608, -43.55394, -43.54254, -43.53217, -43.52277, 
        -43.51417, -43.50631, -43.49823, -43.48967, -43.48035, -43.47049, 
        -43.46019, -43.44936, -43.43821, -43.42673, -43.41483, -43.4029, 
        -43.39085, -43.37857, -43.36589, -43.35262, -43.33944, -43.32493, 
        -43.3117, -43.29869, -43.28592, -43.27391, -43.26253, -43.25262, 
        -43.24498, -43.23943, -43.23584, -43.23392, -43.23277, -43.23243, 
        -43.23267, -43.23318, -43.23361, -43.23388, -43.23361, -43.23277, 
        -43.23124, -43.22887, -43.22535, -43.22069, -43.21525, -43.20971, 
        -43.20478, -43.20057, -43.19702, -43.19416, -43.19162, -43.18925, 
        -43.18682, -43.18431, -43.18206, -43.17896, -43.17812, -43.1783, 
        -43.17932, -43.18038, -43.18168, -43.1828, -43.18376, -43.18387, 
        -43.18281, -43.18042, -43.17715, -43.17272, -43.16771, -43.16255, 
        -43.1576, -43.15319, -43.14902, -43.14448, -43.13882, -43.13128, 
        -43.12063, -43.10546, -43.08482, -43.05777, -43.02337, -42.98125, 
        -42.93059, -42.87066, -42.80042, -42.71878, -42.62448, -42.51653, 
        -42.39457, -42.25966, -42.114, -41.96102, -41.80607, -41.65433, 
        -41.51027, -41.37735, -41.25708, -41.14985, -41.05378, -40.96573, 
        -40.88532,
  -40.58743, -40.6362, -40.68668, -40.73708, -40.78697, -40.83566, 
        -40.8833, -40.93034, -40.97717, -41.0239, -41.07053, -41.11691, 
        -41.16309, -41.20888, -41.25424, -41.29803, -41.34238, -41.38599, 
        -41.42851, -41.46928, -41.50794, -41.54467, -41.5791, -41.61181, 
        -41.64304, -41.67311, -41.70203, -41.73011, -41.75706, -41.78235, 
        -41.80449, -41.82497, -41.84256, -41.85721, -41.86909, -41.8789, 
        -41.88654, -41.8923, -41.89688, -41.90122, -41.90543, -41.91025, 
        -41.91629, -41.92294, -41.93061, -41.93852, -41.94518, -41.95243, 
        -41.95908, -41.96505, -41.97113, -41.9772, -41.98367, -41.99057, 
        -41.99826, -42.00651, -42.01587, -42.02608, -42.03661, -42.04664, 
        -42.05531, -42.06335, -42.07077, -42.08009, -42.09021, -42.10092, 
        -42.11141, -42.12119, -42.13028, -42.13885, -42.14717, -42.15623, 
        -42.16608, -42.17665, -42.18804, -42.20038, -42.21372, -42.22872, 
        -42.24518, -42.26167, -42.27949, -42.29668, -42.31235, -42.32692, 
        -42.34066, -42.35359, -42.3666, -42.38021, -42.39473, -42.41072, 
        -42.42796, -42.44615, -42.46521, -42.48472, -42.50451, -42.52437, 
        -42.54488, -42.56476, -42.58622, -42.60849, -42.63147, -42.65539, 
        -42.67968, -42.70411, -42.72943, -42.75518, -42.78086, -42.80503, 
        -42.82709, -42.84532, -42.86184, -42.87659, -42.89167, -42.90712, 
        -42.92389, -42.94146, -42.95821, -42.97569, -42.99228, -43.00773, 
        -43.02206, -43.03526, -43.04727, -43.05843, -43.06902, -43.07944, 
        -43.08995, -43.1002, -43.11018, -43.11978, -43.12934, -43.13883, 
        -43.14821, -43.15812, -43.16869, -43.18027, -43.19249, -43.20472, 
        -43.21864, -43.23311, -43.24797, -43.26344, -43.279, -43.29433, 
        -43.30933, -43.32399, -43.33815, -43.35184, -43.36556, -43.37953, 
        -43.39391, -43.40855, -43.42315, -43.43702, -43.44958, -43.46067, 
        -43.4703, -43.47899, -43.48745, -43.49447, -43.5028, -43.51125, 
        -43.52028, -43.52953, -43.53927, -43.54957, -43.5596, -43.56979, 
        -43.57958, -43.58912, -43.59834, -43.60685, -43.61453, -43.62153, 
        -43.62785, -43.63354, -43.63859, -43.64297, -43.64611, -43.64822, 
        -43.64925, -43.64953, -43.64913, -43.64758, -43.64649, -43.6448, 
        -43.64228, -43.63891, -43.63422, -43.62921, -43.62251, -43.61464, 
        -43.60572, -43.59573, -43.58473, -43.57317, -43.56113, -43.54868, 
        -43.5361, -43.52366, -43.51196, -43.50126, -43.49154, -43.4829, 
        -43.47536, -43.46817, -43.46049, -43.45216, -43.4429, -43.43294, 
        -43.42272, -43.41092, -43.39957, -43.38803, -43.37627, -43.36483, 
        -43.35364, -43.34219, -43.33026, -43.31791, -43.30518, -43.29229, 
        -43.2799, -43.26777, -43.25618, -43.24545, -43.23575, -43.22813, 
        -43.22252, -43.21894, -43.21733, -43.21651, -43.21648, -43.21686, 
        -43.21757, -43.2184, -43.21916, -43.21996, -43.22054, -43.22087, 
        -43.22063, -43.21957, -43.21704, -43.21211, -43.20725, -43.20221, 
        -43.19741, -43.19325, -43.18965, -43.18709, -43.18483, -43.18275, 
        -43.18052, -43.17805, -43.17508, -43.17255, -43.17054, -43.1694, 
        -43.16879, -43.16876, -43.16914, -43.16963, -43.16975, -43.16914, 
        -43.16751, -43.16518, -43.16168, -43.1571, -43.15171, -43.14548, 
        -43.13914, -43.13321, -43.12767, -43.12219, -43.1161, -43.10858, 
        -43.09811, -43.08315, -43.0623, -43.03458, -42.99973, -42.95651, 
        -42.90527, -42.84403, -42.77405, -42.69314, -42.5999, -42.49343, 
        -42.37351, -42.24082, -42.09718, -41.9458, -41.79157, -41.63961, 
        -41.4944, -41.3595, -41.23705, -41.12714, -41.02861, -40.93946, 
        -40.85739,
  -40.47594, -40.52677, -40.57833, -40.62966, -40.68016, -40.72924, 
        -40.77708, -40.82409, -40.87069, -40.91706, -40.96247, -41.00873, 
        -41.055, -41.10121, -41.1472, -41.19281, -41.23766, -41.28151, 
        -41.32395, -41.36433, -41.40265, -41.43864, -41.47267, -41.50473, 
        -41.53568, -41.5643, -41.5929, -41.62044, -41.647, -41.67217, 
        -41.69525, -41.71592, -41.73412, -41.74955, -41.76252, -41.77311, 
        -41.78175, -41.78878, -41.79483, -41.80051, -41.8054, -41.8121, 
        -41.81977, -41.82835, -41.8378, -41.84734, -41.85665, -41.86528, 
        -41.87289, -41.88007, -41.8869, -41.89408, -41.90171, -41.90993, 
        -41.91864, -41.92783, -41.93674, -41.94728, -41.95792, -41.96793, 
        -41.97683, -41.98507, -41.99376, -42.0034, -42.01369, -42.02404, 
        -42.03407, -42.04342, -42.05182, -42.06027, -42.06883, -42.07798, 
        -42.08825, -42.09858, -42.11068, -42.12333, -42.13695, -42.15195, 
        -42.1685, -42.18589, -42.20357, -42.22061, -42.23625, -42.25085, 
        -42.26451, -42.27786, -42.29115, -42.30535, -42.32053, -42.33689, 
        -42.35456, -42.37219, -42.39125, -42.41057, -42.4302, -42.45014, 
        -42.47008, -42.49059, -42.51158, -42.53351, -42.55656, -42.58014, 
        -42.60413, -42.62818, -42.65246, -42.67722, -42.70178, -42.72498, 
        -42.74597, -42.76358, -42.7779, -42.79205, -42.8064, -42.82166, 
        -42.83796, -42.85484, -42.8722, -42.88889, -42.90462, -42.91913, 
        -42.93244, -42.94436, -42.9552, -42.96516, -42.97465, -42.98399, 
        -42.9935, -43.00319, -43.01278, -43.02197, -43.0299, -43.03909, 
        -43.04826, -43.05802, -43.06878, -43.0803, -43.09299, -43.10666, 
        -43.12116, -43.13624, -43.15162, -43.16719, -43.18287, -43.19828, 
        -43.21375, -43.22849, -43.24294, -43.25724, -43.27109, -43.28534, 
        -43.29987, -43.31398, -43.32884, -43.34316, -43.35596, -43.36718, 
        -43.37706, -43.38586, -43.39466, -43.4033, -43.41196, -43.42073, 
        -43.43039, -43.44085, -43.45237, -43.46398, -43.47584, -43.48819, 
        -43.50008, -43.51182, -43.52261, -43.53272, -43.54155, -43.54887, 
        -43.55536, -43.56017, -43.56547, -43.57021, -43.57405, -43.57673, 
        -43.57848, -43.5798, -43.58076, -43.58196, -43.5826, -43.58256, 
        -43.58184, -43.57965, -43.57698, -43.57331, -43.56823, -43.56171, 
        -43.55413, -43.5455, -43.53574, -43.52522, -43.5137, -43.50166, 
        -43.48926, -43.47715, -43.46563, -43.45417, -43.4449, -43.43681, 
        -43.42992, -43.42311, -43.41578, -43.40762, -43.39852, -43.3888, 
        -43.37873, -43.36812, -43.35703, -43.34559, -43.33434, -43.32356, 
        -43.31301, -43.30228, -43.29137, -43.27996, -43.26785, -43.256, 
        -43.24448, -43.23331, -43.22301, -43.21371, -43.20608, -43.20051, 
        -43.19697, -43.19534, -43.19499, -43.19433, -43.19498, -43.1959, 
        -43.19677, -43.19745, -43.19836, -43.19941, -43.20066, -43.20179, 
        -43.20278, -43.2028, -43.20139, -43.19848, -43.19461, -43.19031, 
        -43.18585, -43.18198, -43.17893, -43.17642, -43.17451, -43.1731, 
        -43.17118, -43.16851, -43.16558, -43.16238, -43.15911, -43.15617, 
        -43.15405, -43.1527, -43.15187, -43.15125, -43.15027, -43.1489, 
        -43.14717, -43.14491, -43.14173, -43.13749, -43.13101, -43.12433, 
        -43.11715, -43.11018, -43.10366, -43.09732, -43.09074, -43.0829, 
        -43.0724, -43.05748, -43.03614, -43.0078, -42.97216, -42.92838, 
        -42.8772, -42.81706, -42.7473, -42.66717, -42.57524, -42.47062, 
        -42.35309, -42.22296, -42.08178, -41.93242, -41.77918, -41.62727, 
        -41.48123, -41.34468, -41.22004, -41.10755, -41.0066, -40.91536, 
        -40.83159,
  -40.35786, -40.40981, -40.4623, -40.51438, -40.56546, -40.614, 
        -40.66174, -40.70854, -40.75477, -40.80079, -40.84702, -40.89342, 
        -40.93996, -40.98656, -41.03314, -41.07932, -41.12454, -41.1683, 
        -41.21028, -41.24978, -41.28638, -41.32187, -41.35552, -41.38774, 
        -41.41844, -41.44818, -41.47672, -41.50404, -41.53036, -41.55538, 
        -41.57842, -41.5994, -41.61787, -41.63411, -41.64786, -41.65831, 
        -41.66805, -41.67632, -41.68385, -41.69127, -41.69899, -41.70738, 
        -41.71669, -41.72708, -41.73797, -41.74885, -41.75952, -41.76943, 
        -41.77857, -41.78693, -41.79491, -41.80204, -41.81086, -41.82029, 
        -41.83014, -41.84034, -41.85068, -41.86073, -41.87069, -41.8806, 
        -41.88956, -41.89815, -41.90728, -41.91702, -41.92754, -41.9379, 
        -41.94771, -41.9557, -41.96417, -41.97229, -41.98106, -41.99099, 
        -42.00183, -42.01396, -42.02684, -42.04037, -42.05458, -42.06993, 
        -42.08633, -42.1036, -42.12103, -42.13781, -42.15359, -42.16817, 
        -42.18213, -42.19493, -42.20918, -42.22414, -42.24001, -42.25696, 
        -42.27489, -42.29368, -42.31315, -42.33263, -42.35221, -42.37218, 
        -42.39239, -42.41274, -42.43361, -42.45535, -42.47783, -42.50113, 
        -42.52506, -42.54789, -42.57172, -42.59552, -42.61908, -42.64121, 
        -42.66094, -42.67799, -42.69268, -42.70642, -42.72002, -42.73455, 
        -42.75027, -42.76668, -42.78329, -42.79933, -42.8143, -42.82773, 
        -42.83979, -42.85051, -42.86005, -42.86772, -42.87606, -42.88414, 
        -42.89239, -42.90088, -42.90968, -42.91847, -42.92691, -42.93567, 
        -42.94498, -42.95468, -42.9654, -42.97714, -42.99026, -43.00447, 
        -43.01942, -43.03497, -43.05074, -43.06666, -43.08256, -43.09828, 
        -43.11285, -43.12814, -43.14291, -43.15739, -43.17163, -43.18612, 
        -43.2007, -43.21568, -43.23074, -43.24502, -43.25784, -43.26925, 
        -43.27931, -43.28859, -43.2976, -43.3069, -43.31604, -43.32532, 
        -43.33555, -43.34703, -43.35948, -43.37242, -43.38622, -43.39939, 
        -43.41372, -43.4271, -43.43991, -43.45129, -43.46078, -43.46886, 
        -43.47577, -43.48177, -43.48739, -43.49244, -43.49673, -43.50011, 
        -43.50281, -43.50515, -43.5077, -43.51056, -43.51313, -43.51509, 
        -43.51603, -43.516, -43.51479, -43.51252, -43.50888, -43.50382, 
        -43.49665, -43.48928, -43.48087, -43.47119, -43.46074, -43.44931, 
        -43.4373, -43.42545, -43.41402, -43.40354, -43.39437, -43.38669, 
        -43.38008, -43.37358, -43.36654, -43.35874, -43.34985, -43.34056, 
        -43.33087, -43.32084, -43.31023, -43.29938, -43.28878, -43.2785, 
        -43.26844, -43.2585, -43.24831, -43.2376, -43.22664, -43.21481, 
        -43.20422, -43.19415, -43.18528, -43.17755, -43.17191, -43.16825, 
        -43.16661, -43.1665, -43.16739, -43.16872, -43.16997, -43.17114, 
        -43.17205, -43.17273, -43.17367, -43.17492, -43.17636, -43.17817, 
        -43.17992, -43.18093, -43.18078, -43.17929, -43.17662, -43.17315, 
        -43.16944, -43.16624, -43.16365, -43.16161, -43.16014, -43.15898, 
        -43.15723, -43.15501, -43.15184, -43.14683, -43.14234, -43.13798, 
        -43.13443, -43.13165, -43.12918, -43.12698, -43.12476, -43.12293, 
        -43.12109, -43.11894, -43.11633, -43.1125, -43.10741, -43.10081, 
        -43.09346, -43.08569, -43.07834, -43.07146, -43.06434, -43.05609, 
        -43.04519, -43.0296, -43.00787, -42.97904, -42.94273, -42.89891, 
        -42.84742, -42.78765, -42.71881, -42.6396, -42.54933, -42.447, 
        -42.33228, -42.20523, -42.06697, -41.91984, -41.76809, -41.61662, 
        -41.47015, -41.33223, -41.20555, -41.09053, -40.98746, -40.8931, 
        -40.80805,
  -40.23254, -40.2848, -40.33829, -40.39115, -40.44277, -40.4924, 
        -40.54026, -40.58685, -40.63264, -40.67831, -40.72432, -40.77085, 
        -40.8177, -40.8648, -40.91186, -40.95737, -41.00255, -41.0458, 
        -41.08693, -41.12585, -41.16245, -41.19722, -41.23078, -41.26302, 
        -41.29422, -41.32423, -41.35303, -41.38052, -41.40682, -41.43157, 
        -41.45372, -41.47488, -41.49363, -41.51026, -41.52488, -41.53733, 
        -41.548, -41.55755, -41.56673, -41.57593, -41.58567, -41.59563, 
        -41.60658, -41.61815, -41.63021, -41.64222, -41.65281, -41.66398, 
        -41.67447, -41.68422, -41.69345, -41.70274, -41.71272, -41.72355, 
        -41.73465, -41.74583, -41.75612, -41.76601, -41.77522, -41.78416, 
        -41.79321, -41.80232, -41.81099, -41.82115, -41.83184, -41.84217, 
        -41.85197, -41.86089, -41.86959, -41.87807, -41.88716, -41.89771, 
        -41.90954, -41.92241, -41.93616, -41.95067, -41.96579, -41.9816, 
        -41.99844, -42.01445, -42.03171, -42.04822, -42.06401, -42.07909, 
        -42.0938, -42.10846, -42.12368, -42.13941, -42.15609, -42.17353, 
        -42.19199, -42.21113, -42.23087, -42.25068, -42.27064, -42.2906, 
        -42.31107, -42.33055, -42.35133, -42.37283, -42.39513, -42.41801, 
        -42.44172, -42.46535, -42.48899, -42.51213, -42.5346, -42.55576, 
        -42.57486, -42.59114, -42.60557, -42.61866, -42.63161, -42.64536, 
        -42.66032, -42.67617, -42.69117, -42.70652, -42.72049, -42.73291, 
        -42.74378, -42.75328, -42.76147, -42.76892, -42.77584, -42.78239, 
        -42.78924, -42.79653, -42.80402, -42.81205, -42.82023, -42.82899, 
        -42.8379, -42.84748, -42.85855, -42.87055, -42.88406, -42.89769, 
        -42.91329, -42.92933, -42.94554, -42.96157, -42.97752, -42.99348, 
        -43.00939, -43.02505, -43.04036, -43.05537, -43.06994, -43.08437, 
        -43.09888, -43.11336, -43.12805, -43.14204, -43.15474, -43.16646, 
        -43.17709, -43.18708, -43.19662, -43.20503, -43.21447, -43.22432, 
        -43.23512, -43.24709, -43.26037, -43.27464, -43.29006, -43.30601, 
        -43.32219, -43.33759, -43.35197, -43.36444, -43.37492, -43.38384, 
        -43.39117, -43.39767, -43.4037, -43.40929, -43.4141, -43.41825, 
        -43.42189, -43.42559, -43.42965, -43.43311, -43.4376, -43.44147, 
        -43.44435, -43.44604, -43.44666, -43.44588, -43.44364, -43.43988, 
        -43.43496, -43.42886, -43.42171, -43.41331, -43.40378, -43.39335, 
        -43.38213, -43.37061, -43.35932, -43.34892, -43.3399, -43.33229, 
        -43.3256, -43.31933, -43.31261, -43.30527, -43.29712, -43.28839, 
        -43.27924, -43.26872, -43.25895, -43.24884, -43.23892, -43.229, 
        -43.2194, -43.20992, -43.20022, -43.19038, -43.18051, -43.17059, 
        -43.16093, -43.15189, -43.14428, -43.13836, -43.13457, -43.13268, 
        -43.13274, -43.13403, -43.13588, -43.13806, -43.13998, -43.14138, 
        -43.14252, -43.14335, -43.14443, -43.14574, -43.14753, -43.14977, 
        -43.15191, -43.15395, -43.15404, -43.1538, -43.15216, -43.14985, 
        -43.14733, -43.145, -43.14289, -43.14138, -43.14005, -43.13914, 
        -43.13779, -43.1356, -43.13213, -43.12761, -43.12233, -43.117, 
        -43.11223, -43.10769, -43.10326, -43.09924, -43.09605, -43.09352, 
        -43.09156, -43.08971, -43.08747, -43.08438, -43.07983, -43.07378, 
        -43.06658, -43.05868, -43.05086, -43.04328, -43.03532, -43.02629, 
        -43.0146, -42.99862, -42.9763, -42.94698, -42.91016, -42.8663, 
        -42.81408, -42.75503, -42.68715, -42.60942, -42.52113, -42.42149, 
        -42.31015, -42.18679, -42.0519, -41.90762, -41.75783, -41.60728, 
        -41.46067, -41.32174, -41.19304, -41.07576, -40.97033, -40.87582, 
        -40.78951,
  -40.10052, -40.15451, -40.20866, -40.26229, -40.31426, -40.36428, 
        -40.41229, -40.45877, -40.50446, -40.55005, -40.59489, -40.6414, 
        -40.68853, -40.7359, -40.78299, -40.82946, -40.87426, -40.91689, 
        -40.95716, -40.99512, -41.03098, -41.0654, -41.09874, -41.13128, 
        -41.16294, -41.19234, -41.22136, -41.24896, -41.2752, -41.29998, 
        -41.32312, -41.34431, -41.3636, -41.38067, -41.39568, -41.40907, 
        -41.42096, -41.43191, -41.44295, -41.45397, -41.4644, -41.47565, 
        -41.48809, -41.50074, -41.51364, -41.5266, -41.53923, -41.55139, 
        -41.56289, -41.57398, -41.58447, -41.59506, -41.60623, -41.61821, 
        -41.63061, -41.64244, -41.65261, -41.66232, -41.67117, -41.6798, 
        -41.68851, -41.69809, -41.70825, -41.71902, -41.7299, -41.74042, 
        -41.75026, -41.75966, -41.76872, -41.77797, -41.7877, -41.79869, 
        -41.81105, -41.82384, -41.83837, -41.85369, -41.8699, -41.88653, 
        -41.90376, -41.92093, -41.93816, -41.95495, -41.97113, -41.98687, 
        -42.00257, -42.01833, -42.03428, -42.05056, -42.06791, -42.08614, 
        -42.10507, -42.12384, -42.14392, -42.16409, -42.18463, -42.2048, 
        -42.22532, -42.24634, -42.26711, -42.28869, -42.3107, -42.33335, 
        -42.35653, -42.38011, -42.40351, -42.4264, -42.44788, -42.46805, 
        -42.48666, -42.50261, -42.51549, -42.52815, -42.54053, -42.55354, 
        -42.56776, -42.58274, -42.59806, -42.61261, -42.62551, -42.63686, 
        -42.64654, -42.65473, -42.66175, -42.66787, -42.67345, -42.67845, 
        -42.68391, -42.68961, -42.69593, -42.70294, -42.70969, -42.7182, 
        -42.72709, -42.73698, -42.74787, -42.76009, -42.77391, -42.78902, 
        -42.80503, -42.82158, -42.83799, -42.85418, -42.87022, -42.88625, 
        -42.90229, -42.91828, -42.93387, -42.94913, -42.96402, -42.97845, 
        -42.99295, -43.00608, -43.02026, -43.03392, -43.04681, -43.0588, 
        -43.07018, -43.08081, -43.09091, -43.10073, -43.11069, -43.12077, 
        -43.13184, -43.14416, -43.1578, -43.17301, -43.1895, -43.20687, 
        -43.22453, -43.24155, -43.25724, -43.27105, -43.28278, -43.29274, 
        -43.30087, -43.30715, -43.31392, -43.32004, -43.32571, -43.3308, 
        -43.33565, -43.34058, -43.3463, -43.35248, -43.35839, -43.36388, 
        -43.36853, -43.37215, -43.37439, -43.375, -43.37431, -43.37194, 
        -43.36839, -43.3636, -43.35774, -43.35067, -43.34253, -43.33317, 
        -43.32282, -43.31195, -43.30111, -43.29015, -43.28121, -43.2736, 
        -43.26697, -43.2608, -43.25456, -43.24776, -43.24027, -43.23206, 
        -43.22349, -43.21458, -43.20551, -43.19624, -43.18694, -43.17748, 
        -43.1682, -43.15896, -43.14975, -43.1406, -43.13138, -43.12206, 
        -43.11318, -43.10554, -43.0993, -43.095, -43.0929, -43.09274, 
        -43.09407, -43.09655, -43.09985, -43.10191, -43.10424, -43.10615, 
        -43.10753, -43.10871, -43.10991, -43.11146, -43.11358, -43.11599, 
        -43.11887, -43.12142, -43.12349, -43.12446, -43.12398, -43.12268, 
        -43.12137, -43.11969, -43.11821, -43.11697, -43.11615, -43.11533, 
        -43.11425, -43.11185, -43.10821, -43.1035, -43.09788, -43.0918, 
        -43.08556, -43.07909, -43.07299, -43.06763, -43.06322, -43.06003, 
        -43.0578, -43.05617, -43.05451, -43.05205, -43.04737, -43.04204, 
        -43.03522, -43.02758, -43.01957, -43.01132, -43.00263, -42.99249, 
        -42.97991, -42.96291, -42.94011, -42.91041, -42.87365, -42.82998, 
        -42.7794, -42.72117, -42.6544, -42.57866, -42.49298, -42.39648, 
        -42.28883, -42.16936, -42.03833, -41.89738, -41.75011, -41.60106, 
        -41.4549, -41.31543, -41.18524, -41.0666, -40.95937, -40.86318, 
        -40.7765,
  -39.96465, -40.019, -40.07362, -40.12764, -40.18011, -40.22959, 
        -40.27795, -40.32447, -40.37025, -40.41575, -40.46147, -40.50777, 
        -40.55479, -40.60212, -40.64925, -40.69526, -40.73946, -40.7812, 
        -40.82058, -40.85776, -40.89201, -40.92623, -40.95959, -40.99249, 
        -41.02447, -41.05529, -41.08461, -41.11232, -41.13846, -41.16327, 
        -41.18654, -41.20784, -41.22736, -41.24508, -41.26073, -41.27389, 
        -41.28693, -41.29959, -41.31229, -41.32479, -41.33746, -41.35049, 
        -41.36375, -41.3773, -41.39106, -41.40479, -41.4183, -41.43126, 
        -41.44384, -41.45596, -41.46772, -41.47847, -41.49082, -41.50395, 
        -41.51746, -41.53043, -41.54223, -41.55242, -41.56136, -41.56998, 
        -41.57898, -41.58874, -41.59944, -41.6107, -41.62178, -41.63251, 
        -41.64277, -41.65164, -41.66135, -41.67133, -41.68208, -41.69349, 
        -41.70615, -41.72048, -41.73586, -41.7522, -41.76924, -41.78696, 
        -41.80495, -41.82264, -41.84017, -41.85738, -41.87455, -41.89125, 
        -41.90808, -41.92369, -41.94043, -41.95709, -41.97479, -41.99358, 
        -42.01339, -42.03391, -42.05463, -42.07544, -42.09645, -42.11706, 
        -42.13763, -42.1585, -42.17982, -42.20136, -42.22325, -42.24549, 
        -42.26836, -42.29066, -42.31387, -42.33662, -42.35835, -42.37799, 
        -42.39566, -42.41135, -42.42501, -42.43719, -42.44905, -42.46145, 
        -42.47461, -42.48876, -42.50296, -42.51632, -42.52832, -42.53856, 
        -42.54691, -42.5541, -42.56007, -42.56408, -42.56846, -42.57228, 
        -42.57605, -42.58044, -42.58559, -42.59159, -42.59874, -42.60699, 
        -42.61608, -42.62601, -42.63703, -42.64946, -42.66345, -42.6788, 
        -42.6949, -42.71153, -42.72802, -42.74435, -42.76035, -42.77629, 
        -42.79148, -42.80743, -42.8231, -42.83865, -42.85388, -42.86864, 
        -42.88302, -42.89677, -42.91035, -42.92353, -42.93637, -42.94897, 
        -42.96108, -42.97261, -42.98351, -42.99355, -43.00392, -43.01415, 
        -43.02533, -43.03757, -43.05124, -43.06698, -43.08442, -43.10181, 
        -43.12043, -43.13862, -43.15567, -43.17095, -43.18408, -43.1952, 
        -43.20459, -43.21289, -43.22051, -43.22756, -43.23421, -43.2404, 
        -43.24643, -43.25307, -43.26015, -43.2677, -43.27508, -43.28214, 
        -43.28846, -43.29351, -43.29755, -43.30001, -43.3008, -43.29991, 
        -43.2969, -43.29329, -43.28882, -43.2832, -43.27625, -43.26799, 
        -43.25877, -43.24883, -43.23895, -43.22935, -43.22097, -43.21356, 
        -43.20702, -43.20101, -43.19513, -43.1888, -43.18164, -43.17391, 
        -43.16592, -43.15783, -43.14956, -43.14099, -43.13228, -43.12338, 
        -43.11428, -43.10518, -43.09627, -43.08737, -43.07742, -43.06873, 
        -43.06088, -43.05433, -43.0496, -43.04686, -43.04622, -43.04731, 
        -43.04995, -43.05384, -43.058, -43.06151, -43.06459, -43.06718, 
        -43.06962, -43.07146, -43.07318, -43.07529, -43.07756, -43.08037, 
        -43.08323, -43.08641, -43.08901, -43.09068, -43.09123, -43.09105, 
        -43.09054, -43.08967, -43.08877, -43.08791, -43.08726, -43.08681, 
        -43.08544, -43.08285, -43.07833, -43.07364, -43.06787, -43.06107, 
        -43.05367, -43.04607, -43.03865, -43.03206, -43.02668, -43.02259, 
        -43.02, -43.01827, -43.01695, -43.01527, -43.01221, -43.00775, 
        -43.00176, -42.99449, -42.98655, -42.97784, -42.96824, -42.95704, 
        -42.94335, -42.92559, -42.902, -42.87208, -42.83559, -42.79247, 
        -42.74244, -42.68508, -42.61992, -42.54626, -42.46337, -42.37051, 
        -42.2669, -42.15166, -42.02483, -41.88772, -41.74346, -41.59661, 
        -41.45153, -41.31212, -41.18143, -41.0615, -40.95353, -40.85556, 
        -40.76812,
  -39.82521, -39.87827, -39.93285, -39.98698, -40.03978, -40.09053, 
        -40.13917, -40.18611, -40.23203, -40.27766, -40.32315, -40.36935, 
        -40.41605, -40.463, -40.50965, -40.55408, -40.59758, -40.63857, 
        -40.67722, -40.71386, -40.74877, -40.78294, -40.81649, -40.84962, 
        -40.88198, -40.91319, -40.94281, -40.97071, -40.99669, -41.02146, 
        -41.04397, -41.06544, -41.08522, -41.10335, -41.11972, -41.1349, 
        -41.14893, -41.16276, -41.17682, -41.19085, -41.2051, -41.21943, 
        -41.23347, -41.24769, -41.26215, -41.27658, -41.28995, -41.30383, 
        -41.31713, -41.33024, -41.34296, -41.35571, -41.3693, -41.38353, 
        -41.39795, -41.4122, -41.42499, -41.43606, -41.44591, -41.45496, 
        -41.46431, -41.47471, -41.48483, -41.49637, -41.50785, -41.51886, 
        -41.52945, -41.53995, -41.55051, -41.5612, -41.57244, -41.5844, 
        -41.59776, -41.61248, -41.6285, -41.64592, -41.66411, -41.68259, 
        -41.70132, -41.71874, -41.73701, -41.75528, -41.77359, -41.79184, 
        -41.80969, -41.82718, -41.84439, -41.86174, -41.87986, -41.89918, 
        -41.91978, -41.94118, -41.96246, -41.9836, -42.00501, -42.02591, 
        -42.04682, -42.06673, -42.08811, -42.11001, -42.13161, -42.15373, 
        -42.17635, -42.19924, -42.22242, -42.24529, -42.26708, -42.28661, 
        -42.30437, -42.31972, -42.33305, -42.34507, -42.3564, -42.36794, 
        -42.38008, -42.39295, -42.40496, -42.41725, -42.42806, -42.43708, 
        -42.44431, -42.45045, -42.45547, -42.45951, -42.4629, -42.46565, 
        -42.46845, -42.47158, -42.47559, -42.48091, -42.48756, -42.49555, 
        -42.50471, -42.51487, -42.52631, -42.53905, -42.5529, -42.56709, 
        -42.58316, -42.59952, -42.61587, -42.63179, -42.64771, -42.66353, 
        -42.67947, -42.69537, -42.71119, -42.72683, -42.74227, -42.75727, 
        -42.77169, -42.78521, -42.79826, -42.81097, -42.82375, -42.83674, 
        -42.84975, -42.86216, -42.87374, -42.88335, -42.89362, -42.90383, 
        -42.91504, -42.92714, -42.941, -42.95668, -42.97428, -42.99329, 
        -43.01267, -43.03191, -43.05011, -43.06673, -43.08146, -43.09406, 
        -43.10495, -43.1145, -43.12331, -43.13151, -43.13922, -43.14673, 
        -43.15423, -43.16227, -43.17094, -43.17894, -43.18769, -43.19626, 
        -43.20382, -43.21032, -43.2159, -43.22012, -43.22253, -43.22343, 
        -43.22283, -43.22121, -43.21799, -43.21357, -43.20774, -43.20067, 
        -43.19252, -43.18388, -43.175, -43.1664, -43.15865, -43.15171, 
        -43.14556, -43.13989, -43.13428, -43.12803, -43.12117, -43.11387, 
        -43.10545, -43.09806, -43.09053, -43.08267, -43.07415, -43.06577, 
        -43.05665, -43.04771, -43.03896, -43.03015, -43.02151, -43.01358, 
        -43.00665, -43.00127, -42.99791, -42.99662, -42.99704, -42.99924, 
        -43.00314, -43.00791, -43.01293, -43.01743, -43.02177, -43.02537, 
        -43.02849, -43.03123, -43.03377, -43.03636, -43.03891, -43.04171, 
        -43.04489, -43.04811, -43.04993, -43.05222, -43.05376, -43.0546, 
        -43.05478, -43.05471, -43.05468, -43.05369, -43.05312, -43.05258, 
        -43.05095, -43.04839, -43.04499, -43.04028, -43.03433, -43.02724, 
        -43.01938, -43.0111, -43.00281, -42.99521, -42.98883, -42.98419, 
        -42.98103, -42.97909, -42.97791, -42.97651, -42.97431, -42.97071, 
        -42.96525, -42.95856, -42.95065, -42.94175, -42.93147, -42.91963, 
        -42.90489, -42.88615, -42.86212, -42.83201, -42.7956, -42.75279, 
        -42.70242, -42.64601, -42.58234, -42.51102, -42.43119, -42.34214, 
        -42.24245, -42.13154, -42.00906, -41.87609, -41.73561, -41.59172, 
        -41.44868, -41.31026, -41.17993, -41.06008, -40.95177, -40.8546, 
        -40.7673,
  -39.68191, -39.73518, -39.78911, -39.84292, -39.89571, -39.94663, 
        -39.99564, -40.04303, -40.08934, -40.13503, -40.17952, -40.22533, 
        -40.27158, -40.31798, -40.36396, -40.40871, -40.4514, -40.49184, 
        -40.52991, -40.56626, -40.60131, -40.63541, -40.66932, -40.7029, 
        -40.73561, -40.76615, -40.79596, -40.82411, -40.85034, -40.87504, 
        -40.89851, -40.92028, -40.94024, -40.95854, -40.97552, -40.99132, 
        -41.00657, -41.02151, -41.03664, -41.05206, -41.06643, -41.08155, 
        -41.09636, -41.11151, -41.12671, -41.14204, -41.15707, -41.17199, 
        -41.18655, -41.20029, -41.2138, -41.22744, -41.24193, -41.2572, 
        -41.27288, -41.28813, -41.30112, -41.31328, -41.32411, -41.33432, 
        -41.34449, -41.35559, -41.36734, -41.37931, -41.39104, -41.40254, 
        -41.41368, -41.42459, -41.43574, -41.44725, -41.45926, -41.47198, 
        -41.48588, -41.50024, -41.51696, -41.53528, -41.5544, -41.57369, 
        -41.593, -41.61239, -41.63181, -41.65129, -41.67111, -41.6909, 
        -41.71006, -41.72828, -41.746, -41.76376, -41.78249, -41.80214, 
        -41.8233, -41.84452, -41.86662, -41.88828, -41.90968, -41.93089, 
        -41.95206, -41.97314, -41.99451, -42.01603, -42.03795, -42.06008, 
        -42.08247, -42.10522, -42.12813, -42.15103, -42.173, -42.19331, 
        -42.21122, -42.22641, -42.23867, -42.25031, -42.26143, -42.27226, 
        -42.28337, -42.29485, -42.30632, -42.31724, -42.32689, -42.33467, 
        -42.34111, -42.3463, -42.35039, -42.35358, -42.35637, -42.35858, 
        -42.36042, -42.36261, -42.36593, -42.37062, -42.37609, -42.38412, 
        -42.39335, -42.4039, -42.41556, -42.42843, -42.44241, -42.45711, 
        -42.47261, -42.48858, -42.50428, -42.51982, -42.53539, -42.55092, 
        -42.56657, -42.58208, -42.59783, -42.61354, -42.62931, -42.64449, 
        -42.6588, -42.67117, -42.68373, -42.69619, -42.70893, -42.72228, 
        -42.73576, -42.74875, -42.76064, -42.77168, -42.78213, -42.79245, 
        -42.80328, -42.81544, -42.82893, -42.84457, -42.86194, -42.88102, 
        -42.90119, -42.92117, -42.94048, -42.9586, -42.9748, -42.98903, 
        -43.00153, -43.01171, -43.02171, -43.03134, -43.04053, -43.04944, 
        -43.05876, -43.06833, -43.07845, -43.08888, -43.09904, -43.10877, 
        -43.1176, -43.12539, -43.13245, -43.13832, -43.14262, -43.14536, 
        -43.14653, -43.14633, -43.14466, -43.14141, -43.13675, -43.13072, 
        -43.1238, -43.11634, -43.10876, -43.10052, -43.09361, -43.08744, 
        -43.08207, -43.07661, -43.0712, -43.06514, -43.05851, -43.05154, 
        -43.04463, -43.03764, -43.03042, -43.02311, -43.0151, -43.00695, 
        -42.99797, -42.98909, -42.98014, -42.97159, -42.96371, -42.95665, 
        -42.95065, -42.94645, -42.94419, -42.94381, -42.94534, -42.94875, 
        -42.95346, -42.95908, -42.96506, -42.96982, -42.97522, -42.98004, 
        -42.98412, -42.98766, -42.9908, -42.99372, -42.99657, -42.99953, 
        -43.00274, -43.00577, -43.00886, -43.01181, -43.01393, -43.0157, 
        -43.01693, -43.01743, -43.01731, -43.0172, -43.01635, -43.01574, 
        -43.01394, -43.01148, -43.00779, -43.00281, -42.99691, -42.98992, 
        -42.98203, -42.97355, -42.96495, -42.95678, -42.94975, -42.94451, 
        -42.94086, -42.93879, -42.93727, -42.93602, -42.93326, -42.93033, 
        -42.92583, -42.9197, -42.9119, -42.90272, -42.8921, -42.87937, 
        -42.86388, -42.84455, -42.82021, -42.78997, -42.75354, -42.7108, 
        -42.66175, -42.60619, -42.54409, -42.47488, -42.3979, -42.31221, 
        -42.21648, -42.10972, -41.99164, -41.86313, -41.72685, -41.58668, 
        -41.44668, -41.31081, -41.18188, -41.06311, -40.9554, -40.85866, 
        -40.77168,
  -39.53722, -39.58945, -39.64235, -39.69548, -39.74771, -39.79758, 
        -39.84684, -39.89451, -39.94107, -39.98693, -40.03245, -40.07799, 
        -40.12382, -40.16955, -40.21471, -40.25869, -40.30067, -40.34066, 
        -40.37871, -40.41496, -40.44911, -40.48359, -40.51778, -40.55176, 
        -40.58503, -40.61696, -40.6472, -40.67546, -40.70193, -40.72693, 
        -40.75039, -40.77201, -40.79209, -40.81054, -40.8277, -40.84311, 
        -40.85902, -40.87495, -40.89117, -40.9076, -40.92387, -40.93979, 
        -40.95583, -40.97154, -40.98792, -41.0042, -41.02034, -41.03636, 
        -41.05157, -41.06614, -41.08059, -41.09411, -41.10959, -41.12586, 
        -41.14256, -41.15899, -41.17403, -41.18738, -41.19928, -41.21061, 
        -41.22228, -41.2341, -41.24633, -41.25884, -41.27119, -41.28321, 
        -41.2951, -41.30577, -41.31745, -41.32944, -41.34226, -41.35583, 
        -41.37057, -41.38684, -41.40459, -41.4237, -41.44342, -41.46341, 
        -41.48357, -41.50376, -41.52431, -41.54543, -41.56665, -41.58765, 
        -41.60788, -41.6261, -41.64449, -41.66272, -41.682, -41.70235, 
        -41.72412, -41.74666, -41.76949, -41.79181, -41.81348, -41.83466, 
        -41.85579, -41.87696, -41.89835, -41.91973, -41.94155, -41.96368, 
        -41.98613, -42.00786, -42.03066, -42.05342, -42.07556, -42.09623, 
        -42.11481, -42.13034, -42.14353, -42.15511, -42.16597, -42.17638, 
        -42.18658, -42.19665, -42.20651, -42.21593, -42.22429, -42.2313, 
        -42.23677, -42.24107, -42.24446, -42.24619, -42.24831, -42.24989, 
        -42.25154, -42.25315, -42.25607, -42.26058, -42.2671, -42.27527, 
        -42.28476, -42.29549, -42.30751, -42.3205, -42.33429, -42.34864, 
        -42.36345, -42.37821, -42.39314, -42.40799, -42.42312, -42.43842, 
        -42.45279, -42.46804, -42.48358, -42.4994, -42.51516, -42.53025, 
        -42.54441, -42.5573, -42.56953, -42.58161, -42.59436, -42.60786, 
        -42.62149, -42.63484, -42.64702, -42.65822, -42.66864, -42.67901, 
        -42.68977, -42.70146, -42.71471, -42.72993, -42.74741, -42.76572, 
        -42.78622, -42.80708, -42.82737, -42.84687, -42.86472, -42.88062, 
        -42.89464, -42.90729, -42.91897, -42.93, -42.94059, -42.95142, 
        -42.96225, -42.97371, -42.98555, -42.99751, -43.00907, -43.01994, 
        -43.02991, -43.03902, -43.04732, -43.05469, -43.06065, -43.06509, 
        -43.06721, -43.06871, -43.0684, -43.06651, -43.06297, -43.05789, 
        -43.05206, -43.04579, -43.03965, -43.03364, -43.02801, -43.02306, 
        -43.0182, -43.01337, -43.00792, -43.00221, -42.99598, -42.98955, 
        -42.98292, -42.97609, -42.96907, -42.96177, -42.9543, -42.94623, 
        -42.9375, -42.92844, -42.91964, -42.91172, -42.90357, -42.8975, 
        -42.89288, -42.88967, -42.88811, -42.88867, -42.89122, -42.8953, 
        -42.90094, -42.90743, -42.91439, -42.92122, -42.92781, -42.93365, 
        -42.93869, -42.94288, -42.94621, -42.94921, -42.95236, -42.95543, 
        -42.95847, -42.96185, -42.9654, -42.96865, -42.9718, -42.97432, 
        -42.9762, -42.97713, -42.97788, -42.97758, -42.9775, -42.97634, 
        -42.97419, -42.97134, -42.96645, -42.96144, -42.95559, -42.94879, 
        -42.94109, -42.93261, -42.92414, -42.91598, -42.90878, -42.90317, 
        -42.89927, -42.89651, -42.89481, -42.89345, -42.8918, -42.88953, 
        -42.88559, -42.87994, -42.87236, -42.86315, -42.85229, -42.83904, 
        -42.82298, -42.80317, -42.77853, -42.74823, -42.71194, -42.66908, 
        -42.62018, -42.56527, -42.50429, -42.43682, -42.36216, -42.27938, 
        -42.18699, -42.08416, -41.97043, -41.84637, -41.71472, -41.57888, 
        -41.44276, -41.31044, -41.18468, -41.068, -40.96186, -40.86509, 
        -40.77858,
  -39.39111, -39.44108, -39.49267, -39.54468, -39.59604, -39.64625, 
        -39.69531, -39.74313, -39.78978, -39.83584, -39.88134, -39.92664, 
        -39.97199, -40.01719, -40.0617, -40.10394, -40.14551, -40.18517, 
        -40.22316, -40.25964, -40.29517, -40.33024, -40.36502, -40.39948, 
        -40.4332, -40.46561, -40.49624, -40.52491, -40.55167, -40.57658, 
        -40.59882, -40.62023, -40.64008, -40.65847, -40.6757, -40.69234, 
        -40.70885, -40.72567, -40.74272, -40.76002, -40.77733, -40.79457, 
        -40.81149, -40.82859, -40.84587, -40.86335, -40.87961, -40.89653, 
        -40.91288, -40.9287, -40.94425, -40.96001, -40.9763, -40.99321, 
        -41.0107, -41.02791, -41.04393, -41.0584, -41.07161, -41.08426, 
        -41.09676, -41.1096, -41.12159, -41.13464, -41.14776, -41.16075, 
        -41.17353, -41.18592, -41.19835, -41.21111, -41.2245, -41.23921, 
        -41.25522, -41.27279, -41.29173, -41.31143, -41.33146, -41.35204, 
        -41.37288, -41.39299, -41.41488, -41.43725, -41.45971, -41.48167, 
        -41.50274, -41.5228, -41.54209, -41.56107, -41.58074, -41.60167, 
        -41.62414, -41.64726, -41.67085, -41.69348, -41.71553, -41.73674, 
        -41.75773, -41.77784, -41.7992, -41.82082, -41.84255, -41.86465, 
        -41.88724, -41.90979, -41.93226, -41.9549, -41.97691, -41.99797, 
        -42.01716, -42.03346, -42.04695, -42.05841, -42.06908, -42.07904, 
        -42.08847, -42.0975, -42.10504, -42.11305, -42.12016, -42.12627, 
        -42.13096, -42.13458, -42.13726, -42.13931, -42.14091, -42.14232, 
        -42.1438, -42.14589, -42.14879, -42.15341, -42.15993, -42.16809, 
        -42.1778, -42.18881, -42.20093, -42.21392, -42.22754, -42.24038, 
        -42.25435, -42.26815, -42.28201, -42.29629, -42.31089, -42.32581, 
        -42.34082, -42.35616, -42.3716, -42.3873, -42.40269, -42.41749, 
        -42.43097, -42.44326, -42.45497, -42.46679, -42.47953, -42.49282, 
        -42.50637, -42.51971, -42.53206, -42.54234, -42.55285, -42.56316, 
        -42.5738, -42.58529, -42.59839, -42.61338, -42.63075, -42.65025, 
        -42.6713, -42.69299, -42.71457, -42.73515, -42.75429, -42.77166, 
        -42.7873, -42.80149, -42.81461, -42.82713, -42.83939, -42.85179, 
        -42.86454, -42.87797, -42.89154, -42.90411, -42.91708, -42.92929, 
        -42.94048, -42.95073, -42.96009, -42.96862, -42.97607, -42.98233, 
        -42.98717, -42.9902, -42.99145, -42.99072, -42.98811, -42.98426, 
        -42.97948, -42.97464, -42.96965, -42.96519, -42.96099, -42.95712, 
        -42.95327, -42.94883, -42.944, -42.93872, -42.933, -42.92675, 
        -42.91914, -42.91255, -42.90561, -42.89857, -42.89103, -42.88296, 
        -42.87429, -42.86551, -42.85749, -42.85007, -42.84389, -42.83894, 
        -42.83528, -42.83302, -42.83233, -42.83385, -42.83705, -42.84191, 
        -42.84812, -42.85539, -42.86312, -42.87102, -42.87852, -42.88524, 
        -42.89082, -42.89518, -42.89858, -42.90168, -42.90502, -42.90818, 
        -42.91175, -42.91548, -42.91845, -42.9225, -42.92633, -42.92954, 
        -42.93185, -42.93357, -42.93471, -42.93541, -42.93526, -42.93419, 
        -42.93144, -42.92825, -42.92413, -42.91913, -42.91338, -42.90685, 
        -42.89952, -42.89125, -42.8829, -42.87484, -42.86798, -42.86211, 
        -42.85779, -42.85472, -42.85244, -42.85095, -42.84947, -42.84747, 
        -42.84415, -42.83891, -42.83186, -42.82277, -42.81153, -42.79794, 
        -42.78127, -42.76095, -42.73607, -42.70566, -42.66945, -42.62695, 
        -42.57732, -42.52299, -42.46257, -42.39635, -42.32348, -42.24272, 
        -42.153, -42.05343, -41.94359, -41.82391, -41.69692, -41.56595, 
        -41.43473, -41.3068, -41.18532, -41.07195, -40.96825, -40.87412, 
        -40.78851,
  -39.24218, -39.29234, -39.3429, -39.39364, -39.44401, -39.49337, 
        -39.54174, -39.58891, -39.63534, -39.68116, -39.72557, -39.77078, 
        -39.8159, -39.86077, -39.90488, -39.94767, -39.9888, -40.02829, 
        -40.06627, -40.10299, -40.13895, -40.17459, -40.20991, -40.24503, 
        -40.27928, -40.31128, -40.34237, -40.37139, -40.39808, -40.42282, 
        -40.44547, -40.46645, -40.48593, -40.50431, -40.52167, -40.53864, 
        -40.55577, -40.57337, -40.59131, -40.60969, -40.62733, -40.64565, 
        -40.66403, -40.68227, -40.70077, -40.71936, -40.73774, -40.75594, 
        -40.77355, -40.79082, -40.80762, -40.8246, -40.84188, -40.85949, 
        -40.8774, -40.89512, -40.91092, -40.92623, -40.94057, -40.9542, 
        -40.96785, -40.98163, -40.99554, -41.0094, -41.02337, -41.03748, 
        -41.05144, -41.06491, -41.0784, -41.09213, -41.10665, -41.12254, 
        -41.13986, -41.15748, -41.17722, -41.19779, -41.21844, -41.23927, 
        -41.26058, -41.28274, -41.30561, -41.32903, -41.3526, -41.37547, 
        -41.3972, -41.41788, -41.43793, -41.45809, -41.47866, -41.50012, 
        -41.52308, -41.54591, -41.56989, -41.59299, -41.61518, -41.63661, 
        -41.65756, -41.67847, -41.69984, -41.72137, -41.74327, -41.76548, 
        -41.78787, -41.81057, -41.83289, -41.855, -41.87682, -41.89785, 
        -41.91728, -41.93423, -41.94765, -41.95942, -41.96981, -41.97923, 
        -41.98812, -41.99635, -42.00379, -42.01056, -42.01667, -42.02198, 
        -42.02605, -42.02885, -42.0309, -42.03246, -42.03377, -42.03515, 
        -42.03668, -42.03915, -42.04252, -42.04742, -42.05319, -42.06143, 
        -42.07126, -42.08245, -42.09465, -42.10748, -42.12083, -42.134, 
        -42.14711, -42.16001, -42.17313, -42.18668, -42.20081, -42.21548, 
        -42.23047, -42.24558, -42.26083, -42.27617, -42.29107, -42.30511, 
        -42.31788, -42.32853, -42.33976, -42.35118, -42.36337, -42.3765, 
        -42.38976, -42.40292, -42.41539, -42.42679, -42.43726, -42.4476, 
        -42.45823, -42.46989, -42.4829, -42.49797, -42.51545, -42.53537, 
        -42.55703, -42.57951, -42.60214, -42.62406, -42.6445, -42.66317, 
        -42.67987, -42.69428, -42.70872, -42.72265, -42.73638, -42.75034, 
        -42.76473, -42.77996, -42.79544, -42.81058, -42.82518, -42.83873, 
        -42.85112, -42.8625, -42.87268, -42.88229, -42.8912, -42.89902, 
        -42.90546, -42.91007, -42.91258, -42.91305, -42.91146, -42.90873, 
        -42.90534, -42.9017, -42.89815, -42.89423, -42.8914, -42.88868, 
        -42.88561, -42.88218, -42.87802, -42.87353, -42.86827, -42.86218, 
        -42.85583, -42.84923, -42.84224, -42.83498, -42.82734, -42.81911, 
        -42.81086, -42.80276, -42.79524, -42.78884, -42.78353, -42.77964, 
        -42.77686, -42.77533, -42.77576, -42.77783, -42.78176, -42.78742, 
        -42.79441, -42.80212, -42.81057, -42.818, -42.82588, -42.83311, 
        -42.83876, -42.84315, -42.84675, -42.85004, -42.85343, -42.85732, 
        -42.86169, -42.86658, -42.87129, -42.87588, -42.87997, -42.88339, 
        -42.88632, -42.88876, -42.89054, -42.8914, -42.89148, -42.89021, 
        -42.88788, -42.88475, -42.88063, -42.87573, -42.87011, -42.86377, 
        -42.85692, -42.84909, -42.84101, -42.83337, -42.82625, -42.82026, 
        -42.8154, -42.81171, -42.80906, -42.80728, -42.80484, -42.80312, 
        -42.8003, -42.79583, -42.78921, -42.78042, -42.76915, -42.75521, 
        -42.73811, -42.71724, -42.69182, -42.66129, -42.62525, -42.58313, 
        -42.53526, -42.48154, -42.42192, -42.35655, -42.28459, -42.20528, 
        -42.11764, -42.0206, -41.914, -41.79825, -41.6758, -41.5498, 
        -41.42366, -41.30079, -41.18381, -41.07481, -40.97437, -40.88251, 
        -40.79791,
  -39.09349, -39.14294, -39.19267, -39.24231, -39.29141, -39.33858, 
        -39.38581, -39.43214, -39.47787, -39.52314, -39.56833, -39.61331, 
        -39.65823, -39.70294, -39.74683, -39.78942, -39.83043, -39.86982, 
        -39.90771, -39.94467, -39.97998, -40.01603, -40.05193, -40.08751, 
        -40.12234, -40.15571, -40.18724, -40.21622, -40.24294, -40.26714, 
        -40.28913, -40.30967, -40.32883, -40.34706, -40.3647, -40.38126, 
        -40.39919, -40.41771, -40.43697, -40.45675, -40.47658, -40.49631, 
        -40.51591, -40.53536, -40.55491, -40.57457, -40.59418, -40.61361, 
        -40.63292, -40.65156, -40.67006, -40.68728, -40.70538, -40.72369, 
        -40.74211, -40.7601, -40.7775, -40.79366, -40.80886, -40.8237, 
        -40.83847, -40.85319, -40.8679, -40.8827, -40.89771, -40.91292, 
        -40.92795, -40.94193, -40.95664, -40.97184, -40.98751, -41.00468, 
        -41.02288, -41.04259, -41.06312, -41.08431, -41.10566, -41.12732, 
        -41.1492, -41.17219, -41.19601, -41.22041, -41.24474, -41.26838, 
        -41.29092, -41.31124, -41.332, -41.35287, -41.37458, -41.39689, 
        -41.42029, -41.44455, -41.46902, -41.49243, -41.51484, -41.53645, 
        -41.55768, -41.57878, -41.60013, -41.62171, -41.64377, -41.66629, 
        -41.68856, -41.71004, -41.73216, -41.75367, -41.77505, -41.79579, 
        -41.81527, -41.83263, -41.84749, -41.86012, -41.8707, -41.87983, 
        -41.88778, -41.89496, -41.90148, -41.90743, -41.91282, -41.9174, 
        -41.92068, -41.92297, -41.9244, -41.92459, -41.9257, -41.92715, 
        -41.929, -41.93167, -41.93562, -41.94109, -41.94812, -41.95659, 
        -41.96658, -41.9775, -41.98967, -42.00235, -42.0152, -42.02778, 
        -42.04021, -42.05241, -42.06495, -42.07792, -42.09158, -42.10602, 
        -42.1199, -42.13495, -42.1501, -42.1649, -42.17923, -42.19251, 
        -42.20444, -42.21541, -42.22611, -42.23714, -42.24888, -42.26135, 
        -42.27451, -42.28748, -42.29979, -42.3112, -42.322, -42.33245, 
        -42.34328, -42.35501, -42.3684, -42.38383, -42.40167, -42.42108, 
        -42.44331, -42.46677, -42.49041, -42.51352, -42.53497, -42.55463, 
        -42.57233, -42.58875, -42.60415, -42.61902, -42.63392, -42.64926, 
        -42.66517, -42.68191, -42.69905, -42.716, -42.73212, -42.74706, 
        -42.76063, -42.7729, -42.78415, -42.79483, -42.80491, -42.81434, 
        -42.82104, -42.827, -42.83072, -42.83213, -42.83212, -42.83059, 
        -42.82845, -42.82611, -42.82418, -42.82257, -42.82102, -42.81945, 
        -42.81767, -42.81503, -42.812, -42.80804, -42.80346, -42.79793, 
        -42.79171, -42.78507, -42.77794, -42.77029, -42.76259, -42.75446, 
        -42.74663, -42.73914, -42.73236, -42.72668, -42.72121, -42.71779, 
        -42.71588, -42.71531, -42.71666, -42.71959, -42.72462, -42.73084, 
        -42.73841, -42.74654, -42.75538, -42.76405, -42.77213, -42.77912, 
        -42.78473, -42.78913, -42.79289, -42.79666, -42.80059, -42.80552, 
        -42.81077, -42.8165, -42.82185, -42.82684, -42.83133, -42.83533, 
        -42.83875, -42.84148, -42.84355, -42.84491, -42.84519, -42.84449, 
        -42.84253, -42.83966, -42.83492, -42.83034, -42.8251, -42.81909, 
        -42.81239, -42.80511, -42.79752, -42.78984, -42.78285, -42.77647, 
        -42.77097, -42.76654, -42.76329, -42.76104, -42.75949, -42.75795, 
        -42.75562, -42.75159, -42.74557, -42.73725, -42.72623, -42.7123, 
        -42.69497, -42.67364, -42.64791, -42.61746, -42.58158, -42.54033, 
        -42.49323, -42.44043, -42.38166, -42.31702, -42.24561, -42.16718, 
        -42.08079, -41.98589, -41.88199, -41.7699, -41.65173, -41.53051, 
        -41.4096, -41.29147, -41.1792, -41.07415, -40.97716, -40.88704, 
        -40.80465,
  -38.94424, -38.99235, -39.04131, -39.08977, -39.13765, -39.18436, 
        -39.2301, -39.27508, -39.31976, -39.36456, -39.40932, -39.45416, 
        -39.49901, -39.54361, -39.58739, -39.62894, -39.66992, -39.70927, 
        -39.74717, -39.78413, -39.82058, -39.85691, -39.89318, -39.92915, 
        -39.96428, -39.99802, -40.02964, -40.05869, -40.08482, -40.10833, 
        -40.12864, -40.14875, -40.16784, -40.18618, -40.20427, -40.22251, 
        -40.24142, -40.26139, -40.28202, -40.30323, -40.32463, -40.34589, 
        -40.36677, -40.38741, -40.40798, -40.42874, -40.44851, -40.46925, 
        -40.49007, -40.51077, -40.53069, -40.55021, -40.56918, -40.58818, 
        -40.60691, -40.62531, -40.64316, -40.66005, -40.67624, -40.69207, 
        -40.70793, -40.72359, -40.73819, -40.75393, -40.76996, -40.78608, 
        -40.80249, -40.81882, -40.83535, -40.85205, -40.86954, -40.88745, 
        -40.90675, -40.92723, -40.94843, -40.96988, -40.99192, -41.01438, 
        -41.03763, -41.06046, -41.08525, -41.1106, -41.13556, -41.1596, 
        -41.18262, -41.20454, -41.22596, -41.24752, -41.27003, -41.29327, 
        -41.31726, -41.34208, -41.36657, -41.39031, -41.41339, -41.43555, 
        -41.45713, -41.47765, -41.49926, -41.52108, -41.54345, -41.56617, 
        -41.58887, -41.61125, -41.63309, -41.65425, -41.67484, -41.69507, 
        -41.71412, -41.73141, -41.74687, -41.76012, -41.77112, -41.77985, 
        -41.78716, -41.7936, -41.79817, -41.80322, -41.80781, -41.8115, 
        -41.81424, -41.81592, -41.81695, -41.81776, -41.81869, -41.82004, 
        -41.82224, -41.82538, -41.82973, -41.83563, -41.84302, -41.85163, 
        -41.86165, -41.87263, -41.8843, -41.89661, -41.90929, -41.92038, 
        -41.93233, -41.94416, -41.95621, -41.96889, -41.9823, -41.99647, 
        -42.01128, -42.0263, -42.04112, -42.0556, -42.06916, -42.08154, 
        -42.09289, -42.1035, -42.11388, -42.12476, -42.13618, -42.14816, 
        -42.16083, -42.17327, -42.18551, -42.19613, -42.20714, -42.21817, 
        -42.22946, -42.24176, -42.2554, -42.27129, -42.28947, -42.31041, 
        -42.33332, -42.35756, -42.38205, -42.40589, -42.4282, -42.44845, 
        -42.4668, -42.48391, -42.5001, -42.51579, -42.5315, -42.54794, 
        -42.56501, -42.58317, -42.60177, -42.61916, -42.63674, -42.65291, 
        -42.66731, -42.68068, -42.69304, -42.70474, -42.71608, -42.72671, 
        -42.73551, -42.74277, -42.74727, -42.74998, -42.75111, -42.75103, 
        -42.75029, -42.74969, -42.74931, -42.74924, -42.74912, -42.74875, 
        -42.74801, -42.7465, -42.74411, -42.74106, -42.73706, -42.73218, 
        -42.72527, -42.71861, -42.7111, -42.70331, -42.69576, -42.68816, 
        -42.68098, -42.67413, -42.66804, -42.66282, -42.65847, -42.65548, 
        -42.65409, -42.65444, -42.65681, -42.66105, -42.66695, -42.67408, 
        -42.68208, -42.69056, -42.69961, -42.70829, -42.71611, -42.72275, 
        -42.7284, -42.73307, -42.737, -42.74097, -42.74578, -42.75146, 
        -42.75756, -42.76371, -42.76855, -42.77402, -42.77905, -42.78382, 
        -42.78723, -42.79051, -42.79274, -42.79425, -42.79539, -42.79537, 
        -42.79443, -42.79225, -42.789, -42.78503, -42.78034, -42.77475, 
        -42.76852, -42.76166, -42.75433, -42.74682, -42.73954, -42.73258, 
        -42.72628, -42.72083, -42.71696, -42.71439, -42.71268, -42.71119, 
        -42.70899, -42.7056, -42.70014, -42.69247, -42.6818, -42.66809, 
        -42.6507, -42.62922, -42.60338, -42.57302, -42.53773, -42.49717, 
        -42.45026, -42.39851, -42.34091, -42.27689, -42.20605, -42.12838, 
        -42.04304, -41.94989, -41.84863, -41.73993, -41.62578, -41.50878, 
        -41.39219, -41.27836, -41.17005, -41.06907, -40.97566, -40.88917, 
        -40.80938,
  -38.79336, -38.84224, -38.89047, -38.93779, -38.98422, -39.02948, 
        -39.07386, -39.11764, -39.16135, -39.20522, -39.24854, -39.29309, 
        -39.33781, -39.38232, -39.42617, -39.46867, -39.50968, -39.54905, 
        -39.58698, -39.6239, -39.66034, -39.69662, -39.73286, -39.76887, 
        -39.80404, -39.83673, -39.86829, -39.89687, -39.92247, -39.94554, 
        -39.96666, -39.98665, -40.00572, -40.02447, -40.04325, -40.06245, 
        -40.08263, -40.10389, -40.12629, -40.14913, -40.17109, -40.1937, 
        -40.21575, -40.23751, -40.25893, -40.28036, -40.30233, -40.32467, 
        -40.34716, -40.3696, -40.39118, -40.41199, -40.43216, -40.45187, 
        -40.47112, -40.49003, -40.5073, -40.52466, -40.54178, -40.5588, 
        -40.57577, -40.5924, -40.60892, -40.62554, -40.64257, -40.65995, 
        -40.67757, -40.69546, -40.71341, -40.73148, -40.75005, -40.76926, 
        -40.7893, -40.80934, -40.83105, -40.85334, -40.87621, -40.8997, 
        -40.92414, -40.94926, -40.97491, -41.00088, -41.02652, -41.05096, 
        -41.0745, -41.09694, -41.11919, -41.1415, -41.16437, -41.18816, 
        -41.21264, -41.23679, -41.26202, -41.28653, -41.31028, -41.33307, 
        -41.35534, -41.37725, -41.39932, -41.42154, -41.44438, -41.46744, 
        -41.49037, -41.51288, -41.53477, -41.55569, -41.57605, -41.59561, 
        -41.61404, -41.6311, -41.64544, -41.6588, -41.67002, -41.67902, 
        -41.68578, -41.69148, -41.69624, -41.70022, -41.70396, -41.7069, 
        -41.70886, -41.71001, -41.7106, -41.71131, -41.71215, -41.71364, 
        -41.71598, -41.71945, -41.72429, -41.73042, -41.73699, -41.74561, 
        -41.75544, -41.76631, -41.77787, -41.78981, -41.80196, -41.81421, 
        -41.82597, -41.83759, -41.8493, -41.86181, -41.87482, -41.88888, 
        -41.90361, -41.91833, -41.93292, -41.94682, -41.95982, -41.97186, 
        -41.98283, -41.99211, -42.00249, -42.0132, -42.02426, -42.03598, 
        -42.04821, -42.06041, -42.0727, -42.08477, -42.09636, -42.10785, 
        -42.11991, -42.13261, -42.14685, -42.16306, -42.18179, -42.20313, 
        -42.22658, -42.25134, -42.27635, -42.30038, -42.32289, -42.34363, 
        -42.36236, -42.37889, -42.39536, -42.41195, -42.42829, -42.44574, 
        -42.46386, -42.48292, -42.50259, -42.52204, -42.5404, -42.55747, 
        -42.57311, -42.58758, -42.60148, -42.61457, -42.62695, -42.63863, 
        -42.64867, -42.65675, -42.66255, -42.66649, -42.66873, -42.66992, 
        -42.67072, -42.67151, -42.6726, -42.67301, -42.67434, -42.6752, 
        -42.67558, -42.67504, -42.67345, -42.67117, -42.66764, -42.66319, 
        -42.65759, -42.65105, -42.64368, -42.63635, -42.62914, -42.62202, 
        -42.61565, -42.60958, -42.60374, -42.59857, -42.59421, -42.59154, 
        -42.5908, -42.59212, -42.59573, -42.60099, -42.6081, -42.61606, 
        -42.6245, -42.63338, -42.64241, -42.64964, -42.65711, -42.6638, 
        -42.66954, -42.6744, -42.67876, -42.6834, -42.68873, -42.69478, 
        -42.70099, -42.70741, -42.7136, -42.71967, -42.72537, -42.73012, 
        -42.73434, -42.73801, -42.74092, -42.74288, -42.74432, -42.74544, 
        -42.74534, -42.74387, -42.74181, -42.73869, -42.73461, -42.72967, 
        -42.72373, -42.71724, -42.71027, -42.70271, -42.69493, -42.68727, 
        -42.68016, -42.67406, -42.66953, -42.66652, -42.66344, -42.66187, 
        -42.65986, -42.65669, -42.65168, -42.6444, -42.63427, -42.62083, 
        -42.60381, -42.58267, -42.5571, -42.52735, -42.49288, -42.45329, 
        -42.40807, -42.35735, -42.30049, -42.23761, -42.16798, -42.09139, 
        -42.00742, -41.91612, -41.81727, -41.71169, -41.60107, -41.4878, 
        -41.37493, -41.26487, -41.15973, -41.06205, -40.9714, -40.88742, 
        -40.81019,
  -38.64285, -38.6912, -38.73866, -38.78492, -38.83001, -38.87303, 
        -38.91625, -38.9591, -39.00199, -39.04533, -39.08934, -39.13351, 
        -39.17799, -39.22212, -39.2656, -39.30803, -39.34903, -39.38845, 
        -39.42646, -39.46335, -39.49856, -39.53456, -39.57046, -39.606, 
        -39.64085, -39.67423, -39.70545, -39.73395, -39.75957, -39.78247, 
        -39.8034, -39.82346, -39.84282, -39.86211, -39.88148, -39.90082, 
        -39.9224, -39.94527, -39.96925, -39.99389, -40.01828, -40.04239, 
        -40.06561, -40.08786, -40.11016, -40.13277, -40.15597, -40.17975, 
        -40.2038, -40.22773, -40.25087, -40.27205, -40.29343, -40.31393, 
        -40.33365, -40.35283, -40.37166, -40.38992, -40.40786, -40.42575, 
        -40.44358, -40.46168, -40.47921, -40.49679, -40.51475, -40.53322, 
        -40.55216, -40.57117, -40.58952, -40.60886, -40.62844, -40.64873, 
        -40.66964, -40.69151, -40.71394, -40.73693, -40.76078, -40.78541, 
        -40.81094, -40.83729, -40.86403, -40.89043, -40.91602, -40.94107, 
        -40.9649, -40.98712, -41.01002, -41.03327, -41.05695, -41.08096, 
        -41.10593, -41.13148, -41.15726, -41.18272, -41.20747, -41.23121, 
        -41.25413, -41.27662, -41.29903, -41.3218, -41.34512, -41.36842, 
        -41.392, -41.41399, -41.4363, -41.45755, -41.47754, -41.49665, 
        -41.51459, -41.53088, -41.54573, -41.55881, -41.56977, -41.57874, 
        -41.58558, -41.59084, -41.59466, -41.59763, -41.60049, -41.60263, 
        -41.60421, -41.6049, -41.60529, -41.60476, -41.60544, -41.60715, 
        -41.60954, -41.61346, -41.6186, -41.62479, -41.63219, -41.64069, 
        -41.65033, -41.66087, -41.6721, -41.68397, -41.69614, -41.70825, 
        -41.72004, -41.73174, -41.74351, -41.75563, -41.76852, -41.78221, 
        -41.79556, -41.81025, -41.82454, -41.8382, -41.85089, -41.86255, 
        -41.87341, -41.88379, -41.89407, -41.90474, -41.9159, -41.92767, 
        -41.93987, -41.95225, -41.96471, -41.97728, -41.98979, -42.00196, 
        -42.01444, -42.02777, -42.04241, -42.05914, -42.07826, -42.09886, 
        -42.12248, -42.14713, -42.17208, -42.19632, -42.21882, -42.23936, 
        -42.25835, -42.27594, -42.29303, -42.30985, -42.32704, -42.34527, 
        -42.36433, -42.38423, -42.40418, -42.42389, -42.44274, -42.46039, 
        -42.47713, -42.49301, -42.50838, -42.52304, -42.53686, -42.54958, 
        -42.55962, -42.56882, -42.57576, -42.58072, -42.58405, -42.58665, 
        -42.58892, -42.59124, -42.59369, -42.59636, -42.59893, -42.60115, 
        -42.60266, -42.60305, -42.60209, -42.59999, -42.59685, -42.59254, 
        -42.58721, -42.58094, -42.57444, -42.56774, -42.56134, -42.55539, 
        -42.54965, -42.54399, -42.53816, -42.53282, -42.52861, -42.52494, 
        -42.52486, -42.52705, -42.53185, -42.53844, -42.54657, -42.55552, 
        -42.56465, -42.57378, -42.58257, -42.5907, -42.59806, -42.60478, 
        -42.61053, -42.61575, -42.62079, -42.62596, -42.63169, -42.6377, 
        -42.64388, -42.64993, -42.6566, -42.66292, -42.66862, -42.67382, 
        -42.67839, -42.68272, -42.68649, -42.68942, -42.69238, -42.69411, 
        -42.69483, -42.69468, -42.69321, -42.69012, -42.6867, -42.68225, 
        -42.67716, -42.67082, -42.66397, -42.65622, -42.64797, -42.63974, 
        -42.63195, -42.62529, -42.62043, -42.61701, -42.61461, -42.61272, 
        -42.61053, -42.60734, -42.6026, -42.59567, -42.58585, -42.57291, 
        -42.55616, -42.53555, -42.51083, -42.48185, -42.44828, -42.40948, 
        -42.36521, -42.31557, -42.25986, -42.19829, -42.13026, -42.05521, 
        -41.9732, -41.88414, -41.78794, -41.68524, -41.57779, -41.46785, 
        -41.3579, -41.25054, -41.14753, -41.0518, -40.96383, -40.88122, 
        -40.80591,
  -38.49075, -38.53743, -38.58385, -38.629, -38.67321, -38.71659, 
        -38.75922, -38.80171, -38.84441, -38.88752, -38.93113, -38.97517, 
        -39.01904, -39.06255, -39.10539, -39.14637, -39.18717, -39.22658, 
        -39.26459, -39.30146, -39.33759, -39.37327, -39.40851, -39.44339, 
        -39.47756, -39.51031, -39.54129, -39.56985, -39.59566, -39.61876, 
        -39.63906, -39.6594, -39.67912, -39.69881, -39.7192, -39.74064, 
        -39.76355, -39.78794, -39.81358, -39.83979, -39.86565, -39.89086, 
        -39.91486, -39.93819, -39.96151, -39.98534, -40.00868, -40.03384, 
        -40.0593, -40.08456, -40.10915, -40.13259, -40.15502, -40.17628, 
        -40.19672, -40.2163, -40.23563, -40.25442, -40.27334, -40.29239, 
        -40.31128, -40.33019, -40.34795, -40.36697, -40.38591, -40.40531, 
        -40.42524, -40.44521, -40.46539, -40.48581, -40.5067, -40.52815, 
        -40.55027, -40.57322, -40.59667, -40.62071, -40.6452, -40.67081, 
        -40.69722, -40.72328, -40.75073, -40.77779, -40.80378, -40.8289, 
        -40.8532, -40.87713, -40.901, -40.92507, -40.94965, -40.97454, 
        -40.99981, -41.02563, -41.05167, -41.07788, -41.10358, -41.12846, 
        -41.15232, -41.17448, -41.19733, -41.22059, -41.24446, -41.26836, 
        -41.29263, -41.31631, -41.3393, -41.36096, -41.3809, -41.39993, 
        -41.41734, -41.43278, -41.44698, -41.45936, -41.46967, -41.47857, 
        -41.48514, -41.49038, -41.49266, -41.49484, -41.49669, -41.49805, 
        -41.49914, -41.49981, -41.49995, -41.50041, -41.50128, -41.50282, 
        -41.50566, -41.50974, -41.51471, -41.52103, -41.52822, -41.53654, 
        -41.54572, -41.55585, -41.5668, -41.57829, -41.59051, -41.60191, 
        -41.61414, -41.62619, -41.63788, -41.64969, -41.66228, -41.67573, 
        -41.68972, -41.704, -41.71821, -41.73172, -41.74419, -41.75571, 
        -41.76656, -41.77712, -41.78777, -41.79882, -41.81047, -41.82241, 
        -41.83475, -41.84768, -41.86097, -41.87337, -41.88642, -41.89946, 
        -41.91254, -41.92639, -41.94147, -41.95845, -41.97782, -41.99935, 
        -42.02277, -42.04708, -42.07167, -42.0953, -42.11761, -42.13806, 
        -42.15702, -42.17484, -42.19202, -42.20932, -42.22714, -42.246, 
        -42.26549, -42.28575, -42.30571, -42.32436, -42.34296, -42.36112, 
        -42.37896, -42.39633, -42.41357, -42.43003, -42.4455, -42.45951, 
        -42.47178, -42.48169, -42.48946, -42.49546, -42.50012, -42.50409, 
        -42.50775, -42.51143, -42.51503, -42.51904, -42.52279, -42.52606, 
        -42.5284, -42.52917, -42.52851, -42.52653, -42.52364, -42.51964, 
        -42.51475, -42.50811, -42.50254, -42.49658, -42.49125, -42.48625, 
        -42.48121, -42.47606, -42.47044, -42.46512, -42.46094, -42.45866, 
        -42.45884, -42.46181, -42.46764, -42.47553, -42.48473, -42.49443, 
        -42.50434, -42.51394, -42.52267, -42.53091, -42.53839, -42.54495, 
        -42.55089, -42.5565, -42.56187, -42.56728, -42.57297, -42.57883, 
        -42.58476, -42.59097, -42.59655, -42.60289, -42.6087, -42.61428, 
        -42.61946, -42.62431, -42.62909, -42.63332, -42.63698, -42.63954, 
        -42.64138, -42.64262, -42.64237, -42.64112, -42.63863, -42.63499, 
        -42.63041, -42.62439, -42.61737, -42.60958, -42.60085, -42.59218, 
        -42.58419, -42.57744, -42.57237, -42.56867, -42.56583, -42.56341, 
        -42.56083, -42.55736, -42.55255, -42.54575, -42.53627, -42.52367, 
        -42.50762, -42.48769, -42.46386, -42.4358, -42.4032, -42.36523, 
        -42.32101, -42.27192, -42.21755, -42.15754, -42.09144, -42.01894, 
        -41.93961, -41.85328, -41.76029, -41.66082, -41.55642, -41.44915, 
        -41.34134, -41.23573, -41.13483, -41.04025, -40.95244, -40.87236, 
        -40.7985,
  -38.33597, -38.38273, -38.42815, -38.47262, -38.51605, -38.55926, 
        -38.60195, -38.64465, -38.68758, -38.73071, -38.77344, -38.81671, 
        -38.85994, -38.90269, -38.94477, -38.98607, -39.02644, -39.06571, 
        -39.10378, -39.14071, -39.17679, -39.21216, -39.247, -39.28111, 
        -39.31434, -39.34573, -39.37631, -39.40474, -39.43079, -39.45433, 
        -39.47614, -39.49669, -39.51693, -39.53754, -39.55896, -39.58179, 
        -39.60594, -39.63179, -39.65892, -39.68645, -39.71251, -39.73852, 
        -39.76349, -39.78765, -39.81186, -39.83673, -39.86234, -39.8887, 
        -39.91552, -39.94217, -39.96818, -39.99292, -40.01626, -40.03853, 
        -40.05949, -40.0796, -40.09821, -40.11772, -40.13753, -40.15738, 
        -40.17735, -40.19714, -40.21715, -40.23725, -40.25754, -40.27804, 
        -40.29865, -40.31936, -40.3405, -40.36202, -40.38424, -40.40713, 
        -40.43075, -40.45392, -40.47859, -40.50344, -40.52877, -40.55493, 
        -40.58196, -40.60971, -40.63755, -40.66491, -40.69167, -40.71749, 
        -40.74215, -40.76671, -40.79153, -40.81651, -40.84173, -40.86727, 
        -40.89359, -40.91866, -40.9447, -40.97125, -40.99757, -41.02349, 
        -41.04852, -41.07283, -41.0966, -41.12036, -41.14465, -41.16902, 
        -41.19392, -41.21825, -41.2417, -41.26365, -41.28407, -41.3027, 
        -41.31981, -41.3349, -41.34747, -41.3593, -41.36945, -41.37749, 
        -41.38382, -41.38906, -41.3924, -41.39408, -41.39506, -41.39587, 
        -41.39634, -41.39664, -41.39703, -41.39721, -41.398, -41.39984, 
        -41.40265, -41.40669, -41.41198, -41.41788, -41.42396, -41.43182, 
        -41.44079, -41.4508, -41.46159, -41.47302, -41.48505, -41.49761, 
        -41.51015, -41.5225, -41.53431, -41.54622, -41.55843, -41.57147, 
        -41.58516, -41.59923, -41.61327, -41.62653, -41.63898, -41.65052, 
        -41.66161, -41.67144, -41.68264, -41.69434, -41.70652, -41.71889, 
        -41.73201, -41.74585, -41.75998, -41.77435, -41.78837, -41.80214, 
        -41.81577, -41.8299, -41.84544, -41.86271, -41.88192, -41.90338, 
        -41.92635, -41.95005, -41.97353, -41.99624, -42.01796, -42.03825, 
        -42.0572, -42.07431, -42.09211, -42.10983, -42.1279, -42.14691, 
        -42.16685, -42.18687, -42.20649, -42.22573, -42.24446, -42.26307, 
        -42.28173, -42.30088, -42.31994, -42.33826, -42.35564, -42.37114, 
        -42.38388, -42.39464, -42.40336, -42.41055, -42.41609, -42.4213, 
        -42.42635, -42.43166, -42.43655, -42.44066, -42.44533, -42.44947, 
        -42.45209, -42.45304, -42.4522, -42.45039, -42.44757, -42.44408, 
        -42.44009, -42.43571, -42.43088, -42.42599, -42.42137, -42.41703, 
        -42.41253, -42.40752, -42.40233, -42.39744, -42.39355, -42.39148, 
        -42.39206, -42.39561, -42.40216, -42.41096, -42.42122, -42.43215, 
        -42.44268, -42.45273, -42.46219, -42.46953, -42.47672, -42.48319, 
        -42.48937, -42.49545, -42.50117, -42.50677, -42.51226, -42.51771, 
        -42.52356, -42.52959, -42.53592, -42.54201, -42.54811, -42.55409, 
        -42.55997, -42.56564, -42.5713, -42.5765, -42.58142, -42.58534, 
        -42.58855, -42.5906, -42.59146, -42.59127, -42.58977, -42.58699, 
        -42.58278, -42.57714, -42.57029, -42.56223, -42.55347, -42.54473, 
        -42.53692, -42.53025, -42.52508, -42.52116, -42.51695, -42.51397, 
        -42.51085, -42.50687, -42.50199, -42.49519, -42.48583, -42.47324, 
        -42.45754, -42.4383, -42.41533, -42.38836, -42.3567, -42.31974, 
        -42.27724, -42.22915, -42.17635, -42.11821, -42.05461, -41.98483, 
        -41.90879, -41.82586, -41.73615, -41.64001, -41.53846, -41.4337, 
        -41.328, -41.22382, -41.12331, -41.02861, -40.94075, -40.86055, 
        -40.78682,
  -38.18027, -38.22598, -38.27055, -38.31425, -38.35758, -38.40083, 
        -38.44334, -38.4869, -38.53065, -38.57425, -38.61765, -38.66077, 
        -38.70342, -38.7452, -38.78609, -38.82649, -38.86626, -38.90528, 
        -38.94336, -38.98055, -39.01578, -39.05109, -39.08552, -39.11894, 
        -39.15143, -39.18283, -39.21285, -39.24109, -39.26749, -39.29154, 
        -39.31391, -39.33525, -39.35638, -39.3779, -39.40053, -39.4235, 
        -39.44911, -39.47628, -39.50475, -39.5334, -39.56149, -39.58842, 
        -39.61412, -39.63917, -39.66438, -39.69006, -39.71663, -39.74401, 
        -39.77187, -39.79974, -39.8268, -39.85163, -39.87606, -39.89916, 
        -39.92088, -39.94157, -39.96188, -39.98208, -40.00254, -40.02331, 
        -40.04414, -40.06491, -40.08597, -40.10717, -40.12876, -40.15034, 
        -40.17189, -40.19333, -40.21425, -40.23692, -40.26067, -40.28518, 
        -40.31046, -40.33601, -40.36169, -40.38746, -40.41341, -40.43999, 
        -40.4674, -40.49524, -40.52367, -40.55151, -40.57878, -40.60555, 
        -40.63174, -40.65636, -40.68174, -40.70755, -40.73343, -40.75961, 
        -40.78584, -40.81226, -40.83867, -40.86523, -40.89182, -40.91842, 
        -40.94431, -40.9698, -40.99472, -41.01933, -41.04387, -41.06874, 
        -41.09393, -41.11765, -41.14175, -41.16417, -41.18486, -41.20352, 
        -41.22035, -41.23534, -41.24866, -41.2601, -41.26973, -41.27778, 
        -41.28425, -41.28896, -41.29203, -41.29364, -41.29437, -41.29464, 
        -41.29488, -41.29511, -41.29535, -41.29495, -41.29588, -41.29772, 
        -41.30055, -41.30432, -41.30896, -41.31461, -41.32132, -41.32914, 
        -41.338, -41.34809, -41.35865, -41.37001, -41.38204, -41.39452, 
        -41.40724, -41.41986, -41.43202, -41.4439, -41.45609, -41.46878, 
        -41.48116, -41.49503, -41.50872, -41.52213, -41.5346, -41.54642, 
        -41.55796, -41.56937, -41.5811, -41.5934, -41.60621, -41.61921, 
        -41.63317, -41.64808, -41.66364, -41.67913, -41.69389, -41.70815, 
        -41.7223, -41.73693, -41.75277, -41.77023, -41.78955, -41.80952, 
        -41.83184, -41.85444, -41.87667, -41.89845, -41.91946, -41.93977, 
        -41.9588, -41.97733, -41.9953, -42.01335, -42.03197, -42.05135, 
        -42.07116, -42.0909, -42.11004, -42.12865, -42.14714, -42.1659, 
        -42.1859, -42.20652, -42.22757, -42.2479, -42.26658, -42.28319, 
        -42.29619, -42.30788, -42.31762, -42.32549, -42.33229, -42.33838, 
        -42.34476, -42.35119, -42.35746, -42.36355, -42.36898, -42.3733, 
        -42.3761, -42.3768, -42.37595, -42.37376, -42.37123, -42.36848, 
        -42.36537, -42.36198, -42.35839, -42.35484, -42.35108, -42.34717, 
        -42.34285, -42.33823, -42.3334, -42.3288, -42.32542, -42.32294, 
        -42.32398, -42.328, -42.33517, -42.34477, -42.35603, -42.36777, 
        -42.37931, -42.39008, -42.3998, -42.40788, -42.41519, -42.42166, 
        -42.42818, -42.43456, -42.4406, -42.44628, -42.45181, -42.45742, 
        -42.46294, -42.46852, -42.4744, -42.48045, -42.48654, -42.49283, 
        -42.49908, -42.50539, -42.51202, -42.51849, -42.52454, -42.52993, 
        -42.53454, -42.53789, -42.54011, -42.53994, -42.53948, -42.53753, 
        -42.53389, -42.52871, -42.52184, -42.51369, -42.50503, -42.4966, 
        -42.48911, -42.48277, -42.47789, -42.47361, -42.46999, -42.46645, 
        -42.46262, -42.45825, -42.453, -42.44614, -42.4369, -42.42451, 
        -42.40907, -42.39038, -42.36806, -42.3418, -42.31089, -42.27479, 
        -42.23309, -42.18621, -42.1347, -42.07893, -42.01796, -41.95172, 
        -41.87911, -41.7998, -41.71364, -41.62084, -41.52224, -41.41993, 
        -41.31607, -41.2127, -41.11223, -41.01656, -40.92727, -40.84446, 
        -40.76979,
  -38.0232, -38.06677, -38.11062, -38.15403, -38.19752, -38.24144, 
        -38.28595, -38.33042, -38.37458, -38.41868, -38.46235, -38.50507, 
        -38.54706, -38.58803, -38.62809, -38.66671, -38.70604, -38.74483, 
        -38.78294, -38.82032, -38.85666, -38.89202, -38.92622, -38.95919, 
        -38.99096, -39.02162, -39.05103, -39.07912, -39.10558, -39.12992, 
        -39.15195, -39.17406, -39.1961, -39.21891, -39.24289, -39.26831, 
        -39.29531, -39.32383, -39.35335, -39.38298, -39.41193, -39.43979, 
        -39.46632, -39.49238, -39.51845, -39.545, -39.57146, -39.59962, 
        -39.62821, -39.65722, -39.6851, -39.71181, -39.73709, -39.76101, 
        -39.78359, -39.80498, -39.82593, -39.84679, -39.86794, -39.88934, 
        -39.91081, -39.93247, -39.95337, -39.97574, -39.99828, -40.0208, 
        -40.04345, -40.06603, -40.08918, -40.11326, -40.13839, -40.16446, 
        -40.19138, -40.21821, -40.24483, -40.27142, -40.29778, -40.32498, 
        -40.35314, -40.3805, -40.40912, -40.43762, -40.46585, -40.49345, 
        -40.52048, -40.54727, -40.57395, -40.60013, -40.6264, -40.65252, 
        -40.67868, -40.70513, -40.73212, -40.75932, -40.78617, -40.81316, 
        -40.83979, -40.86484, -40.89044, -40.91561, -40.94071, -40.96577, 
        -40.99104, -41.01598, -41.04005, -41.06284, -41.08404, -41.10321, 
        -41.12033, -41.13538, -41.14876, -41.16025, -41.1699, -41.17789, 
        -41.18427, -41.18892, -41.19083, -41.19243, -41.19299, -41.19305, 
        -41.19323, -41.19353, -41.19414, -41.19487, -41.19608, -41.19793, 
        -41.20042, -41.20348, -41.20758, -41.2126, -41.21886, -41.22661, 
        -41.23573, -41.24593, -41.25657, -41.26788, -41.27986, -41.29148, 
        -41.30431, -41.31716, -41.32957, -41.34166, -41.35386, -41.3666, 
        -41.38004, -41.39389, -41.40766, -41.42094, -41.43361, -41.44587, 
        -41.4581, -41.4702, -41.48239, -41.49523, -41.50844, -41.52258, 
        -41.53759, -41.5536, -41.57038, -41.58577, -41.60131, -41.61633, 
        -41.63084, -41.6458, -41.66184, -41.6796, -41.69872, -41.71903, 
        -41.74012, -41.76147, -41.7826, -41.80342, -41.82396, -41.84406, 
        -41.86362, -41.88244, -41.9009, -41.9196, -41.93877, -41.95837, 
        -41.97809, -41.99747, -42.01617, -42.03299, -42.05128, -42.07066, 
        -42.09155, -42.11363, -42.13614, -42.15785, -42.17788, -42.1954, 
        -42.2106, -42.22313, -42.23343, -42.24224, -42.24991, -42.25714, 
        -42.26453, -42.27232, -42.27993, -42.28665, -42.29258, -42.29715, 
        -42.29993, -42.30034, -42.29926, -42.29736, -42.29486, -42.29242, 
        -42.29, -42.28656, -42.28422, -42.28178, -42.27892, -42.2755, 
        -42.27156, -42.26704, -42.26261, -42.25864, -42.25575, -42.25501, 
        -42.25661, -42.26115, -42.26879, -42.27906, -42.29094, -42.30385, 
        -42.31632, -42.32738, -42.33678, -42.3451, -42.35233, -42.35936, 
        -42.36606, -42.37268, -42.37904, -42.38517, -42.39097, -42.39656, 
        -42.40193, -42.40719, -42.41242, -42.41709, -42.42311, -42.42941, 
        -42.43612, -42.44345, -42.45091, -42.45855, -42.46595, -42.47299, 
        -42.47916, -42.48394, -42.48732, -42.48929, -42.48968, -42.48862, 
        -42.48574, -42.48086, -42.47427, -42.46641, -42.45813, -42.4503, 
        -42.44329, -42.43753, -42.43277, -42.42842, -42.42415, -42.41999, 
        -42.41566, -42.41086, -42.40538, -42.39858, -42.38937, -42.37724, 
        -42.36193, -42.3434, -42.3213, -42.29533, -42.265, -42.22957, 
        -42.18798, -42.14261, -42.09278, -42.0388, -41.98064, -41.91748, 
        -41.84853, -41.77274, -41.69017, -41.60086, -41.50536, -41.40554, 
        -41.30345, -41.20103, -41.09991, -41.0026, -40.91135, -40.82702, 
        -40.75046,
  -37.86467, -37.90819, -37.95128, -37.99459, -38.03848, -38.08292, 
        -38.12803, -38.17332, -38.2183, -38.2627, -38.30527, -38.3479, 
        -38.38933, -38.4298, -38.46939, -38.50859, -38.54763, -38.5863, 
        -38.62447, -38.66199, -38.69862, -38.73418, -38.76822, -38.80095, 
        -38.83243, -38.86157, -38.8907, -38.91851, -38.94453, -38.9691, 
        -38.9928, -39.01569, -39.03888, -39.06282, -39.08799, -39.11464, 
        -39.14299, -39.17274, -39.20332, -39.23396, -39.26384, -39.29165, 
        -39.31925, -39.34635, -39.37346, -39.4008, -39.42894, -39.45764, 
        -39.4871, -39.51639, -39.54517, -39.57266, -39.59882, -39.62342, 
        -39.64665, -39.6689, -39.69059, -39.71107, -39.73277, -39.75481, 
        -39.77694, -39.79929, -39.82191, -39.84505, -39.86853, -39.892, 
        -39.91553, -39.93956, -39.96423, -39.98986, -40.01657, -40.04415, 
        -40.07221, -40.09925, -40.12685, -40.15406, -40.18118, -40.20886, 
        -40.23752, -40.26669, -40.29624, -40.32567, -40.3546, -40.38312, 
        -40.41111, -40.43868, -40.46574, -40.49263, -40.51884, -40.54491, 
        -40.57109, -40.59679, -40.62429, -40.65191, -40.67967, -40.70717, 
        -40.7342, -40.76065, -40.78641, -40.81157, -40.83657, -40.86166, 
        -40.88693, -40.91189, -40.93584, -40.95895, -40.98041, -40.99998, 
        -41.01791, -41.03383, -41.04678, -41.05869, -41.06863, -41.07642, 
        -41.0827, -41.08711, -41.08986, -41.09135, -41.09204, -41.09238, 
        -41.09266, -41.0931, -41.09414, -41.09546, -41.09707, -41.09913, 
        -41.10144, -41.1041, -41.10732, -41.11168, -41.11666, -41.12411, 
        -41.13313, -41.14311, -41.15391, -41.16549, -41.17744, -41.19012, 
        -41.20326, -41.21645, -41.22925, -41.24158, -41.25396, -41.26681, 
        -41.2803, -41.29444, -41.30856, -41.32225, -41.33537, -41.34811, 
        -41.36075, -41.37225, -41.38523, -41.39856, -41.41268, -41.42765, 
        -41.44394, -41.46095, -41.47849, -41.49538, -41.51182, -41.52736, 
        -41.54234, -41.5579, -41.5741, -41.59155, -41.61017, -41.62947, 
        -41.64955, -41.66988, -41.68993, -41.70993, -41.72992, -41.74994, 
        -41.76992, -41.78841, -41.80774, -41.82711, -41.84672, -41.86665, 
        -41.88633, -41.90551, -41.92364, -41.94122, -41.95931, -41.97916, 
        -42.00092, -42.02409, -42.04769, -42.07053, -42.0917, -42.11026, 
        -42.12636, -42.13977, -42.15064, -42.15981, -42.16811, -42.17638, 
        -42.18494, -42.19374, -42.20231, -42.20882, -42.21506, -42.21975, 
        -42.22247, -42.22288, -42.22182, -42.21977, -42.21719, -42.21495, 
        -42.21311, -42.21151, -42.21014, -42.20871, -42.20672, -42.20403, 
        -42.20042, -42.19634, -42.19248, -42.18924, -42.18736, -42.18732, 
        -42.18953, -42.19481, -42.20284, -42.21357, -42.22623, -42.23953, 
        -42.2521, -42.26316, -42.27274, -42.28008, -42.28762, -42.29469, 
        -42.30167, -42.30898, -42.3161, -42.32292, -42.32908, -42.33456, 
        -42.33985, -42.34455, -42.34952, -42.35463, -42.36037, -42.36658, 
        -42.37364, -42.38138, -42.38994, -42.39888, -42.40788, -42.41653, 
        -42.42434, -42.43054, -42.43509, -42.43814, -42.43957, -42.4392, 
        -42.43714, -42.43298, -42.42713, -42.41991, -42.41245, -42.4053, 
        -42.39884, -42.39329, -42.3884, -42.38369, -42.37799, -42.3733, 
        -42.3687, -42.36383, -42.35829, -42.35168, -42.34269, -42.33087, 
        -42.31556, -42.29696, -42.27472, -42.24866, -42.2184, -42.1835, 
        -42.14385, -42.09954, -42.05145, -41.99933, -41.94379, -41.88342, 
        -41.81767, -41.74545, -41.66647, -41.58077, -41.48855, -41.39138, 
        -41.29113, -41.18921, -41.08775, -40.98858, -40.89469, -40.80778, 
        -40.72854,
  -37.70686, -37.7495, -37.79216, -37.83551, -37.8799, -37.92477, 
        -37.96918, -38.01475, -38.06001, -38.10442, -38.14772, -38.19034, 
        -38.23163, -38.27193, -38.31156, -38.35079, -38.38963, -38.42841, 
        -38.46677, -38.50454, -38.54027, -38.57594, -38.6102, -38.64297, 
        -38.67423, -38.70416, -38.73292, -38.76043, -38.78669, -38.81142, 
        -38.83538, -38.8591, -38.88322, -38.90812, -38.93444, -38.96115, 
        -38.99063, -39.02145, -39.05302, -39.08457, -39.11538, -39.14525, 
        -39.17405, -39.2024, -39.23066, -39.25897, -39.28771, -39.31716, 
        -39.34719, -39.37704, -39.40638, -39.4335, -39.46024, -39.48561, 
        -39.50956, -39.53262, -39.55522, -39.5774, -39.59973, -39.6222, 
        -39.64481, -39.6677, -39.69095, -39.71477, -39.73897, -39.76335, 
        -39.78798, -39.81316, -39.83839, -39.8658, -39.89426, -39.92325, 
        -39.95224, -39.98104, -40.00935, -40.03728, -40.06521, -40.09378, 
        -40.12312, -40.15296, -40.18337, -40.21392, -40.24405, -40.2734, 
        -40.30211, -40.32906, -40.35634, -40.38278, -40.40891, -40.43525, 
        -40.46175, -40.48878, -40.51691, -40.54519, -40.57375, -40.60204, 
        -40.62963, -40.65622, -40.68188, -40.7067, -40.73108, -40.75557, 
        -40.78033, -40.80424, -40.82866, -40.85198, -40.87426, -40.8946, 
        -40.91332, -40.93026, -40.94512, -40.95789, -40.96822, -40.97633, 
        -40.98216, -40.98598, -40.98818, -40.98937, -40.99012, -40.99081, 
        -40.99168, -40.99286, -40.9943, -40.99509, -40.9971, -40.99928, 
        -41.00171, -41.00444, -41.00765, -41.01162, -41.01703, -41.02396, 
        -41.03278, -41.04272, -41.05344, -41.06503, -41.07702, -41.08968, 
        -41.10307, -41.11653, -41.1296, -41.14237, -41.15543, -41.16872, 
        -41.18162, -41.19608, -41.21046, -41.22469, -41.23844, -41.25194, 
        -41.26512, -41.27837, -41.29177, -41.30562, -41.32017, -41.33616, 
        -41.3532, -41.37071, -41.38913, -41.40684, -41.42376, -41.43973, 
        -41.45523, -41.47103, -41.48736, -41.50448, -41.52241, -41.54, 
        -41.55909, -41.57844, -41.5974, -41.61648, -41.63604, -41.65606, 
        -41.67614, -41.69604, -41.71632, -41.73652, -41.75719, -41.77775, 
        -41.79741, -41.81596, -41.83379, -41.85133, -41.86985, -41.89006, 
        -41.91227, -41.93654, -41.96121, -41.98517, -42.00726, -42.0266, 
        -42.04226, -42.05625, -42.0676, -42.07717, -42.08631, -42.09533, 
        -42.1048, -42.11429, -42.1235, -42.13152, -42.13806, -42.14285, 
        -42.14553, -42.14597, -42.14471, -42.14272, -42.14038, -42.13825, 
        -42.13681, -42.13631, -42.13624, -42.13551, -42.13461, -42.13239, 
        -42.12908, -42.1256, -42.12236, -42.11994, -42.1191, -42.11893, 
        -42.12205, -42.12793, -42.13694, -42.14839, -42.16118, -42.17459, 
        -42.18673, -42.19743, -42.20691, -42.21516, -42.22287, -42.23013, 
        -42.23783, -42.24596, -42.25368, -42.2611, -42.2679, -42.27362, 
        -42.27865, -42.2834, -42.28798, -42.29279, -42.29819, -42.30434, 
        -42.31172, -42.32017, -42.3296, -42.33965, -42.34979, -42.36004, 
        -42.36928, -42.37692, -42.38286, -42.38597, -42.38833, -42.38903, 
        -42.38771, -42.38453, -42.37947, -42.37317, -42.36642, -42.36001, 
        -42.35409, -42.34855, -42.34347, -42.33859, -42.33373, -42.32878, 
        -42.32406, -42.31923, -42.31402, -42.30775, -42.29898, -42.2872, 
        -42.27172, -42.25251, -42.22972, -42.20305, -42.17255, -42.13797, 
        -42.09898, -42.05587, -42.00895, -41.95901, -41.9054, -41.84778, 
        -41.78488, -41.7158, -41.64055, -41.55843, -41.46973, -41.37565, 
        -41.27737, -41.17646, -41.07433, -40.97357, -40.87689, -40.78577, 
        -40.70369,
  -37.5495, -37.59039, -37.63278, -37.67624, -37.72046, -37.76575, 
        -37.81112, -37.85634, -37.90107, -37.94523, -37.98885, -38.03157, 
        -38.07322, -38.11355, -38.15333, -38.19176, -38.23104, -38.27014, 
        -38.30872, -38.34661, -38.38351, -38.41928, -38.45372, -38.48657, 
        -38.51793, -38.54798, -38.57656, -38.60407, -38.63029, -38.65549, 
        -38.67899, -38.70331, -38.72811, -38.75396, -38.78101, -38.8096, 
        -38.8398, -38.87137, -38.90376, -38.93605, -38.96783, -38.99886, 
        -39.02913, -39.05886, -39.08831, -39.11777, -39.14653, -39.17682, 
        -39.20744, -39.23791, -39.26764, -39.29638, -39.32379, -39.34971, 
        -39.37484, -39.39865, -39.42194, -39.44491, -39.46761, -39.49049, 
        -39.51362, -39.53709, -39.56007, -39.58447, -39.6092, -39.63438, 
        -39.65986, -39.6863, -39.71381, -39.74277, -39.77269, -39.80292, 
        -39.83308, -39.86254, -39.89146, -39.92001, -39.94905, -39.97863, 
        -40.00888, -40.03867, -40.0699, -40.10125, -40.13227, -40.16245, 
        -40.19163, -40.21947, -40.24653, -40.27275, -40.29875, -40.325, 
        -40.35191, -40.37983, -40.4085, -40.43789, -40.46757, -40.49646, 
        -40.5248, -40.55081, -40.57643, -40.60071, -40.62437, -40.6479, 
        -40.67178, -40.69619, -40.72078, -40.74463, -40.76788, -40.78947, 
        -40.80938, -40.82739, -40.84333, -40.85716, -40.86828, -40.87636, 
        -40.88229, -40.88591, -40.8864, -40.88671, -40.88713, -40.88766, 
        -40.88897, -40.89071, -40.89301, -40.89548, -40.89777, -40.90053, 
        -40.90354, -40.90653, -40.90975, -40.91389, -40.91928, -40.92603, 
        -40.93432, -40.94388, -40.95434, -40.96578, -40.97805, -40.98979, 
        -41.00323, -41.01695, -41.03045, -41.04382, -41.05752, -41.07154, 
        -41.08602, -41.10082, -41.11554, -41.13008, -41.14446, -41.15857, 
        -41.17261, -41.18657, -41.20074, -41.21516, -41.23046, -41.2468, 
        -41.26423, -41.28255, -41.30112, -41.31837, -41.33566, -41.35191, 
        -41.36782, -41.38376, -41.40008, -41.41681, -41.43418, -41.45216, 
        -41.47019, -41.48837, -41.50657, -41.52504, -41.54387, -41.56341, 
        -41.58361, -41.604, -41.62526, -41.64657, -41.66798, -41.68873, 
        -41.70863, -41.72717, -41.74461, -41.76118, -41.77995, -41.80095, 
        -41.82408, -41.84932, -41.87504, -41.89985, -41.92278, -41.94291, 
        -41.96006, -41.97443, -41.98607, -41.99625, -42.00576, -42.01555, 
        -42.02535, -42.03545, -42.04485, -42.05308, -42.05991, -42.06482, 
        -42.06749, -42.06819, -42.06702, -42.0651, -42.06281, -42.0612, 
        -42.06029, -42.05959, -42.06055, -42.06103, -42.06088, -42.05928, 
        -42.05703, -42.05421, -42.05166, -42.05033, -42.05029, -42.05202, 
        -42.05597, -42.06282, -42.07264, -42.08439, -42.09711, -42.10991, 
        -42.12161, -42.13206, -42.14104, -42.14931, -42.15706, -42.16496, 
        -42.17337, -42.18211, -42.19063, -42.19866, -42.20589, -42.21238, 
        -42.21801, -42.22288, -42.22752, -42.23111, -42.2363, -42.24244, 
        -42.24992, -42.25879, -42.26881, -42.27986, -42.29138, -42.30301, 
        -42.31344, -42.3223, -42.32934, -42.33454, -42.33787, -42.3394, 
        -42.33901, -42.33695, -42.33306, -42.32809, -42.32244, -42.31647, 
        -42.31085, -42.30544, -42.30014, -42.29518, -42.29025, -42.28533, 
        -42.28057, -42.27571, -42.27092, -42.26448, -42.25571, -42.24373, 
        -42.22786, -42.208, -42.18428, -42.15693, -42.12592, -42.0912, 
        -42.0531, -42.01026, -41.96475, -41.91615, -41.86475, -41.80908, 
        -41.74868, -41.68264, -41.61073, -41.5324, -41.44754, -41.35658, 
        -41.26049, -41.16039, -41.05807, -40.95614, -40.85729, -40.76408, 
        -40.67867,
  -37.3918, -37.43335, -37.47563, -37.51875, -37.56279, -37.6077, 
        -37.65249, -37.69709, -37.74136, -37.78554, -37.82885, -37.87083, 
        -37.91316, -37.95437, -37.99455, -38.03455, -38.07432, -38.11367, 
        -38.1524, -38.19017, -38.22694, -38.26266, -38.29718, -38.33034, 
        -38.36208, -38.39143, -38.42029, -38.44785, -38.47439, -38.50005, 
        -38.52514, -38.55013, -38.57557, -38.60187, -38.62943, -38.65842, 
        -38.68905, -38.72105, -38.75402, -38.78713, -38.81987, -38.85109, 
        -38.88277, -38.91404, -38.945, -38.97588, -39.0069, -39.0382, 
        -39.06958, -39.10054, -39.13073, -39.16006, -39.1882, -39.21522, 
        -39.24104, -39.26592, -39.28992, -39.31257, -39.33577, -39.35898, 
        -39.38251, -39.40663, -39.43124, -39.45608, -39.48133, -39.507, 
        -39.53344, -39.56092, -39.58977, -39.61999, -39.65125, -39.68264, 
        -39.71369, -39.74295, -39.77256, -39.80209, -39.83196, -39.8624, 
        -39.89344, -39.92533, -39.95747, -39.98952, -40.02095, -40.05167, 
        -40.08093, -40.10857, -40.13505, -40.1613, -40.18741, -40.21379, 
        -40.24143, -40.2692, -40.29899, -40.3294, -40.35974, -40.38963, 
        -40.41859, -40.44611, -40.4719, -40.49624, -40.51942, -40.54222, 
        -40.56538, -40.5892, -40.61351, -40.63779, -40.66157, -40.68401, 
        -40.7051, -40.72419, -40.74044, -40.75513, -40.7673, -40.7761, 
        -40.78228, -40.78536, -40.78652, -40.78624, -40.78601, -40.78615, 
        -40.78724, -40.78943, -40.79227, -40.79543, -40.79899, -40.80232, 
        -40.80619, -40.80983, -40.81367, -40.81797, -40.82213, -40.82854, 
        -40.83631, -40.84536, -40.85563, -40.86714, -40.8798, -40.89281, 
        -40.9065, -40.92014, -40.93407, -40.94805, -40.96243, -40.9773, 
        -40.99243, -41.00784, -41.02309, -41.03813, -41.05293, -41.06773, 
        -41.0824, -41.09704, -41.11079, -41.12611, -41.14219, -41.15907, 
        -41.17688, -41.1953, -41.21375, -41.23196, -41.24939, -41.26609, 
        -41.28229, -41.29864, -41.31464, -41.33113, -41.34776, -41.36461, 
        -41.38175, -41.39899, -41.41649, -41.43417, -41.45267, -41.47213, 
        -41.49226, -41.51225, -41.53417, -41.55664, -41.57829, -41.5994, 
        -41.61887, -41.6372, -41.65434, -41.672, -41.69153, -41.71342, 
        -41.73779, -41.76369, -41.79026, -41.81612, -41.83999, -41.8611, 
        -41.87875, -41.89347, -41.90568, -41.91614, -41.92598, -41.93595, 
        -41.94597, -41.95605, -41.96564, -41.9732, -41.98025, -41.98528, 
        -41.98813, -41.98896, -41.98794, -41.98608, -41.98397, -41.98249, 
        -41.98228, -41.98327, -41.98495, -41.98662, -41.9876, -41.98737, 
        -41.98605, -41.9844, -41.98297, -41.98221, -41.98294, -41.98563, 
        -41.99083, -41.99849, -42.00861, -42.02052, -42.03297, -42.04498, 
        -42.05606, -42.06564, -42.07404, -42.08216, -42.08917, -42.09762, 
        -42.10653, -42.11576, -42.12493, -42.13377, -42.14198, -42.1493, 
        -42.1557, -42.16122, -42.16611, -42.17077, -42.1759, -42.18213, 
        -42.18991, -42.19919, -42.20985, -42.22173, -42.2344, -42.24697, 
        -42.25846, -42.26822, -42.27635, -42.28251, -42.28693, -42.28961, 
        -42.29059, -42.28981, -42.28734, -42.28366, -42.2788, -42.2734, 
        -42.26778, -42.26239, -42.25683, -42.2515, -42.24551, -42.24062, 
        -42.23586, -42.23114, -42.22596, -42.21946, -42.21051, -42.19825, 
        -42.18208, -42.16152, -42.13694, -42.10876, -42.07714, -42.04263, 
        -42.00507, -41.96436, -41.92048, -41.87378, -41.82353, -41.76948, 
        -41.71137, -41.64799, -41.57917, -41.50439, -41.42314, -41.33533, 
        -41.24147, -41.14272, -41.04092, -40.93793, -40.83731, -40.74158, 
        -40.65311,
  -37.23612, -37.27721, -37.31932, -37.36215, -37.40588, -37.44987, 
        -37.49318, -37.5371, -37.58074, -37.62451, -37.66794, -37.71144, 
        -37.75402, -37.79617, -37.83742, -37.87806, -37.91832, -37.95793, 
        -37.99666, -38.03426, -38.06975, -38.10526, -38.13973, -38.17313, 
        -38.20525, -38.23594, -38.26508, -38.29316, -38.32024, -38.34666, 
        -38.3723, -38.39796, -38.42405, -38.45082, -38.47871, -38.50794, 
        -38.53773, -38.56998, -38.6032, -38.63694, -38.67059, -38.70402, 
        -38.73713, -38.76991, -38.80252, -38.83493, -38.86734, -38.89976, 
        -38.932, -38.9635, -38.99416, -39.02296, -39.05183, -39.07999, 
        -39.10685, -39.13292, -39.15784, -39.18203, -39.20571, -39.22943, 
        -39.2533, -39.27795, -39.30298, -39.32847, -39.35432, -39.38057, 
        -39.40764, -39.43607, -39.46522, -39.49674, -39.52911, -39.56153, 
        -39.59326, -39.62428, -39.65493, -39.68534, -39.71624, -39.74765, 
        -39.77929, -39.81167, -39.84432, -39.87714, -39.90938, -39.94007, 
        -39.96911, -39.9956, -40.02197, -40.04803, -40.07439, -40.10159, 
        -40.13017, -40.15992, -40.19062, -40.2217, -40.25274, -40.28313, 
        -40.3126, -40.34076, -40.36693, -40.39155, -40.41496, -40.43803, 
        -40.4611, -40.48457, -40.50764, -40.53197, -40.55594, -40.57893, 
        -40.60028, -40.62004, -40.63793, -40.65365, -40.66663, -40.67651, 
        -40.68299, -40.68659, -40.6876, -40.68705, -40.68663, -40.68625, 
        -40.68686, -40.68876, -40.6914, -40.69424, -40.69861, -40.70322, 
        -40.70791, -40.71268, -40.71731, -40.72205, -40.72739, -40.73351, 
        -40.74061, -40.74922, -40.75907, -40.77053, -40.7831, -40.79659, 
        -40.81062, -40.8247, -40.8391, -40.85383, -40.86898, -40.88449, 
        -40.89941, -40.91547, -40.9313, -40.94684, -40.96224, -40.97768, 
        -40.99305, -41.00851, -41.02402, -41.04017, -41.05693, -41.07449, 
        -41.09235, -41.11055, -41.12875, -41.1468, -41.1642, -41.18108, 
        -41.19759, -41.21399, -41.23008, -41.24613, -41.26219, -41.27724, 
        -41.29341, -41.30952, -41.32597, -41.34331, -41.36119, -41.38025, 
        -41.40066, -41.42238, -41.44495, -41.46757, -41.48978, -41.51055, 
        -41.52977, -41.54758, -41.56476, -41.58293, -41.6034, -41.62614, 
        -41.65113, -41.67801, -41.70551, -41.73249, -41.75728, -41.77932, 
        -41.79705, -41.81232, -41.82502, -41.83577, -41.8456, -41.85539, 
        -41.86539, -41.87569, -41.8854, -41.89414, -41.9012, -41.90628, 
        -41.90915, -41.90987, -41.9091, -41.90726, -41.90559, -41.90472, 
        -41.90487, -41.9064, -41.90896, -41.91166, -41.91395, -41.9151, 
        -41.915, -41.91422, -41.91383, -41.91415, -41.9159, -41.91857, 
        -41.92471, -41.93312, -41.94386, -41.95575, -41.96776, -41.97903, 
        -41.98896, -41.9975, -42.00548, -42.01325, -42.02106, -42.02974, 
        -42.03897, -42.04865, -42.05858, -42.06827, -42.07742, -42.08585, 
        -42.09336, -42.09993, -42.10551, -42.11058, -42.11592, -42.12246, 
        -42.13049, -42.14031, -42.15171, -42.16449, -42.17765, -42.19089, 
        -42.20303, -42.21337, -42.2223, -42.22864, -42.23428, -42.23832, 
        -42.24072, -42.24117, -42.24016, -42.23766, -42.23375, -42.22892, 
        -42.22337, -42.21772, -42.21209, -42.20643, -42.20116, -42.19597, 
        -42.19093, -42.18594, -42.18043, -42.17371, -42.16449, -42.15208, 
        -42.13558, -42.1147, -42.08935, -42.06071, -42.02866, -41.99414, 
        -41.95715, -41.91758, -41.87557, -41.83002, -41.78148, -41.72903, 
        -41.67236, -41.61111, -41.54509, -41.47339, -41.3954, -41.31047, 
        -41.21898, -41.12214, -41.02113, -40.91838, -40.81649, -40.71775, 
        -40.62648,
  -37.08156, -37.12134, -37.16294, -37.20539, -37.24853, -37.29201, 
        -37.33541, -37.37861, -37.42179, -37.46507, -37.50858, -37.55236, 
        -37.59566, -37.63857, -37.68075, -37.72227, -37.76206, -37.80188, 
        -37.8404, -37.87773, -37.91386, -37.94894, -37.98333, -38.0168, 
        -38.04937, -38.08064, -38.11044, -38.13903, -38.16666, -38.19352, 
        -38.21904, -38.24553, -38.27222, -38.2995, -38.32775, -38.35723, 
        -38.38817, -38.42051, -38.45404, -38.48827, -38.52279, -38.55731, 
        -38.59174, -38.62598, -38.66013, -38.69411, -38.72686, -38.76034, 
        -38.79325, -38.82538, -38.8566, -38.8871, -38.91704, -38.9462, 
        -38.97434, -39.00117, -39.02699, -39.05191, -39.07611, -39.1004, 
        -39.12485, -39.1498, -39.17447, -39.20063, -39.22708, -39.25386, 
        -39.28172, -39.311, -39.34218, -39.37499, -39.40841, -39.4416, 
        -39.47412, -39.50583, -39.53732, -39.56894, -39.6008, -39.6329, 
        -39.66511, -39.69685, -39.73008, -39.76313, -39.79558, -39.82673, 
        -39.85591, -39.88326, -39.9097, -39.93584, -39.96271, -39.99091, 
        -40.0203, -40.05098, -40.08231, -40.11383, -40.14537, -40.17636, 
        -40.20612, -40.23369, -40.26076, -40.28608, -40.30983, -40.33332, 
        -40.35683, -40.38063, -40.40496, -40.42952, -40.45362, -40.47652, 
        -40.49794, -40.5177, -40.53585, -40.55174, -40.56516, -40.57571, 
        -40.58297, -40.58693, -40.58861, -40.58762, -40.58685, -40.58649, 
        -40.58693, -40.58855, -40.59118, -40.59507, -40.6, -40.60544, 
        -40.61131, -40.61714, -40.62265, -40.62792, -40.63342, -40.63951, 
        -40.64631, -40.6543, -40.66373, -40.67487, -40.68725, -40.69969, 
        -40.71395, -40.72864, -40.74406, -40.75985, -40.77595, -40.79233, 
        -40.80883, -40.82536, -40.84162, -40.8577, -40.87371, -40.88981, 
        -40.90615, -40.92265, -40.93946, -40.95667, -40.97399, -40.99147, 
        -41.00928, -41.02712, -41.04485, -41.06127, -41.07846, -41.09565, 
        -41.11255, -41.12887, -41.14487, -41.1609, -41.17656, -41.19192, 
        -41.20701, -41.22206, -41.23796, -41.25477, -41.27264, -41.29147, 
        -41.31189, -41.33364, -41.35606, -41.37854, -41.40042, -41.42097, 
        -41.43972, -41.45744, -41.47517, -41.49365, -41.51366, -41.53699, 
        -41.56282, -41.59071, -41.61902, -41.64696, -41.67302, -41.69629, 
        -41.71613, -41.73218, -41.74519, -41.75611, -41.76627, -41.77618, 
        -41.78609, -41.79601, -41.80596, -41.81458, -41.82199, -41.82706, 
        -41.82978, -41.83078, -41.82996, -41.82856, -41.82736, -41.82694, 
        -41.82768, -41.82883, -41.83208, -41.83563, -41.83882, -41.84099, 
        -41.84184, -41.84213, -41.8426, -41.84401, -41.84682, -41.85165, 
        -41.85863, -41.86797, -41.87918, -41.89108, -41.90272, -41.91313, 
        -41.92208, -41.9299, -41.9371, -41.9444, -41.95211, -41.96055, 
        -41.97003, -41.98023, -41.99077, -42.00136, -42.01156, -42.02129, 
        -42.03016, -42.03781, -42.04439, -42.04919, -42.0551, -42.06216, 
        -42.07078, -42.08129, -42.09351, -42.10684, -42.12048, -42.13364, 
        -42.14591, -42.15675, -42.16632, -42.17464, -42.18159, -42.18686, 
        -42.19048, -42.19239, -42.1928, -42.1916, -42.18874, -42.18438, 
        -42.17915, -42.17342, -42.16769, -42.16199, -42.15625, -42.15064, 
        -42.14514, -42.13965, -42.13363, -42.12645, -42.11694, -42.10423, 
        -42.08752, -42.06631, -42.04081, -42.01163, -41.97953, -41.94525, 
        -41.90894, -41.86966, -41.82894, -41.78481, -41.73741, -41.68616, 
        -41.63098, -41.57159, -41.50777, -41.43855, -41.36333, -41.28134, 
        -41.19235, -41.09768, -40.99825, -40.89609, -40.79386, -40.69452, 
        -40.60074,
  -36.92733, -36.96775, -37.00877, -37.05066, -37.09316, -37.13599, 
        -37.17871, -37.22131, -37.26408, -37.30709, -37.35059, -37.39341, 
        -37.43727, -37.48086, -37.52376, -37.56588, -37.60704, -37.647, 
        -37.68561, -37.72261, -37.75843, -37.79333, -37.82749, -37.86108, 
        -37.89378, -37.9244, -37.95468, -37.98388, -38.01225, -38.0401, 
        -38.06754, -38.09492, -38.12246, -38.15046, -38.17924, -38.20911, 
        -38.24029, -38.27281, -38.30654, -38.34119, -38.37634, -38.41078, 
        -38.4463, -38.48188, -38.51733, -38.55269, -38.58763, -38.62204, 
        -38.6557, -38.68853, -38.72034, -38.75163, -38.78241, -38.81253, 
        -38.84182, -38.86978, -38.8965, -38.92113, -38.94611, -38.97084, 
        -38.99591, -39.02157, -39.04763, -39.07449, -39.10151, -39.12902, 
        -39.15759, -39.18776, -39.21989, -39.25362, -39.28807, -39.32214, 
        -39.35557, -39.38839, -39.41974, -39.45196, -39.48451, -39.51704, 
        -39.54973, -39.58264, -39.61595, -39.64936, -39.68204, -39.71332, 
        -39.74307, -39.77112, -39.79793, -39.82473, -39.85212, -39.88108, 
        -39.91116, -39.94151, -39.97348, -40.00512, -40.03686, -40.06833, 
        -40.09872, -40.12793, -40.15574, -40.18179, -40.20648, -40.23051, 
        -40.25426, -40.27859, -40.30336, -40.32821, -40.35256, -40.37563, 
        -40.39703, -40.41657, -40.43346, -40.44946, -40.46278, -40.47342, 
        -40.48092, -40.48557, -40.4878, -40.48857, -40.48848, -40.48856, 
        -40.48908, -40.49068, -40.4934, -40.4974, -40.50271, -40.50864, 
        -40.51533, -40.52207, -40.52836, -40.53428, -40.53918, -40.54535, 
        -40.55198, -40.55973, -40.56878, -40.57946, -40.59167, -40.60523, 
        -40.61967, -40.63503, -40.65111, -40.66784, -40.68509, -40.70237, 
        -40.7197, -40.73677, -40.75354, -40.76999, -40.78638, -40.80298, 
        -40.82004, -40.83765, -40.85447, -40.87261, -40.89087, -40.90893, 
        -40.92665, -40.94397, -40.96093, -40.97789, -40.99476, -41.01184, 
        -41.02887, -41.04536, -41.06121, -41.077, -41.09242, -41.10716, 
        -41.12182, -41.13641, -41.15185, -41.16803, -41.18528, -41.20411, 
        -41.22433, -41.24487, -41.26695, -41.28909, -41.31049, -41.33058, 
        -41.34904, -41.36662, -41.38456, -41.4035, -41.42463, -41.44859, 
        -41.47494, -41.50331, -41.53272, -41.56158, -41.5887, -41.61295, 
        -41.63361, -41.65035, -41.66403, -41.67566, -41.68627, -41.69645, 
        -41.70656, -41.71692, -41.72692, -41.7359, -41.74223, -41.74717, 
        -41.74983, -41.75079, -41.75075, -41.74948, -41.74868, -41.74876, 
        -41.75011, -41.75265, -41.75632, -41.76046, -41.76414, -41.76686, 
        -41.76848, -41.76978, -41.77109, -41.77325, -41.77726, -41.78336, 
        -41.79154, -41.80163, -41.81326, -41.82496, -41.83587, -41.84554, 
        -41.85406, -41.86137, -41.86808, -41.87492, -41.88132, -41.88989, 
        -41.89952, -41.91016, -41.92126, -41.93273, -41.94397, -41.95491, 
        -41.96509, -41.97418, -41.98193, -41.98877, -41.9956, -42.0035, 
        -42.01286, -42.02397, -42.03667, -42.05029, -42.06399, -42.07723, 
        -42.08947, -42.10064, -42.11088, -42.12016, -42.12808, -42.13448, 
        -42.13927, -42.14251, -42.14415, -42.14411, -42.14226, -42.1387, 
        -42.13385, -42.12836, -42.12267, -42.117, -42.11014, -42.10427, 
        -42.09833, -42.09219, -42.08545, -42.07763, -42.06784, -42.05471, 
        -42.03759, -42.01609, -41.99035, -41.96107, -41.92908, -41.89515, 
        -41.85946, -41.82241, -41.78292, -41.74032, -41.69415, -41.64418, 
        -41.59017, -41.53211, -41.46991, -41.40266, -41.32985, -41.25038, 
        -41.16383, -41.07138, -40.9738, -40.87289, -40.77084, -40.67027, 
        -40.57444,
  -36.77528, -36.81532, -36.85595, -36.89726, -36.93911, -36.98117, 
        -37.02228, -37.06438, -37.10692, -37.1498, -37.19328, -37.23725, 
        -37.2814, -37.32529, -37.36857, -37.41097, -37.45245, -37.49247, 
        -37.5311, -37.56808, -37.60363, -37.6374, -37.67165, -37.70527, 
        -37.73824, -37.77012, -37.80086, -37.83065, -37.85982, -37.88859, 
        -37.9171, -37.94551, -37.97407, -38.00296, -38.03255, -38.06308, 
        -38.09371, -38.12653, -38.1605, -38.19546, -38.23114, -38.26733, 
        -38.30386, -38.34062, -38.37717, -38.41351, -38.44931, -38.4844, 
        -38.51863, -38.55195, -38.58461, -38.61567, -38.6473, -38.67834, 
        -38.70863, -38.73759, -38.76521, -38.79172, -38.81744, -38.84291, 
        -38.8685, -38.89468, -38.92121, -38.94847, -38.97647, -39.00476, 
        -39.03421, -39.06538, -39.09728, -39.13176, -39.16713, -39.20236, 
        -39.23691, -39.27065, -39.30381, -39.33676, -39.36954, -39.40224, 
        -39.43498, -39.468, -39.50147, -39.53516, -39.56833, -39.60025, 
        -39.63056, -39.65835, -39.68593, -39.71369, -39.74157, -39.77082, 
        -39.80161, -39.83319, -39.86535, -39.89755, -39.9296, -39.96142, 
        -39.99243, -40.02256, -40.05112, -40.07803, -40.10368, -40.12867, 
        -40.15322, -40.17812, -40.20222, -40.2272, -40.25151, -40.27454, 
        -40.29588, -40.31543, -40.33324, -40.34878, -40.3617, -40.37219, 
        -40.37994, -40.38498, -40.38793, -40.38963, -40.39049, -40.39114, 
        -40.39225, -40.39401, -40.39713, -40.40052, -40.40613, -40.41264, 
        -40.41977, -40.42723, -40.434, -40.4402, -40.44664, -40.45303, 
        -40.45994, -40.46752, -40.47648, -40.48676, -40.49854, -40.51184, 
        -40.52631, -40.54216, -40.55903, -40.57673, -40.59493, -40.61324, 
        -40.63036, -40.64809, -40.66547, -40.68245, -40.69942, -40.71646, 
        -40.73394, -40.75208, -40.7707, -40.78988, -40.80909, -40.8275, 
        -40.84512, -40.86211, -40.87875, -40.8954, -40.91214, -40.929, 
        -40.94582, -40.96217, -40.97779, -40.99313, -41.00818, -41.02174, 
        -41.03609, -41.05022, -41.06524, -41.08121, -41.09831, -41.11661, 
        -41.13654, -41.15771, -41.17933, -41.20115, -41.22233, -41.24218, 
        -41.26036, -41.278, -41.29585, -41.31499, -41.33639, -41.36066, 
        -41.38765, -41.41622, -41.4461, -41.47567, -41.50349, -41.52871, 
        -41.55046, -41.56724, -41.58185, -41.59435, -41.60575, -41.61672, 
        -41.62769, -41.63841, -41.64857, -41.65756, -41.66446, -41.66945, 
        -41.67192, -41.67252, -41.67252, -41.67178, -41.67143, -41.6721, 
        -41.67392, -41.67696, -41.68084, -41.68495, -41.68884, -41.6921, 
        -41.69445, -41.69626, -41.69829, -41.70138, -41.70609, -41.71207, 
        -41.72136, -41.7321, -41.74374, -41.75508, -41.76588, -41.77585, 
        -41.78407, -41.79109, -41.79756, -41.80425, -41.81168, -41.82034, 
        -41.83029, -41.84139, -41.85324, -41.8653, -41.87732, -41.88926, 
        -41.9006, -41.91086, -41.91982, -41.92806, -41.93616, -41.94504, 
        -41.95515, -41.96687, -41.97989, -41.99345, -42.00707, -42.02025, 
        -42.03249, -42.04412, -42.05504, -42.06409, -42.07289, -42.08029, 
        -42.08615, -42.09033, -42.09302, -42.09408, -42.09319, -42.09056, 
        -42.08642, -42.08141, -42.0761, -42.07068, -42.06505, -42.05917, 
        -42.05282, -42.04603, -42.0387, -42.03024, -42.01969, -42.00583, 
        -41.9882, -41.96645, -41.94062, -41.91131, -41.87955, -41.84606, 
        -41.81141, -41.77539, -41.73732, -41.6962, -41.65113, -41.60208, 
        -41.54913, -41.4923, -41.43124, -41.36548, -41.29429, -41.21689, 
        -41.13248, -41.04211, -40.94647, -40.84678, -40.74522, -40.64406, 
        -40.54519,
  -36.62446, -36.66296, -36.7031, -36.74376, -36.78514, -36.8266, 
        -36.86833, -36.91039, -36.95276, -36.99575, -37.03932, -37.08341, 
        -37.12757, -37.17161, -37.21484, -37.25721, -37.29747, -37.33752, 
        -37.37613, -37.41308, -37.44871, -37.48345, -37.51779, -37.55158, 
        -37.58477, -37.61703, -37.64827, -37.67872, -37.70888, -37.73861, 
        -37.76844, -37.79702, -37.82666, -37.85677, -37.88739, -37.91883, 
        -37.9511, -37.98434, -38.01854, -38.05377, -38.08979, -38.12656, 
        -38.16393, -38.2015, -38.23898, -38.27607, -38.31131, -38.34679, 
        -38.38143, -38.41526, -38.44855, -38.48153, -38.5139, -38.54569, 
        -38.57659, -38.60645, -38.63494, -38.66237, -38.68903, -38.71532, 
        -38.74165, -38.7683, -38.79461, -38.8225, -38.8511, -38.88044, 
        -38.91086, -38.94279, -38.97647, -39.01176, -39.0479, -39.08406, 
        -39.11979, -39.15468, -39.18886, -39.2224, -39.2554, -39.28798, 
        -39.32059, -39.35341, -39.38596, -39.41978, -39.45351, -39.4866, 
        -39.51809, -39.54796, -39.5763, -39.60466, -39.63333, -39.6627, 
        -39.69383, -39.72525, -39.75734, -39.78975, -39.82209, -39.85442, 
        -39.88631, -39.91716, -39.94567, -39.97363, -40.00031, -40.02617, 
        -40.0518, -40.07743, -40.10312, -40.12825, -40.15256, -40.17526, 
        -40.19648, -40.2158, -40.23336, -40.24842, -40.2612, -40.27134, 
        -40.2792, -40.28501, -40.28913, -40.29096, -40.29261, -40.29382, 
        -40.29552, -40.29795, -40.3017, -40.30656, -40.31256, -40.31966, 
        -40.32733, -40.33488, -40.34179, -40.34823, -40.35486, -40.36141, 
        -40.36853, -40.37642, -40.38562, -40.39611, -40.40755, -40.41961, 
        -40.43394, -40.44986, -40.46704, -40.48544, -40.50443, -40.52349, 
        -40.54247, -40.56107, -40.57914, -40.59675, -40.61412, -40.63162, 
        -40.64965, -40.66819, -40.68745, -40.70726, -40.72698, -40.74583, 
        -40.76366, -40.78075, -40.7972, -40.81256, -40.829, -40.84542, 
        -40.86162, -40.87746, -40.89295, -40.90817, -40.92298, -40.93739, 
        -40.95149, -40.96558, -40.98032, -40.99597, -41.01295, -41.03113, 
        -41.05038, -41.07095, -41.09195, -41.11313, -41.13372, -41.15279, 
        -41.17105, -41.18901, -41.20714, -41.22656, -41.24759, -41.27208, 
        -41.29916, -41.32828, -41.35836, -41.3882, -41.41691, -41.44304, 
        -41.46575, -41.48473, -41.50061, -41.51432, -41.52687, -41.53907, 
        -41.5508, -41.56197, -41.57204, -41.58098, -41.58788, -41.59237, 
        -41.59471, -41.59517, -41.59475, -41.59448, -41.59477, -41.59605, 
        -41.59839, -41.60042, -41.60437, -41.60854, -41.61282, -41.6164, 
        -41.61915, -41.62145, -41.62399, -41.62765, -41.63316, -41.64083, 
        -41.65039, -41.66137, -41.67315, -41.68489, -41.69588, -41.70561, 
        -41.71392, -41.72117, -41.72795, -41.73494, -41.74284, -41.75196, 
        -41.76234, -41.77396, -41.78612, -41.79882, -41.8118, -41.82421, 
        -41.8363, -41.84736, -41.85756, -41.86611, -41.87566, -41.88548, 
        -41.89634, -41.90839, -41.92142, -41.93495, -41.94852, -41.96171, 
        -41.97419, -41.9863, -41.99791, -42.00875, -42.01812, -42.02647, 
        -42.03297, -42.03783, -42.04119, -42.04308, -42.04329, -42.04186, 
        -42.03888, -42.0348, -42.03016, -42.02523, -42.02008, -42.01437, 
        -42.00793, -42.00088, -41.99266, -41.98341, -41.97186, -41.95751, 
        -41.93922, -41.91695, -41.89098, -41.86174, -41.83043, -41.79758, 
        -41.76393, -41.7281, -41.69156, -41.65176, -41.60791, -41.55958, 
        -41.50737, -41.45142, -41.39138, -41.32674, -41.25671, -41.18052, 
        -41.0978, -41.00909, -40.91478, -40.81632, -40.71493, -40.613, 
        -40.51357,
  -36.47437, -36.51336, -36.55291, -36.59318, -36.63409, -36.67531, 
        -36.71681, -36.75868, -36.80112, -36.84425, -36.88803, -36.93119, 
        -36.97531, -37.01899, -37.0619, -37.10393, -37.14488, -37.18488, 
        -37.22343, -37.26043, -37.29604, -37.33081, -37.36519, -37.39942, 
        -37.4329, -37.46552, -37.49636, -37.52779, -37.55899, -37.58997, 
        -37.6208, -37.65147, -37.68245, -37.71376, -37.74557, -37.77797, 
        -37.81099, -37.84476, -37.87925, -37.91459, -37.95092, -37.98711, 
        -38.02505, -38.06336, -38.10146, -38.13904, -38.17573, -38.21156, 
        -38.24657, -38.28093, -38.31474, -38.34811, -38.381, -38.41331, 
        -38.44477, -38.47528, -38.50473, -38.53209, -38.55982, -38.58716, 
        -38.61445, -38.64193, -38.67001, -38.69866, -38.72799, -38.75825, 
        -38.78958, -38.82245, -38.85699, -38.89309, -38.93001, -38.96704, 
        -39.00376, -39.03982, -39.07381, -39.10795, -39.14122, -39.17386, 
        -39.20631, -39.23918, -39.27251, -39.30656, -39.34053, -39.37417, 
        -39.40672, -39.43786, -39.46739, -39.49611, -39.52494, -39.55437, 
        -39.58519, -39.61691, -39.64808, -39.68058, -39.7133, -39.74616, 
        -39.7788, -39.81057, -39.84075, -39.86983, -39.89757, -39.92438, 
        -39.95112, -39.97775, -40.00393, -40.02936, -40.05344, -40.07607, 
        -40.09687, -40.11575, -40.13185, -40.14667, -40.15916, -40.16953, 
        -40.17796, -40.18467, -40.19006, -40.1941, -40.19707, -40.19937, 
        -40.20186, -40.20469, -40.20887, -40.21436, -40.22087, -40.22819, 
        -40.23603, -40.24375, -40.25098, -40.25776, -40.2633, -40.27027, 
        -40.27777, -40.28601, -40.29547, -40.30596, -40.31785, -40.33088, 
        -40.34541, -40.3615, -40.37873, -40.39713, -40.41644, -40.43606, 
        -40.45559, -40.47483, -40.49355, -40.51183, -40.52979, -40.54776, 
        -40.56612, -40.58513, -40.60373, -40.62381, -40.64381, -40.66292, 
        -40.68085, -40.69786, -40.71428, -40.73043, -40.74662, -40.7625, 
        -40.77821, -40.79371, -40.80885, -40.82401, -40.83879, -40.85326, 
        -40.86752, -40.88204, -40.89695, -40.91254, -40.92898, -40.9464, 
        -40.96497, -40.98342, -41.00339, -41.02361, -41.04374, -41.06279, 
        -41.08118, -41.09943, -41.11805, -41.13784, -41.15998, -41.18476, 
        -41.2122, -41.24162, -41.27199, -41.3023, -41.33145, -41.35806, 
        -41.38167, -41.40175, -41.41893, -41.43427, -41.44838, -41.46175, 
        -41.47455, -41.48626, -41.49671, -41.50542, -41.51107, -41.51534, 
        -41.51717, -41.51743, -41.51713, -41.51714, -41.51786, -41.5197, 
        -41.52222, -41.52553, -41.52958, -41.53381, -41.53796, -41.5417, 
        -41.54461, -41.54733, -41.55053, -41.55479, -41.56076, -41.56857, 
        -41.57848, -41.58989, -41.60177, -41.61354, -41.62463, -41.63438, 
        -41.6431, -41.65097, -41.65843, -41.6662, -41.67387, -41.68373, 
        -41.69484, -41.70675, -41.71953, -41.73264, -41.7459, -41.75882, 
        -41.77139, -41.78323, -41.79454, -41.8053, -41.81603, -41.82689, 
        -41.83842, -41.85064, -41.86377, -41.87716, -41.89058, -41.90369, 
        -41.91645, -41.92914, -41.94146, -41.95291, -41.96311, -41.97192, 
        -41.97886, -41.98405, -41.98784, -41.99015, -41.99147, -41.99135, 
        -41.98986, -41.98712, -41.98353, -41.9794, -41.97472, -41.96832, 
        -41.96191, -41.9544, -41.9457, -41.93544, -41.92323, -41.90812, 
        -41.8895, -41.86696, -41.84082, -41.8118, -41.78099, -41.74913, 
        -41.71655, -41.68305, -41.64772, -41.60934, -41.5667, -41.51908, 
        -41.46717, -41.41183, -41.35251, -41.28862, -41.21943, -41.14419, 
        -41.06263, -40.97475, -40.8812, -40.78292, -40.68137, -40.57844, 
        -40.47704,
  -36.32677, -36.36522, -36.40432, -36.44422, -36.48483, -36.52591, 
        -36.56649, -36.60865, -36.65136, -36.69471, -36.73864, -36.78291, 
        -36.82676, -36.86987, -36.91222, -36.95375, -36.99419, -37.03379, 
        -37.07222, -37.10925, -37.14488, -37.17873, -37.21335, -37.24783, 
        -37.28189, -37.31525, -37.34818, -37.38054, -37.41285, -37.44474, 
        -37.47648, -37.50834, -37.54037, -37.57281, -37.60577, -37.63918, 
        -37.67197, -37.70616, -37.74095, -37.77651, -37.81306, -37.85074, 
        -37.88913, -37.92786, -37.96638, -38.00424, -38.04122, -38.07736, 
        -38.11279, -38.14752, -38.18172, -38.21542, -38.24762, -38.2802, 
        -38.31222, -38.34325, -38.37336, -38.40286, -38.43183, -38.46037, 
        -38.48891, -38.51754, -38.54652, -38.57598, -38.60614, -38.6372, 
        -38.6696, -38.70345, -38.7379, -38.77486, -38.8126, -38.85057, 
        -38.88816, -38.92498, -38.96088, -38.99552, -39.02913, -39.0621, 
        -39.09457, -39.12745, -39.1608, -39.19479, -39.22914, -39.26316, 
        -39.2963, -39.32787, -39.35709, -39.38638, -39.41555, -39.44524, 
        -39.47594, -39.50739, -39.53959, -39.57231, -39.60547, -39.63885, 
        -39.6717, -39.70419, -39.73519, -39.76529, -39.79389, -39.82248, 
        -39.85028, -39.87767, -39.90338, -39.92888, -39.95299, -39.97525, 
        -39.99555, -40.01409, -40.03064, -40.04501, -40.0574, -40.06818, 
        -40.07742, -40.08534, -40.09242, -40.09835, -40.10286, -40.10651, 
        -40.10979, -40.11364, -40.11838, -40.12398, -40.12962, -40.13712, 
        -40.14515, -40.15298, -40.16037, -40.16755, -40.1747, -40.18206, 
        -40.19013, -40.19886, -40.20848, -40.2191, -40.23106, -40.24424, 
        -40.2589, -40.27494, -40.29233, -40.31096, -40.33046, -40.3505, 
        -40.37059, -40.38933, -40.40845, -40.4273, -40.44569, -40.46369, 
        -40.48214, -40.50136, -40.521, -40.54117, -40.5611, -40.58044, 
        -40.59864, -40.61574, -40.63207, -40.64821, -40.66383, -40.67931, 
        -40.69456, -40.70966, -40.72462, -40.73967, -40.75465, -40.76867, 
        -40.78363, -40.79862, -40.81371, -40.8294, -40.84538, -40.86174, 
        -40.87904, -40.89728, -40.91636, -40.93569, -40.95524, -40.97439, 
        -40.99297, -41.01146, -41.03059, -41.05121, -41.07381, -41.09922, 
        -41.12695, -41.15677, -41.18738, -41.21777, -41.24714, -41.27428, 
        -41.29845, -41.31861, -41.33718, -41.35399, -41.36963, -41.38459, 
        -41.39847, -41.41102, -41.42173, -41.4305, -41.43689, -41.44078, 
        -41.44232, -41.44225, -41.44186, -41.44195, -41.44283, -41.44505, 
        -41.4478, -41.45127, -41.45515, -41.45936, -41.46335, -41.46702, 
        -41.47033, -41.47329, -41.47694, -41.48156, -41.48794, -41.49635, 
        -41.50574, -41.51733, -41.52928, -41.54091, -41.55177, -41.56189, 
        -41.57096, -41.57961, -41.58821, -41.59723, -41.60704, -41.61778, 
        -41.62946, -41.642, -41.65501, -41.66832, -41.68181, -41.69519, 
        -41.70824, -41.72087, -41.73313, -41.74501, -41.75663, -41.76839, 
        -41.78028, -41.79277, -41.80571, -41.81891, -41.83237, -41.84568, 
        -41.85892, -41.87219, -41.88515, -41.89724, -41.90706, -41.916, 
        -41.92308, -41.92834, -41.93208, -41.93518, -41.93739, -41.9387, 
        -41.9386, -41.93729, -41.93489, -41.93159, -41.92756, -41.92244, 
        -41.91616, -41.90845, -41.89916, -41.88831, -41.87546, -41.8598, 
        -41.84077, -41.81819, -41.79211, -41.76374, -41.73383, -41.70285, 
        -41.67138, -41.63935, -41.60522, -41.56801, -41.52641, -41.47952, 
        -41.42801, -41.37263, -41.3138, -41.25045, -41.18162, -41.1069, 
        -41.02586, -40.93829, -40.84486, -40.74619, -40.64352, -40.53892, 
        -40.43391,
  -36.18062, -36.21745, -36.25613, -36.2957, -36.3362, -36.37749, 
        -36.41939, -36.46194, -36.50515, -36.5489, -36.59304, -36.63697, 
        -36.68042, -36.72289, -36.76467, -36.80552, -36.8446, -36.88383, 
        -36.9221, -36.95901, -36.99472, -37.02969, -37.06451, -37.09926, 
        -37.13378, -37.16835, -37.20241, -37.23586, -37.26888, -37.30162, 
        -37.33414, -37.3657, -37.39864, -37.43205, -37.46607, -37.50056, 
        -37.53514, -37.5699, -37.60505, -37.64091, -37.67779, -37.71572, 
        -37.75444, -37.79353, -37.83232, -37.87032, -37.90654, -37.94293, 
        -37.97855, -38.01367, -38.04815, -38.082, -38.11532, -38.14817, 
        -38.18046, -38.21191, -38.243, -38.27374, -38.3039, -38.3339, 
        -38.3639, -38.39384, -38.42396, -38.4533, -38.48438, -38.51635, 
        -38.54967, -38.58461, -38.62128, -38.65911, -38.69779, -38.73658, 
        -38.77478, -38.81225, -38.84852, -38.88374, -38.91772, -38.95092, 
        -38.98367, -39.01672, -39.04906, -39.08319, -39.11756, -39.15174, 
        -39.18505, -39.21728, -39.24801, -39.27771, -39.30715, -39.33699, 
        -39.36774, -39.39943, -39.4318, -39.46466, -39.49789, -39.53136, 
        -39.56477, -39.59748, -39.62875, -39.65936, -39.6893, -39.71849, 
        -39.7472, -39.77549, -39.80282, -39.82871, -39.85283, -39.87476, 
        -39.89472, -39.91265, -39.9287, -39.94265, -39.95509, -39.96624, 
        -39.97639, -39.98584, -39.99444, -40.00085, -40.00729, -40.01283, 
        -40.01777, -40.0228, -40.02828, -40.03447, -40.04134, -40.0487, 
        -40.05657, -40.0642, -40.07187, -40.07948, -40.08729, -40.09539, 
        -40.10426, -40.11364, -40.12358, -40.13441, -40.14631, -40.15842, 
        -40.17318, -40.18947, -40.20713, -40.22614, -40.24588, -40.26625, 
        -40.28656, -40.3066, -40.32605, -40.34498, -40.36354, -40.38197, 
        -40.40055, -40.41961, -40.43904, -40.45894, -40.47871, -40.49806, 
        -40.51646, -40.53394, -40.55038, -40.5663, -40.58068, -40.59549, 
        -40.61016, -40.62501, -40.64013, -40.65538, -40.67076, -40.6861, 
        -40.70165, -40.71737, -40.73286, -40.74804, -40.76325, -40.77861, 
        -40.79479, -40.81174, -40.82973, -40.84848, -40.86752, -40.88655, 
        -40.90541, -40.92444, -40.94432, -40.96587, -40.98832, -41.01431, 
        -41.04274, -41.07293, -41.10376, -41.13406, -41.16327, -41.19047, 
        -41.2153, -41.23752, -41.25747, -41.27574, -41.29304, -41.30945, 
        -41.32434, -41.33775, -41.34895, -41.35769, -41.36407, -41.3675, 
        -41.36853, -41.36822, -41.36768, -41.36775, -41.36886, -41.3709, 
        -41.37388, -41.37735, -41.38021, -41.38429, -41.38837, -41.39209, 
        -41.39538, -41.39867, -41.40253, -41.40779, -41.41545, -41.42455, 
        -41.4352, -41.44644, -41.45822, -41.4694, -41.48009, -41.49044, 
        -41.49997, -41.5094, -41.51911, -41.5295, -41.54065, -41.55256, 
        -41.56487, -41.57785, -41.59112, -41.60479, -41.61855, -41.63234, 
        -41.64588, -41.65911, -41.67216, -41.68488, -41.69652, -41.70865, 
        -41.72089, -41.73336, -41.74615, -41.75946, -41.77312, -41.78687, 
        -41.80077, -41.81462, -41.82824, -41.84092, -41.85217, -41.86136, 
        -41.86831, -41.87336, -41.87722, -41.8807, -41.88363, -41.88596, 
        -41.88716, -41.88708, -41.88585, -41.88334, -41.8796, -41.87477, 
        -41.86858, -41.86104, -41.85187, -41.84074, -41.82754, -41.81159, 
        -41.79261, -41.77015, -41.74463, -41.71688, -41.68769, -41.65784, 
        -41.6276, -41.59666, -41.56274, -41.52623, -41.48529, -41.4391, 
        -41.38817, -41.3332, -41.2744, -41.21115, -41.14251, -41.06789, 
        -40.98684, -40.89907, -40.805, -40.70518, -40.60073, -40.49359, 
        -40.38662,
  -36.03423, -36.07157, -36.10989, -36.14943, -36.19015, -36.23186, 
        -36.27439, -36.31758, -36.36133, -36.40546, -36.44956, -36.4922, 
        -36.53502, -36.57692, -36.61793, -36.6581, -36.69764, -36.73666, 
        -36.77459, -36.81153, -36.8476, -36.88302, -36.91825, -36.95358, 
        -36.98886, -37.02412, -37.05792, -37.09248, -37.12637, -37.15968, 
        -37.19247, -37.2254, -37.25884, -37.29294, -37.32795, -37.36326, 
        -37.39883, -37.43452, -37.47045, -37.50688, -37.54435, -37.5816, 
        -37.6204, -37.65934, -37.69802, -37.73605, -37.77324, -37.80963, 
        -37.84547, -37.8808, -37.91561, -37.94985, -37.98345, -38.01655, 
        -38.04901, -38.08136, -38.11342, -38.14406, -38.17554, -38.20678, 
        -38.23785, -38.26897, -38.30038, -38.33189, -38.36404, -38.39719, 
        -38.43172, -38.46793, -38.50567, -38.54457, -38.5841, -38.62344, 
        -38.66219, -38.70004, -38.73565, -38.77108, -38.8054, -38.83899, 
        -38.87228, -38.90553, -38.93926, -38.97335, -39.00777, -39.04217, 
        -39.07579, -39.10791, -39.13905, -39.16943, -39.1991, -39.22915, 
        -39.26014, -39.29174, -39.32343, -39.35654, -39.39012, -39.4236, 
        -39.45726, -39.49055, -39.52315, -39.55463, -39.58547, -39.61559, 
        -39.64492, -39.67381, -39.7015, -39.72741, -39.75169, -39.77361, 
        -39.79351, -39.81123, -39.82693, -39.83992, -39.85247, -39.86413, 
        -39.87527, -39.88594, -39.89583, -39.90476, -39.91269, -39.92, 
        -39.92676, -39.9333, -39.93984, -39.94683, -39.95395, -39.96125, 
        -39.96883, -39.97641, -39.98421, -39.99213, -40.00044, -40.0085, 
        -40.01793, -40.02808, -40.03881, -40.05022, -40.06262, -40.07602, 
        -40.09076, -40.10731, -40.12522, -40.1447, -40.16478, -40.18539, 
        -40.20589, -40.22615, -40.24569, -40.26451, -40.28311, -40.30146, 
        -40.31998, -40.33884, -40.3572, -40.3769, -40.39659, -40.41583, 
        -40.43438, -40.45208, -40.46872, -40.48458, -40.49953, -40.51381, 
        -40.52814, -40.54245, -40.55725, -40.57256, -40.58825, -40.6041, 
        -40.62005, -40.63591, -40.65171, -40.66662, -40.68116, -40.69558, 
        -40.71051, -40.72626, -40.74226, -40.76024, -40.77869, -40.79776, 
        -40.81698, -40.83685, -40.85793, -40.88052, -40.90495, -40.93233, 
        -40.96118, -40.9915, -41.02232, -41.05245, -41.08122, -41.10838, 
        -41.13342, -41.15665, -41.17811, -41.19812, -41.21697, -41.2349, 
        -41.25111, -41.26514, -41.27703, -41.28587, -41.29115, -41.29449, 
        -41.29543, -41.29503, -41.29446, -41.29417, -41.29499, -41.29679, 
        -41.29955, -41.30301, -41.30681, -41.31078, -41.31462, -41.31835, 
        -41.32186, -41.32566, -41.33032, -41.33648, -41.34447, -41.35423, 
        -41.36513, -41.37607, -41.38745, -41.39859, -41.4091, -41.41927, 
        -41.42919, -41.43944, -41.4502, -41.46198, -41.47335, -41.48637, 
        -41.49941, -41.51289, -41.52673, -41.5408, -41.55501, -41.56926, 
        -41.58326, -41.59706, -41.61063, -41.62406, -41.63707, -41.64981, 
        -41.6623, -41.67487, -41.68779, -41.70117, -41.71511, -41.72934, 
        -41.74371, -41.75824, -41.77252, -41.7859, -41.79765, -41.80717, 
        -41.8142, -41.81918, -41.82301, -41.82648, -41.82984, -41.83276, 
        -41.83483, -41.83573, -41.83538, -41.83371, -41.83085, -41.82535, 
        -41.81992, -41.81241, -41.80326, -41.79201, -41.77873, -41.76264, 
        -41.74377, -41.72179, -41.69687, -41.66987, -41.64183, -41.61317, 
        -41.58408, -41.55387, -41.52209, -41.48664, -41.4465, -41.401, 
        -41.35024, -41.29533, -41.23647, -41.17329, -41.1044, -41.02942, 
        -40.94815, -40.85983, -40.76471, -40.66309, -40.55609, -40.4458, 
        -40.33491,
  -35.88999, -35.92688, -35.965, -36.00463, -36.04574, -36.08806, 
        -36.13031, -36.1743, -36.21866, -36.2631, -36.30712, -36.35032, 
        -36.39246, -36.43359, -36.47387, -36.5134, -36.55239, -36.59088, 
        -36.62879, -36.66599, -36.70243, -36.73768, -36.77369, -36.80954, 
        -36.84543, -36.88134, -36.91691, -36.95199, -36.98634, -37.02003, 
        -37.053, -37.08599, -37.1196, -37.15421, -37.18971, -37.22604, 
        -37.26156, -37.29836, -37.33523, -37.37252, -37.4105, -37.44895, 
        -37.48805, -37.52692, -37.56524, -37.60295, -37.63992, -37.67635, 
        -37.7123, -37.74784, -37.78312, -37.81805, -37.85124, -37.88486, 
        -37.91796, -37.95096, -37.9837, -38.0162, -38.04862, -38.08091, 
        -38.11323, -38.14545, -38.17784, -38.21056, -38.24389, -38.27834, 
        -38.31434, -38.35179, -38.38973, -38.42971, -38.46996, -38.50983, 
        -38.5488, -38.58686, -38.62363, -38.65918, -38.69388, -38.72775, 
        -38.76128, -38.79511, -38.82925, -38.86376, -38.89843, -38.93285, 
        -38.96644, -38.99923, -39.02968, -39.06019, -39.09058, -39.12094, 
        -39.15199, -39.18425, -39.21708, -39.25036, -39.28394, -39.31767, 
        -39.35127, -39.38471, -39.41755, -39.44983, -39.48155, -39.51242, 
        -39.54242, -39.57153, -39.59827, -39.62445, -39.64881, -39.67109, 
        -39.69101, -39.70881, -39.72467, -39.73901, -39.75226, -39.765, 
        -39.7769, -39.78867, -39.7997, -39.80996, -39.81923, -39.82782, 
        -39.83588, -39.84374, -39.85157, -39.85924, -39.86563, -39.87306, 
        -39.88056, -39.88788, -39.89574, -39.90382, -39.91258, -39.9222, 
        -39.93239, -39.94354, -39.95533, -39.96768, -39.98082, -39.99491, 
        -40.01024, -40.0271, -40.0454, -40.06521, -40.08583, -40.10678, 
        -40.12761, -40.14695, -40.16653, -40.18549, -40.20387, -40.22208, 
        -40.24031, -40.25897, -40.27804, -40.2973, -40.31654, -40.33548, 
        -40.35395, -40.37168, -40.38838, -40.40409, -40.41874, -40.43267, 
        -40.44639, -40.46036, -40.47493, -40.49007, -40.5057, -40.52192, 
        -40.53729, -40.5533, -40.5689, -40.58378, -40.59774, -40.61128, 
        -40.6252, -40.64011, -40.6561, -40.67319, -40.69118, -40.71027, 
        -40.72997, -40.7506, -40.77283, -40.79645, -40.8223, -40.85005, 
        -40.87989, -40.91024, -40.94097, -40.9706, -40.99905, -41.02625, 
        -41.05169, -41.07486, -41.09783, -41.11957, -41.14005, -41.15929, 
        -41.17677, -41.19185, -41.20401, -41.21327, -41.21919, -41.22253, 
        -41.22359, -41.22376, -41.22316, -41.2226, -41.22319, -41.22482, 
        -41.22728, -41.23039, -41.23401, -41.2378, -41.24169, -41.24558, 
        -41.24958, -41.25398, -41.2593, -41.26624, -41.27473, -41.28492, 
        -41.29481, -41.30619, -41.31736, -41.32779, -41.33803, -41.34798, 
        -41.35804, -41.36874, -41.38036, -41.39318, -41.40672, -41.42082, 
        -41.43481, -41.44893, -41.46313, -41.47778, -41.49232, -41.50706, 
        -41.52143, -41.53565, -41.54993, -41.56381, -41.57737, -41.5906, 
        -41.60346, -41.61625, -41.62935, -41.64295, -41.65722, -41.672, 
        -41.68707, -41.70219, -41.71708, -41.73121, -41.7426, -41.75261, 
        -41.75986, -41.76484, -41.76851, -41.77187, -41.77534, -41.77851, 
        -41.78092, -41.78243, -41.78275, -41.7819, -41.77969, -41.77598, 
        -41.77113, -41.76432, -41.75557, -41.74438, -41.73082, -41.71522, 
        -41.69644, -41.67491, -41.65098, -41.62498, -41.59792, -41.57048, 
        -41.54244, -41.51316, -41.48171, -41.44696, -41.40776, -41.36314, 
        -41.31326, -41.25871, -41.19976, -41.13625, -41.06704, -40.99168, 
        -40.90988, -40.82083, -40.72432, -40.62041, -40.51041, -40.39618, 
        -40.28086,
  -35.74701, -35.78362, -35.8207, -35.86058, -35.9022, -35.94526, 
        -35.98933, -36.03404, -36.07893, -36.12352, -36.16736, -36.21, 
        -36.25139, -36.29171, -36.33124, -36.37018, -36.40772, -36.44595, 
        -36.48386, -36.52139, -36.55854, -36.59554, -36.63208, -36.66862, 
        -36.70511, -36.7415, -36.77758, -36.81305, -36.84761, -36.88134, 
        -36.91439, -36.94637, -36.98012, -37.01505, -37.05122, -37.08831, 
        -37.1259, -37.1636, -37.2014, -37.23962, -37.27825, -37.31721, 
        -37.35616, -37.39484, -37.43289, -37.47021, -37.50692, -37.54221, 
        -37.57837, -37.6144, -37.65036, -37.68591, -37.72092, -37.75533, 
        -37.78918, -37.82278, -37.85616, -37.88935, -37.92252, -37.95566, 
        -37.9888, -38.02202, -38.0555, -38.0885, -38.12313, -38.15892, 
        -38.19614, -38.23487, -38.27493, -38.31581, -38.35663, -38.39706, 
        -38.43637, -38.47444, -38.51124, -38.54699, -38.58174, -38.61578, 
        -38.64975, -38.68401, -38.71772, -38.75263, -38.78763, -38.82232, 
        -38.85634, -38.88936, -38.9216, -38.95293, -38.98391, -39.01486, 
        -39.04626, -39.0785, -39.11139, -39.14478, -39.17846, -39.21233, 
        -39.24614, -39.27977, -39.31195, -39.34479, -39.37687, -39.40824, 
        -39.43866, -39.46778, -39.49557, -39.5218, -39.54638, -39.56886, 
        -39.58912, -39.60752, -39.62411, -39.63916, -39.6533, -39.66684, 
        -39.68017, -39.69314, -39.70528, -39.71535, -39.72564, -39.73542, 
        -39.74482, -39.75406, -39.76303, -39.77145, -39.77911, -39.78642, 
        -39.79356, -39.80059, -39.80811, -39.81632, -39.82539, -39.83534, 
        -39.84624, -39.85812, -39.87072, -39.88405, -39.89843, -39.91367, 
        -39.92887, -39.94641, -39.96526, -39.98542, -40.00624, -40.02744, 
        -40.04849, -40.06903, -40.08892, -40.10824, -40.12678, -40.14487, 
        -40.16281, -40.18092, -40.19938, -40.21803, -40.23687, -40.2553, 
        -40.27339, -40.29062, -40.3071, -40.32249, -40.33596, -40.34976, 
        -40.36333, -40.3772, -40.39154, -40.40661, -40.42245, -40.43899, 
        -40.45561, -40.47196, -40.48781, -40.50235, -40.51599, -40.52892, 
        -40.54217, -40.5562, -40.57137, -40.5877, -40.60499, -40.62356, 
        -40.64337, -40.66456, -40.68753, -40.71243, -40.73825, -40.76686, 
        -40.79688, -40.82751, -40.85811, -40.88773, -40.91607, -40.94321, 
        -40.96929, -40.99446, -41.01865, -41.04192, -41.06392, -41.08444, 
        -41.10307, -41.11902, -41.13197, -41.14155, -41.1479, -41.15167, 
        -41.15316, -41.15348, -41.15323, -41.15289, -41.15311, -41.15418, 
        -41.15603, -41.1587, -41.16112, -41.16497, -41.16908, -41.17327, 
        -41.17751, -41.18245, -41.1884, -41.1959, -41.20508, -41.21559, 
        -41.22667, -41.23794, -41.24889, -41.25917, -41.26889, -41.27855, 
        -41.28857, -41.2996, -41.31187, -41.32558, -41.34015, -41.35494, 
        -41.36977, -41.38438, -41.39903, -41.41378, -41.42878, -41.44387, 
        -41.4589, -41.47386, -41.48873, -41.50338, -41.51663, -41.53035, 
        -41.54348, -41.55657, -41.56998, -41.58403, -41.59877, -41.61403, 
        -41.62969, -41.64544, -41.661, -41.67574, -41.68885, -41.69944, 
        -41.7071, -41.71217, -41.71568, -41.71874, -41.72193, -41.72506, 
        -41.72776, -41.72974, -41.7307, -41.73065, -41.72935, -41.72661, 
        -41.72229, -41.71616, -41.70801, -41.69735, -41.68406, -41.66818, 
        -41.64978, -41.62886, -41.60569, -41.58095, -41.5551, -41.52877, 
        -41.50161, -41.47316, -41.44119, -41.40698, -41.36821, -41.32473, 
        -41.27593, -41.2222, -41.16343, -41.09962, -41.03029, -40.95453, 
        -40.87217, -40.78228, -40.68429, -40.57805, -40.46469, -40.34626, 
        -40.2258,
  -35.60487, -35.64136, -35.67952, -35.71965, -35.76172, -35.80542, 
        -35.85017, -35.89552, -35.9408, -35.98539, -36.02884, -36.06981, 
        -36.11048, -36.15003, -36.18893, -36.22742, -36.26575, -36.30394, 
        -36.34202, -36.38, -36.41776, -36.45535, -36.49276, -36.52987, 
        -36.5668, -36.60357, -36.63883, -36.6744, -36.70899, -36.74259, 
        -36.77592, -36.80927, -36.84327, -36.87851, -36.91511, -36.95277, 
        -36.99107, -37.02958, -37.06837, -37.10732, -37.14651, -37.18472, 
        -37.22379, -37.26231, -37.30006, -37.33706, -37.37355, -37.40981, 
        -37.44633, -37.48287, -37.51983, -37.55641, -37.59235, -37.62757, 
        -37.66219, -37.69633, -37.73017, -37.76275, -37.79629, -37.83003, 
        -37.86398, -37.89816, -37.93279, -37.96788, -38.00386, -38.04096, 
        -38.07933, -38.1192, -38.16004, -38.20158, -38.24306, -38.28379, 
        -38.32335, -38.36158, -38.39758, -38.43342, -38.46825, -38.50254, 
        -38.53676, -38.57141, -38.60648, -38.64189, -38.6773, -38.71245, 
        -38.74697, -38.78069, -38.81374, -38.84624, -38.87817, -38.90978, 
        -38.94153, -38.97371, -39.00548, -39.039, -39.07282, -39.10685, 
        -39.14108, -39.17494, -39.20843, -39.24197, -39.27459, -39.30631, 
        -39.33677, -39.36568, -39.39339, -39.41937, -39.44383, -39.46657, 
        -39.48735, -39.50658, -39.52423, -39.53924, -39.55434, -39.56917, 
        -39.58345, -39.59709, -39.61003, -39.62181, -39.63276, -39.64346, 
        -39.6543, -39.66488, -39.67509, -39.68438, -39.69259, -39.69981, 
        -39.70655, -39.71341, -39.72078, -39.72901, -39.73831, -39.74751, 
        -39.75864, -39.77077, -39.784, -39.79836, -39.81366, -39.82999, 
        -39.84722, -39.86546, -39.88508, -39.90568, -39.92692, -39.94833, 
        -39.96955, -39.99032, -40.01039, -40.02983, -40.0486, -40.0671, 
        -40.08514, -40.10305, -40.12002, -40.13828, -40.15664, -40.17455, 
        -40.19189, -40.20852, -40.22434, -40.23912, -40.25325, -40.26713, 
        -40.28075, -40.29482, -40.30935, -40.32446, -40.34053, -40.3572, 
        -40.37425, -40.39102, -40.40687, -40.42144, -40.43481, -40.44748, 
        -40.46013, -40.47334, -40.48664, -40.50203, -40.51861, -40.53667, 
        -40.55642, -40.57793, -40.60149, -40.62724, -40.65504, -40.68434, 
        -40.71467, -40.74542, -40.77603, -40.80572, -40.83422, -40.86171, 
        -40.88853, -40.91463, -40.93993, -40.96444, -40.98762, -41.00921, 
        -41.02872, -41.04554, -41.05917, -41.06938, -41.07552, -41.08016, 
        -41.08252, -41.08351, -41.08358, -41.08324, -41.08315, -41.08372, 
        -41.08509, -41.08753, -41.09082, -41.09454, -41.09873, -41.10292, 
        -41.10749, -41.11296, -41.11933, -41.12742, -41.13691, -41.14793, 
        -41.15915, -41.17034, -41.18114, -41.19109, -41.2005, -41.20982, 
        -41.21974, -41.23107, -41.24395, -41.25826, -41.27335, -41.28769, 
        -41.30291, -41.31772, -41.3327, -41.34776, -41.36319, -41.37879, 
        -41.39457, -41.41033, -41.42606, -41.44162, -41.45671, -41.47104, 
        -41.48481, -41.49825, -41.51196, -41.52634, -41.54151, -41.55727, 
        -41.57344, -41.58981, -41.60592, -41.62123, -41.63503, -41.64629, 
        -41.65448, -41.65974, -41.66321, -41.66588, -41.66881, -41.67171, 
        -41.67464, -41.67705, -41.67871, -41.67948, -41.679, -41.67728, 
        -41.67277, -41.66724, -41.65944, -41.64927, -41.63635, -41.62074, 
        -41.60248, -41.58213, -41.56004, -41.53651, -41.51213, -41.48693, 
        -41.46077, -41.43274, -41.4021, -41.36798, -41.33005, -41.28745, 
        -41.24021, -41.18774, -41.12968, -41.06593, -40.99648, -40.92071, 
        -40.83805, -40.74747, -40.64816, -40.53969, -40.42309, -40.30048, 
        -40.17488,
  -35.46586, -35.50256, -35.54088, -35.58125, -35.62358, -35.66758, 
        -35.71278, -35.75747, -35.80291, -35.84733, -35.89031, -35.9317, 
        -35.9717, -36.01071, -36.04918, -36.08745, -36.12564, -36.16393, 
        -36.2022, -36.24045, -36.27864, -36.31575, -36.35376, -36.39141, 
        -36.42865, -36.46537, -36.50177, -36.53744, -36.57226, -36.60615, 
        -36.63965, -36.67359, -36.70833, -36.74362, -36.78061, -36.81866, 
        -36.85646, -36.89567, -36.93521, -36.9748, -37.0146, -37.05432, 
        -37.09342, -37.13176, -37.1691, -37.20584, -37.24224, -37.27888, 
        -37.31573, -37.35323, -37.39103, -37.42862, -37.46443, -37.50052, 
        -37.53585, -37.57056, -37.60479, -37.63874, -37.67268, -37.70689, 
        -37.74147, -37.77641, -37.81188, -37.84795, -37.88502, -37.92325, 
        -37.96269, -38.00327, -38.04484, -38.08592, -38.12797, -38.16911, 
        -38.20907, -38.24756, -38.28475, -38.32079, -38.3559, -38.39058, 
        -38.42503, -38.45984, -38.49542, -38.53126, -38.56718, -38.60286, 
        -38.63803, -38.67273, -38.70583, -38.73944, -38.7724, -38.80481, 
        -38.83695, -38.86929, -38.90202, -38.93527, -38.96917, -39.0032, 
        -39.03738, -39.07207, -39.10591, -39.13941, -39.17262, -39.20477, 
        -39.23549, -39.26458, -39.29105, -39.31701, -39.34159, -39.3647, 
        -39.38597, -39.40618, -39.42459, -39.4416, -39.45765, -39.4731, 
        -39.48815, -39.50212, -39.51535, -39.52764, -39.53925, -39.55079, 
        -39.5626, -39.57429, -39.58548, -39.59562, -39.60337, -39.61105, 
        -39.618, -39.62485, -39.63234, -39.64046, -39.64975, -39.66015, 
        -39.67119, -39.68353, -39.69736, -39.71243, -39.72869, -39.74609, 
        -39.76448, -39.78366, -39.80358, -39.82442, -39.84585, -39.86768, 
        -39.88938, -39.90962, -39.93018, -39.95004, -39.96928, -39.98789, 
        -40.00616, -40.0243, -40.0423, -40.06009, -40.07774, -40.09506, 
        -40.11169, -40.12741, -40.14252, -40.15718, -40.17137, -40.18507, 
        -40.19911, -40.21337, -40.22809, -40.24355, -40.25975, -40.27658, 
        -40.2928, -40.30966, -40.3258, -40.3405, -40.35355, -40.36586, 
        -40.37799, -40.39045, -40.40409, -40.41854, -40.43431, -40.452, 
        -40.47165, -40.49353, -40.51788, -40.54436, -40.5729, -40.60275, 
        -40.63348, -40.66461, -40.69522, -40.7251, -40.75393, -40.78195, 
        -40.80934, -40.83506, -40.86109, -40.88616, -40.90998, -40.93228, 
        -40.95254, -40.97034, -40.98506, -40.99643, -41.00468, -41.0103, 
        -41.01332, -41.01501, -41.01547, -41.01539, -41.01524, -41.01556, 
        -41.01651, -41.01867, -41.02172, -41.02529, -41.02945, -41.03395, 
        -41.03878, -41.04444, -41.05121, -41.05986, -41.06968, -41.08053, 
        -41.0905, -41.10161, -41.11228, -41.12192, -41.13146, -41.14079, 
        -41.15109, -41.16261, -41.17583, -41.19045, -41.20583, -41.22143, 
        -41.23675, -41.25178, -41.26683, -41.2822, -41.29805, -41.31439, 
        -41.33097, -41.34779, -41.36458, -41.3812, -41.39716, -41.41212, 
        -41.42636, -41.44021, -41.45419, -41.46887, -41.48442, -41.50069, 
        -41.51738, -41.53415, -41.5507, -41.5665, -41.58076, -41.59152, 
        -41.60027, -41.60569, -41.60918, -41.6119, -41.61446, -41.61734, 
        -41.62032, -41.6232, -41.62572, -41.62736, -41.62801, -41.62753, 
        -41.62447, -41.61941, -41.61237, -41.60259, -41.59014, -41.57486, 
        -41.55709, -41.53735, -41.51629, -41.49408, -41.47107, -41.44727, 
        -41.42195, -41.39455, -41.36418, -41.33017, -41.2926, -41.25085, 
        -41.20484, -41.15361, -41.09686, -41.03374, -40.96461, -40.88932, 
        -40.80683, -40.71601, -40.61592, -40.50575, -40.38648, -40.26012, 
        -40.12994,
  -35.32919, -35.36631, -35.40389, -35.44434, -35.48664, -35.53077, 
        -35.57604, -35.62175, -35.66704, -35.71115, -35.75359, -35.79444, 
        -35.83402, -35.87275, -35.91105, -35.94937, -35.98672, -36.02507, 
        -36.06353, -36.10192, -36.14029, -36.17868, -36.21691, -36.25492, 
        -36.29239, -36.32951, -36.36618, -36.40197, -36.43699, -36.47145, 
        -36.50572, -36.53931, -36.57449, -36.61025, -36.64726, -36.68549, 
        -36.72446, -36.76413, -36.80415, -36.84447, -36.88503, -36.92513, 
        -36.96433, -37.00249, -37.0398, -37.07647, -37.11299, -37.14888, 
        -37.18638, -37.22491, -37.26347, -37.30184, -37.33973, -37.37663, 
        -37.4126, -37.44773, -37.48227, -37.51648, -37.55061, -37.58524, 
        -37.62038, -37.65594, -37.69211, -37.72814, -37.76606, -37.8051, 
        -37.84523, -37.88648, -37.92857, -37.9712, -38.01356, -38.05513, 
        -38.09553, -38.13449, -38.17213, -38.20865, -38.24417, -38.27922, 
        -38.31401, -38.34937, -38.38429, -38.42053, -38.45704, -38.49324, 
        -38.52914, -38.56471, -38.59977, -38.63447, -38.66839, -38.70158, 
        -38.73423, -38.76677, -38.79962, -38.83289, -38.86676, -38.90091, 
        -38.9351, -38.96952, -39.00294, -39.03704, -39.07068, -39.1034, 
        -39.13426, -39.16343, -39.19091, -39.21711, -39.2419, -39.26531, 
        -39.28738, -39.30823, -39.32745, -39.34543, -39.36214, -39.37817, 
        -39.39343, -39.40789, -39.42134, -39.43291, -39.44479, -39.45689, 
        -39.46919, -39.48149, -39.49335, -39.50414, -39.5137, -39.52209, 
        -39.52967, -39.53699, -39.54465, -39.55309, -39.56255, -39.57307, 
        -39.58454, -39.59703, -39.61136, -39.62707, -39.64424, -39.66262, 
        -39.68069, -39.70044, -39.72086, -39.74194, -39.76339, -39.78538, 
        -39.80742, -39.82911, -39.85041, -39.87103, -39.89091, -39.90995, 
        -39.92803, -39.94587, -39.9636, -39.98116, -39.99837, -40.01522, 
        -40.03138, -40.0467, -40.06123, -40.07561, -40.08875, -40.1029, 
        -40.1174, -40.1321, -40.14719, -40.16283, -40.17923, -40.19625, 
        -40.21336, -40.23045, -40.24657, -40.26125, -40.27462, -40.28677, 
        -40.2986, -40.31049, -40.32334, -40.33704, -40.35249, -40.36986, 
        -40.38964, -40.41197, -40.4369, -40.46437, -40.49355, -40.52258, 
        -40.55353, -40.58469, -40.61517, -40.64502, -40.6743, -40.70287, 
        -40.73054, -40.7577, -40.78405, -40.80941, -40.8334, -40.85619, 
        -40.87719, -40.89575, -40.91137, -40.92374, -40.9331, -40.93972, 
        -40.94411, -40.94673, -40.94788, -40.94804, -40.94807, -40.94821, 
        -40.94894, -40.95081, -40.95259, -40.95599, -40.96003, -40.96455, 
        -40.96971, -40.97575, -40.98292, -40.99137, -41.00088, -41.01151, 
        -41.0224, -41.03289, -41.04374, -41.05376, -41.06338, -41.07333, 
        -41.08415, -41.09609, -41.10962, -41.12432, -41.13979, -41.15539, 
        -41.17059, -41.18558, -41.20071, -41.2164, -41.23289, -41.25014, 
        -41.26786, -41.28584, -41.30381, -41.32141, -41.33725, -41.35276, 
        -41.36744, -41.38151, -41.39577, -41.41072, -41.42654, -41.44307, 
        -41.46005, -41.47717, -41.49398, -41.51004, -41.52463, -41.53687, 
        -41.54605, -41.55217, -41.55611, -41.55875, -41.56133, -41.56424, 
        -41.56736, -41.57063, -41.57386, -41.57667, -41.57827, -41.57829, 
        -41.57618, -41.57203, -41.56527, -41.5559, -41.54426, -41.52938, 
        -41.51237, -41.49335, -41.47322, -41.45247, -41.43111, -41.40886, 
        -41.38451, -41.35751, -41.3274, -41.29278, -41.25546, -41.21439, 
        -41.16926, -41.11947, -41.06395, -41.00198, -40.93364, -40.85936, 
        -40.77765, -40.68719, -40.58699, -40.47607, -40.35513, -40.22596, 
        -40.09216,
  -35.1935, -35.23123, -35.27015, -35.31063, -35.3529, -35.39676, 
        -35.44179, -35.48727, -35.5323, -35.57598, -35.61797, -35.65744, 
        -35.69681, -35.73552, -35.77396, -35.81239, -35.85094, -35.88945, 
        -35.92789, -35.96618, -36.00459, -36.04293, -36.08117, -36.11929, 
        -36.1571, -36.19452, -36.23049, -36.26682, -36.30247, -36.33776, 
        -36.37305, -36.40866, -36.44423, -36.48036, -36.51723, -36.55514, 
        -36.59417, -36.63427, -36.67493, -36.71594, -36.75691, -36.79731, 
        -36.83578, -36.87398, -36.91135, -36.94827, -36.98518, -37.02253, 
        -37.06064, -37.09959, -37.13893, -37.17811, -37.21669, -37.25437, 
        -37.29104, -37.3266, -37.36147, -37.39595, -37.42945, -37.46437, 
        -37.49982, -37.53586, -37.57257, -37.61008, -37.64852, -37.68813, 
        -37.72888, -37.7708, -37.81331, -37.85605, -37.89876, -37.94097, 
        -37.98199, -38.02159, -38.05978, -38.09578, -38.132, -38.16774, 
        -38.20343, -38.23944, -38.27539, -38.31203, -38.34894, -38.38608, 
        -38.42273, -38.45906, -38.49517, -38.5307, -38.56542, -38.59929, 
        -38.63252, -38.66537, -38.69735, -38.73069, -38.76435, -38.79841, 
        -38.83274, -38.86726, -38.90196, -38.93665, -38.97073, -39.00384, 
        -39.03518, -39.0646, -39.09227, -39.11854, -39.14367, -39.16777, 
        -39.19049, -39.21183, -39.23181, -39.2493, -39.26665, -39.28309, 
        -39.2988, -39.31329, -39.3269, -39.3395, -39.35173, -39.36391, 
        -39.37656, -39.38919, -39.40142, -39.41274, -39.42293, -39.43207, 
        -39.44051, -39.4486, -39.45686, -39.46581, -39.47547, -39.48505, 
        -39.49664, -39.50959, -39.52418, -39.54059, -39.55873, -39.57794, 
        -39.59788, -39.61829, -39.63909, -39.6604, -39.68202, -39.70398, 
        -39.72626, -39.74824, -39.77007, -39.79128, -39.8116, -39.83091, 
        -39.84941, -39.86733, -39.88476, -39.90091, -39.9175, -39.93375, 
        -39.94977, -39.96503, -39.97963, -39.99413, -40.00846, -40.02291, 
        -40.03766, -40.05274, -40.06817, -40.08405, -40.10067, -40.11771, 
        -40.13495, -40.15209, -40.16837, -40.18324, -40.19666, -40.20893, 
        -40.22046, -40.232, -40.24326, -40.25665, -40.272, -40.2896, 
        -40.30979, -40.33268, -40.35834, -40.38625, -40.41555, -40.44606, 
        -40.47709, -40.50794, -40.53829, -40.56818, -40.59738, -40.62638, 
        -40.65452, -40.68188, -40.70834, -40.7337, -40.75776, -40.78045, 
        -40.8017, -40.82085, -40.83743, -40.85091, -40.86165, -40.86823, 
        -40.87365, -40.87727, -40.87925, -40.88001, -40.88033, -40.8805, 
        -40.88116, -40.88255, -40.88501, -40.88824, -40.89212, -40.89664, 
        -40.90193, -40.90813, -40.91536, -40.92366, -40.93291, -40.9429, 
        -40.9534, -40.96392, -40.97437, -40.98496, -40.99531, -41.00609, 
        -41.01766, -41.03031, -41.04408, -41.05878, -41.07415, -41.08853, 
        -41.1037, -41.11875, -41.13402, -41.15018, -41.16743, -41.18576, 
        -41.20471, -41.22406, -41.24325, -41.26175, -41.27911, -41.29512, 
        -41.31012, -41.32433, -41.33871, -41.35378, -41.36973, -41.38638, 
        -41.40345, -41.42057, -41.43739, -41.45346, -41.46819, -41.48092, 
        -41.49079, -41.4978, -41.50236, -41.50547, -41.50828, -41.51133, 
        -41.51473, -41.51844, -41.52239, -41.526, -41.52857, -41.5294, 
        -41.52699, -41.52325, -41.51714, -41.50869, -41.49728, -41.48337, 
        -41.4671, -41.44912, -41.43023, -41.41099, -41.39127, -41.37036, 
        -41.34729, -41.32089, -41.29111, -41.25801, -41.22141, -41.18095, 
        -41.13656, -41.08763, -41.03323, -40.97268, -40.90563, -40.83247, 
        -40.75188, -40.66247, -40.56319, -40.45258, -40.33116, -40.20086, 
        -40.06511,
  -35.06044, -35.0989, -35.1382, -35.17879, -35.22089, -35.26444, 
        -35.30912, -35.35318, -35.39771, -35.44093, -35.4826, -35.52293, 
        -35.56234, -35.60126, -35.63997, -35.67859, -35.71718, -35.75563, 
        -35.79401, -35.83208, -35.87018, -35.90726, -35.94536, -35.98351, 
        -36.02149, -36.05927, -36.09672, -36.1339, -36.17057, -36.20723, 
        -36.24378, -36.28025, -36.31659, -36.35279, -36.38942, -36.42696, 
        -36.46621, -36.50559, -36.54681, -36.58841, -36.62991, -36.67061, 
        -36.71014, -36.74859, -36.78619, -36.82342, -36.86077, -36.8986, 
        -36.93721, -36.97655, -37.01644, -37.05612, -37.09434, -37.13264, 
        -37.16998, -37.20618, -37.24145, -37.27622, -37.31096, -37.34602, 
        -37.38165, -37.41795, -37.45499, -37.49286, -37.53175, -37.57182, 
        -37.61313, -37.65535, -37.69815, -37.74022, -37.78325, -37.82573, 
        -37.86741, -37.9076, -37.94643, -37.98422, -38.02128, -38.05805, 
        -38.09444, -38.1311, -38.16832, -38.20529, -38.24277, -38.28049, 
        -38.31807, -38.35508, -38.39108, -38.42733, -38.46276, -38.49715, 
        -38.53075, -38.56395, -38.59722, -38.63054, -38.66417, -38.69804, 
        -38.73222, -38.76675, -38.80185, -38.83693, -38.87157, -38.90521, 
        -38.93707, -38.96685, -38.99489, -39.02062, -39.04633, -39.07079, 
        -39.0941, -39.11587, -39.13618, -39.15482, -39.17277, -39.18956, 
        -39.20531, -39.22059, -39.23432, -39.24705, -39.25937, -39.27179, 
        -39.28442, -39.29704, -39.30941, -39.32104, -39.3307, -39.34069, 
        -39.34998, -39.35877, -39.36783, -39.37725, -39.38735, -39.39808, 
        -39.40988, -39.42303, -39.4381, -39.45515, -39.47401, -39.49412, 
        -39.51487, -39.53596, -39.55723, -39.57862, -39.6005, -39.6226, 
        -39.64502, -39.66635, -39.68864, -39.71023, -39.73095, -39.75074, 
        -39.76949, -39.78754, -39.80487, -39.82158, -39.83795, -39.85389, 
        -39.86964, -39.88493, -39.89968, -39.91425, -39.92897, -39.94372, 
        -39.95885, -39.97422, -39.98983, -40.00608, -40.02275, -40.04007, 
        -40.0565, -40.07359, -40.0896, -40.10461, -40.11813, -40.13053, 
        -40.14227, -40.15379, -40.1659, -40.17967, -40.19524, -40.21337, 
        -40.23405, -40.25756, -40.28374, -40.31206, -40.3419, -40.37266, 
        -40.40384, -40.4344, -40.46434, -40.49396, -40.5233, -40.55217, 
        -40.58048, -40.60794, -40.63342, -40.65866, -40.68256, -40.70515, 
        -40.72625, -40.74566, -40.76276, -40.77709, -40.78874, -40.79776, 
        -40.80431, -40.80882, -40.81161, -40.81306, -40.81365, -40.81393, 
        -40.81458, -40.81599, -40.81797, -40.82067, -40.82426, -40.82867, 
        -40.83391, -40.84032, -40.84748, -40.85569, -40.86462, -40.87415, 
        -40.88395, -40.8932, -40.90371, -40.91454, -40.92567, -40.93756, 
        -40.95018, -40.96362, -40.97796, -40.99284, -41.00811, -41.02338, 
        -41.03849, -41.05362, -41.06937, -41.08609, -41.10429, -41.12376, 
        -41.1441, -41.16483, -41.18506, -41.20433, -41.22211, -41.23832, 
        -41.25351, -41.26777, -41.28225, -41.29727, -41.31311, -41.32972, 
        -41.34663, -41.36346, -41.37991, -41.39561, -41.41031, -41.42235, 
        -41.43306, -41.4411, -41.44666, -41.45074, -41.45408, -41.45772, 
        -41.46151, -41.46587, -41.47031, -41.47451, -41.47781, -41.47931, 
        -41.47855, -41.47546, -41.4701, -41.46244, -41.45193, -41.43894, 
        -41.42376, -41.40689, -41.3895, -41.37181, -41.35359, -41.33389, 
        -41.31176, -41.28651, -41.25729, -41.22497, -41.18935, -41.14968, 
        -41.10601, -41.05796, -41.00426, -40.94489, -40.87934, -40.80745, 
        -40.72818, -40.64046, -40.54262, -40.4335, -40.31305, -40.18311, 
        -40.04703,
  -34.92884, -34.96783, -35.00653, -35.0473, -35.08937, -35.13275, 
        -35.17707, -35.2214, -35.26542, -35.30822, -35.34977, -35.39032, 
        -35.42993, -35.46926, -35.50809, -35.54666, -35.58512, -35.62236, 
        -35.66037, -35.69826, -35.73593, -35.77369, -35.81161, -35.84958, 
        -35.88776, -35.9258, -35.96402, -36.00213, -36.04047, -36.07877, 
        -36.11666, -36.15316, -36.19008, -36.22625, -36.26284, -36.30046, 
        -36.33961, -36.38038, -36.4221, -36.46403, -36.50569, -36.54659, 
        -36.5864, -36.62516, -36.6632, -36.70087, -36.73875, -36.77603, 
        -36.81491, -36.85457, -36.89475, -36.93489, -36.97455, -37.01351, 
        -37.05129, -37.08797, -37.12366, -37.15886, -37.19386, -37.22904, 
        -37.26474, -37.30119, -37.33837, -37.37562, -37.41495, -37.45558, 
        -37.49728, -37.53978, -37.58264, -37.62574, -37.66893, -37.71175, 
        -37.7538, -37.79457, -37.83409, -37.87291, -37.91101, -37.94882, 
        -37.98629, -38.02395, -38.06182, -38.09896, -38.1372, -38.17568, 
        -38.21415, -38.25214, -38.28976, -38.32663, -38.36237, -38.3971, 
        -38.4311, -38.46468, -38.49821, -38.5316, -38.56507, -38.59875, 
        -38.63298, -38.66772, -38.70305, -38.73762, -38.7729, -38.8067, 
        -38.83871, -38.86879, -38.89708, -38.92425, -38.95034, -38.97538, 
        -38.99912, -39.02122, -39.04193, -39.06118, -39.0793, -39.09652, 
        -39.11278, -39.12815, -39.14231, -39.15524, -39.16684, -39.17937, 
        -39.19188, -39.20458, -39.2168, -39.22868, -39.23985, -39.25026, 
        -39.26046, -39.27027, -39.28014, -39.28996, -39.30033, -39.31128, 
        -39.32324, -39.33688, -39.35245, -39.37017, -39.38982, -39.41073, 
        -39.43124, -39.45295, -39.47475, -39.49649, -39.51862, -39.54091, 
        -39.56349, -39.58629, -39.60875, -39.63077, -39.65187, -39.67185, 
        -39.69074, -39.70877, -39.726, -39.74271, -39.75889, -39.7747, 
        -39.79016, -39.80537, -39.8204, -39.83524, -39.85001, -39.86399, 
        -39.87934, -39.89504, -39.91132, -39.92799, -39.94501, -39.96247, 
        -39.97982, -39.99663, -40.01252, -40.02741, -40.0411, -40.05366, 
        -40.06567, -40.07769, -40.0905, -40.10479, -40.12124, -40.1398, 
        -40.16135, -40.18547, -40.21235, -40.24117, -40.27148, -40.30121, 
        -40.33197, -40.36238, -40.39238, -40.42193, -40.45103, -40.47967, 
        -40.50786, -40.53535, -40.56163, -40.58678, -40.61056, -40.63276, 
        -40.65355, -40.6728, -40.68998, -40.70486, -40.71737, -40.72717, 
        -40.73482, -40.74046, -40.74426, -40.74643, -40.7474, -40.74784, 
        -40.74842, -40.7495, -40.75104, -40.75212, -40.75516, -40.75911, 
        -40.76449, -40.77094, -40.77842, -40.78644, -40.79528, -40.80427, 
        -40.81358, -40.82319, -40.8334, -40.84456, -40.8567, -40.86975, 
        -40.88355, -40.89801, -40.91308, -40.92837, -40.94367, -40.95903, 
        -40.97427, -40.98984, -41.00621, -41.02389, -41.04308, -41.06358, 
        -41.08481, -41.10662, -41.12778, -41.14762, -41.16572, -41.18124, 
        -41.19655, -41.21102, -41.22551, -41.24051, -41.25615, -41.27241, 
        -41.2889, -41.3052, -41.32098, -41.33617, -41.35065, -41.36391, 
        -41.37536, -41.38454, -41.39134, -41.39663, -41.40103, -41.4054, 
        -41.40995, -41.41481, -41.41984, -41.42432, -41.42799, -41.42989, 
        -41.42974, -41.42741, -41.42295, -41.41624, -41.40697, -41.39513, 
        -41.3811, -41.36567, -41.34966, -41.33363, -41.31671, -41.29816, 
        -41.27707, -41.25266, -41.22483, -41.19264, -41.15802, -41.11961, 
        -41.07663, -41.02894, -40.97592, -40.91743, -40.85328, -40.78267, 
        -40.70523, -40.61939, -40.52372, -40.4169, -40.29867, -40.17058, 
        -40.03605,
  -34.79742, -34.83693, -34.877, -34.9181, -34.96024, -35.00342, 
        -35.04733, -35.09104, -35.13438, -35.17673, -35.21819, -35.25888, 
        -35.29806, -35.33751, -35.37657, -35.41516, -35.45332, -35.49112, 
        -35.52878, -35.56633, -35.60395, -35.64146, -35.67901, -35.71704, 
        -35.75532, -35.79373, -35.83305, -35.87179, -35.91159, -35.95116, 
        -35.99086, -36.02929, -36.06668, -36.1032, -36.13985, -36.17722, 
        -36.21667, -36.2575, -36.29935, -36.34134, -36.38307, -36.42411, 
        -36.46322, -36.50241, -36.54091, -36.57915, -36.6174, -36.65602, 
        -36.69537, -36.73549, -36.77608, -36.81659, -36.8567, -36.89598, 
        -36.93409, -36.97114, -37.00717, -37.04269, -37.07706, -37.11243, 
        -37.14835, -37.18489, -37.22232, -37.2608, -37.30071, -37.3418, 
        -37.38388, -37.42657, -37.46946, -37.51237, -37.55534, -37.59834, 
        -37.64056, -37.68179, -37.72226, -37.76097, -37.80012, -37.83894, 
        -37.87753, -37.91626, -37.95508, -37.99426, -38.03365, -38.07321, 
        -38.11274, -38.15166, -38.18995, -38.22715, -38.26322, -38.29823, 
        -38.33245, -38.36636, -38.40014, -38.43296, -38.46676, -38.50072, 
        -38.53503, -38.57031, -38.60621, -38.64211, -38.67737, -38.71106, 
        -38.74306, -38.77297, -38.80112, -38.82819, -38.85452, -38.87967, 
        -38.90371, -38.9262, -38.94728, -38.96598, -38.98466, -39.00239, 
        -39.01923, -39.03505, -39.04933, -39.06286, -39.07571, -39.08823, 
        -39.10077, -39.11315, -39.1255, -39.13757, -39.14942, -39.16078, 
        -39.17188, -39.18249, -39.19306, -39.20347, -39.21402, -39.22449, 
        -39.23674, -39.25085, -39.26699, -39.28547, -39.30603, -39.32768, 
        -39.34984, -39.37217, -39.39442, -39.41683, -39.43939, -39.46197, 
        -39.48475, -39.50779, -39.53056, -39.55285, -39.57396, -39.59396, 
        -39.6127, -39.63057, -39.64761, -39.66308, -39.67909, -39.69477, 
        -39.71029, -39.7257, -39.74089, -39.75591, -39.77105, -39.78627, 
        -39.80175, -39.81792, -39.8343, -39.85133, -39.86854, -39.88598, 
        -39.90283, -39.91949, -39.93538, -39.95031, -39.96419, -39.9775, 
        -39.99054, -40.00368, -40.01758, -40.03217, -40.0497, -40.0697, 
        -40.09197, -40.11682, -40.14417, -40.17302, -40.2033, -40.23378, 
        -40.26442, -40.29447, -40.32401, -40.3532, -40.38208, -40.41066, 
        -40.43882, -40.46632, -40.49246, -40.51704, -40.54037, -40.56216, 
        -40.58248, -40.60125, -40.61834, -40.63345, -40.64651, -40.65634, 
        -40.66492, -40.67139, -40.67588, -40.6787, -40.68017, -40.6808, 
        -40.68135, -40.68205, -40.68301, -40.68457, -40.6869, -40.69053, 
        -40.69567, -40.70228, -40.71007, -40.7182, -40.72696, -40.73506, 
        -40.74373, -40.75296, -40.76317, -40.77465, -40.78747, -40.80149, 
        -40.81643, -40.83201, -40.84792, -40.86382, -40.87959, -40.89531, 
        -40.91014, -40.92639, -40.94374, -40.96242, -40.98293, -41.00426, 
        -41.02655, -41.04901, -41.07056, -41.09069, -41.10903, -41.12572, 
        -41.14121, -41.15599, -41.17065, -41.1856, -41.20111, -41.21693, 
        -41.23289, -41.24848, -41.26354, -41.27802, -41.29211, -41.30545, 
        -41.31755, -41.32779, -41.33604, -41.34275, -41.34877, -41.35432, 
        -41.35964, -41.36511, -41.37027, -41.37484, -41.37831, -41.38049, 
        -41.38067, -41.37779, -41.37438, -41.36885, -41.36097, -41.35066, 
        -41.33813, -41.32419, -41.30959, -41.2947, -41.27906, -41.26159, 
        -41.24158, -41.21846, -41.19197, -41.16211, -41.12868, -41.09134, 
        -41.04928, -41.00222, -40.94979, -40.89212, -40.8291, -40.76028, 
        -40.68445, -40.60057, -40.50731, -40.40313, -40.28799, -40.16285, 
        -40.03085,
  -34.66794, -34.70795, -34.74844, -34.78991, -34.83246, -34.87551, 
        -34.91888, -34.96124, -35.00364, -35.04559, -35.08703, -35.12791, 
        -35.16833, -35.20812, -35.24718, -35.28549, -35.32324, -35.36064, 
        -35.3979, -35.43516, -35.47242, -35.50993, -35.54673, -35.58489, 
        -35.62362, -35.66306, -35.70331, -35.74415, -35.7857, -35.82708, 
        -35.86781, -35.90725, -35.94513, -35.98185, -36.01848, -36.05618, 
        -36.0955, -36.13541, -36.17714, -36.21911, -36.26067, -36.30175, 
        -36.34221, -36.38197, -36.4211, -36.45985, -36.49858, -36.53758, 
        -36.5774, -36.61759, -36.65853, -36.69945, -36.73995, -36.77853, 
        -36.8169, -36.85414, -36.89059, -36.92665, -36.96261, -36.99845, 
        -37.03477, -37.07152, -37.10917, -37.14809, -37.18837, -37.22989, 
        -37.27228, -37.31504, -37.35776, -37.39941, -37.44214, -37.48483, 
        -37.52722, -37.56901, -37.61018, -37.65081, -37.69107, -37.73091, 
        -37.77052, -37.8103, -37.8503, -37.89068, -37.93122, -37.9721, 
        -38.0125, -38.05231, -38.09112, -38.12774, -38.16397, -38.19913, 
        -38.23365, -38.26787, -38.30213, -38.33656, -38.37091, -38.40548, 
        -38.44028, -38.47596, -38.51221, -38.54833, -38.58336, -38.61683, 
        -38.64828, -38.67759, -38.70538, -38.73132, -38.75733, -38.78275, 
        -38.80687, -38.82972, -38.85129, -38.87183, -38.89129, -38.90973, 
        -38.92718, -38.94329, -38.95823, -38.97212, -38.98521, -38.99768, 
        -39.01009, -39.02232, -39.03461, -39.04704, -39.05956, -39.07085, 
        -39.08297, -39.09452, -39.10566, -39.1164, -39.12754, -39.13916, 
        -39.15212, -39.16664, -39.18338, -39.20266, -39.22398, -39.24626, 
        -39.26897, -39.29193, -39.3148, -39.33786, -39.36094, -39.38422, 
        -39.40752, -39.43079, -39.45276, -39.47509, -39.49635, -39.51608, 
        -39.53449, -39.55177, -39.56844, -39.58453, -39.6003, -39.61592, 
        -39.63161, -39.6473, -39.66285, -39.67834, -39.69387, -39.70938, 
        -39.72535, -39.74163, -39.75832, -39.77537, -39.79261, -39.80959, 
        -39.82629, -39.84167, -39.85728, -39.87209, -39.88655, -39.9006, 
        -39.91503, -39.92994, -39.94576, -39.96326, -39.98256, -40.00385, 
        -40.02748, -40.05297, -40.08041, -40.10917, -40.13918, -40.16936, 
        -40.19942, -40.22915, -40.25815, -40.28679, -40.31522, -40.34352, 
        -40.37152, -40.39885, -40.42389, -40.44842, -40.47125, -40.49249, 
        -40.51205, -40.53023, -40.54684, -40.56206, -40.57541, -40.58698, 
        -40.59634, -40.6037, -40.609, -40.61238, -40.61423, -40.61515, 
        -40.61562, -40.61604, -40.61657, -40.61737, -40.61909, -40.62233, 
        -40.62734, -40.63393, -40.64156, -40.64999, -40.65808, -40.6662, 
        -40.67461, -40.68225, -40.6922, -40.7039, -40.71706, -40.73188, 
        -40.74786, -40.76455, -40.7815, -40.79841, -40.81499, -40.83149, 
        -40.84818, -40.86569, -40.88422, -40.90417, -40.92566, -40.94819, 
        -40.97116, -40.99384, -41.01551, -41.0356, -41.05395, -41.07069, 
        -41.08649, -41.10174, -41.11669, -41.13174, -41.14706, -41.16269, 
        -41.17794, -41.19289, -41.20732, -41.22111, -41.23481, -41.24814, 
        -41.25976, -41.27091, -41.28043, -41.28842, -41.29587, -41.30264, 
        -41.30896, -41.31483, -41.32002, -41.32433, -41.32776, -41.32977, 
        -41.33026, -41.32929, -41.32674, -41.32262, -41.31646, -41.30781, 
        -41.29693, -41.28445, -41.27112, -41.25726, -41.24265, -41.22629, 
        -41.20736, -41.18545, -41.16034, -41.132, -41.10003, -41.06382, 
        -41.02288, -40.97649, -40.92459, -40.86753, -40.80547, -40.73792, 
        -40.66379, -40.58171, -40.49073, -40.38977, -40.278, -40.1567, 
        -40.02849,
  -34.53925, -34.57968, -34.61969, -34.66164, -34.70456, -34.74773, 
        -34.79065, -34.83325, -34.87513, -34.91667, -34.95792, -34.99892, 
        -35.03947, -35.07933, -35.11829, -35.1563, -35.19359, -35.22952, 
        -35.26639, -35.30347, -35.34082, -35.37861, -35.41679, -35.45551, 
        -35.49503, -35.53551, -35.57696, -35.6193, -35.66214, -35.70474, 
        -35.74618, -35.78627, -35.82359, -35.86052, -35.89716, -35.93516, 
        -35.97456, -36.0153, -36.0568, -36.09845, -36.13993, -36.18117, 
        -36.2221, -36.26251, -36.30228, -36.34153, -36.38059, -36.419, 
        -36.45895, -36.49938, -36.54054, -36.58192, -36.62283, -36.66264, 
        -36.70119, -36.7387, -36.77564, -36.81235, -36.84908, -36.88578, 
        -36.92268, -36.9599, -36.998, -37.03735, -37.07704, -37.11892, 
        -37.16143, -37.20405, -37.24644, -37.28877, -37.33116, -37.37366, 
        -37.41624, -37.45861, -37.50056, -37.54206, -37.58315, -37.62392, 
        -37.66458, -37.70542, -37.74668, -37.78735, -37.82922, -37.871, 
        -37.91234, -37.95281, -37.99215, -38.02992, -38.06631, -38.10164, 
        -38.13643, -38.17125, -38.20598, -38.24096, -38.27603, -38.3115, 
        -38.34735, -38.38359, -38.42008, -38.45512, -38.48995, -38.52278, 
        -38.55336, -38.5819, -38.60912, -38.63579, -38.66163, -38.68678, 
        -38.71121, -38.73459, -38.75673, -38.77813, -38.79872, -38.81803, 
        -38.83619, -38.85291, -38.86811, -38.88222, -38.89453, -38.90705, 
        -38.91922, -38.9314, -38.94385, -38.95669, -38.96987, -38.98326, 
        -38.9963, -39.00884, -39.02052, -39.03178, -39.04306, -39.05499, 
        -39.06817, -39.08331, -39.10081, -39.12074, -39.14254, -39.16541, 
        -39.18868, -39.21125, -39.2348, -39.25851, -39.28244, -39.30639, 
        -39.33037, -39.35411, -39.37735, -39.39978, -39.42071, -39.44017, 
        -39.45808, -39.47464, -39.49061, -39.50611, -39.52164, -39.53736, 
        -39.55341, -39.56949, -39.58557, -39.60155, -39.61763, -39.63259, 
        -39.64869, -39.66511, -39.682, -39.69905, -39.7162, -39.73286, 
        -39.74921, -39.76523, -39.78063, -39.79584, -39.81087, -39.82608, 
        -39.84187, -39.8588, -39.87679, -39.8964, -39.91768, -39.94055, 
        -39.96487, -39.99114, -40.01874, -40.04743, -40.07671, -40.10649, 
        -40.13483, -40.16393, -40.19244, -40.22048, -40.24854, -40.27659, 
        -40.30435, -40.33142, -40.35744, -40.38193, -40.40461, -40.42533, 
        -40.44428, -40.46175, -40.47803, -40.49293, -40.50656, -40.51856, 
        -40.52867, -40.53685, -40.54293, -40.54694, -40.54921, -40.55018, 
        -40.5506, -40.55071, -40.55077, -40.55014, -40.55136, -40.55424, 
        -40.55898, -40.5654, -40.5729, -40.58088, -40.58887, -40.59659, 
        -40.6045, -40.61325, -40.62271, -40.63434, -40.64779, -40.66318, 
        -40.68002, -40.69786, -40.71602, -40.73413, -40.75192, -40.76962, 
        -40.78751, -40.80629, -40.82653, -40.84783, -40.87037, -40.89377, 
        -40.91724, -40.94, -40.96151, -40.98129, -40.9996, -41.0155, 
        -41.03154, -41.04714, -41.06251, -41.0778, -41.09306, -41.10834, 
        -41.12337, -41.13797, -41.15169, -41.16503, -41.17834, -41.1915, 
        -41.20423, -41.21601, -41.22669, -41.23611, -41.24475, -41.25258, 
        -41.25959, -41.26567, -41.27069, -41.27473, -41.27779, -41.27976, 
        -41.28061, -41.28086, -41.27975, -41.2771, -41.27251, -41.26556, 
        -41.25634, -41.24527, -41.23314, -41.22031, -41.20652, -41.19119, 
        -41.17341, -41.15263, -41.12911, -41.10212, -41.07039, -41.03561, 
        -40.99541, -40.94977, -40.89834, -40.84156, -40.78008, -40.71359, 
        -40.64096, -40.56064, -40.4719, -40.37383, -40.26591, -40.14867, 
        -40.02479,
  -34.41016, -34.45107, -34.49259, -34.53501, -34.57811, -34.6213, 
        -34.66412, -34.70624, -34.74768, -34.7888, -34.82979, -34.87064, 
        -34.91009, -34.94972, -34.98858, -35.02633, -35.0634, -35.10011, 
        -35.1369, -35.17399, -35.21159, -35.24982, -35.28876, -35.32848, 
        -35.36913, -35.41087, -35.45361, -35.49611, -35.54002, -35.58335, 
        -35.62537, -35.66557, -35.70392, -35.74107, -35.77794, -35.81581, 
        -35.85513, -35.89563, -35.93677, -35.9782, -36.01964, -36.06113, 
        -36.10165, -36.14283, -36.18335, -36.22306, -36.26244, -36.30186, 
        -36.34201, -36.3828, -36.42426, -36.46588, -36.5071, -36.54714, 
        -36.5859, -36.6237, -36.66122, -36.69876, -36.73549, -36.77318, 
        -36.81089, -36.84891, -36.88759, -36.92739, -36.96851, -37.01057, 
        -37.05311, -37.09555, -37.13758, -37.17965, -37.22189, -37.26448, 
        -37.30735, -37.35038, -37.3931, -37.43423, -37.47606, -37.51764, 
        -37.5592, -37.60115, -37.64353, -37.68629, -37.7292, -37.77183, 
        -37.81392, -37.85496, -37.89452, -37.93251, -37.9691, -38.00468, 
        -38.03997, -38.07523, -38.11072, -38.14546, -38.18142, -38.21774, 
        -38.2544, -38.29126, -38.32808, -38.36401, -38.39836, -38.43045, 
        -38.46019, -38.48804, -38.5146, -38.54057, -38.56621, -38.59167, 
        -38.61597, -38.63992, -38.66331, -38.68567, -38.70629, -38.72695, 
        -38.74557, -38.76288, -38.77864, -38.79278, -38.80603, -38.81865, 
        -38.83076, -38.84292, -38.85549, -38.86882, -38.8829, -38.8972, 
        -38.91122, -38.92437, -38.93651, -38.94813, -38.95967, -38.97195, 
        -38.98459, -39.00021, -39.01828, -39.0388, -39.061, -39.08431, 
        -39.10807, -39.13205, -39.15638, -39.18086, -39.20551, -39.23021, 
        -39.25484, -39.27928, -39.30288, -39.3252, -39.346, -39.36494, 
        -39.38208, -39.39797, -39.41321, -39.42731, -39.44276, -39.45866, 
        -39.47508, -39.49169, -39.50851, -39.52521, -39.54162, -39.55791, 
        -39.57418, -39.59061, -39.60732, -39.62414, -39.64093, -39.65741, 
        -39.67369, -39.68953, -39.70505, -39.72068, -39.73637, -39.75282, 
        -39.77035, -39.78921, -39.80952, -39.83021, -39.8534, -39.87785, 
        -39.90342, -39.92997, -39.95761, -39.98602, -40.01489, -40.04381, 
        -40.07259, -40.10105, -40.12899, -40.15652, -40.18415, -40.21177, 
        -40.23931, -40.26631, -40.2923, -40.31682, -40.33915, -40.3596, 
        -40.37791, -40.39486, -40.41058, -40.42542, -40.439, -40.45158, 
        -40.4615, -40.47047, -40.47721, -40.48173, -40.48441, -40.48544, 
        -40.48574, -40.48552, -40.4852, -40.48525, -40.48633, -40.48903, 
        -40.49355, -40.4996, -40.50647, -40.51373, -40.521, -40.5283, 
        -40.53588, -40.5441, -40.55375, -40.56543, -40.57912, -40.59502, 
        -40.61267, -40.6315, -40.65088, -40.67033, -40.68953, -40.70865, 
        -40.72707, -40.74745, -40.76894, -40.79155, -40.81525, -40.8394, 
        -40.86324, -40.8861, -40.90732, -40.92713, -40.94524, -40.9621, 
        -40.97842, -40.99436, -41.01005, -41.02561, -41.04098, -41.05621, 
        -41.07108, -41.08545, -41.09897, -41.11189, -41.12482, -41.13763, 
        -41.15037, -41.16259, -41.17397, -41.18449, -41.19404, -41.20257, 
        -41.20998, -41.2161, -41.22099, -41.22478, -41.22783, -41.23022, 
        -41.23198, -41.23217, -41.23247, -41.23147, -41.22836, -41.223, 
        -41.21512, -41.20526, -41.19424, -41.18242, -41.16963, -41.15522, 
        -41.13863, -41.11928, -41.09703, -41.07144, -41.04188, -41.00818, 
        -40.96878, -40.92368, -40.87255, -40.81598, -40.75462, -40.6887, 
        -40.61722, -40.53867, -40.45211, -40.35664, -40.25229, -40.13962, 
        -40.02053,
  -34.28282, -34.32418, -34.36607, -34.40877, -34.45203, -34.49531, 
        -34.53805, -34.57896, -34.62016, -34.66097, -34.70161, -34.7421, 
        -34.78221, -34.82166, -34.86023, -34.89796, -34.93503, -34.97182, 
        -35.00872, -35.04607, -35.08416, -35.12317, -35.16219, -35.20319, 
        -35.24519, -35.28822, -35.33213, -35.37661, -35.42103, -35.46456, 
        -35.50657, -35.5467, -35.58504, -35.62223, -35.65925, -35.69706, 
        -35.73612, -35.77531, -35.81623, -35.85754, -35.89913, -35.94102, 
        -35.98307, -36.02486, -36.06594, -36.10619, -36.14589, -36.18558, 
        -36.22579, -36.2668, -36.30854, -36.35052, -36.39198, -36.43126, 
        -36.47028, -36.50854, -36.54669, -36.58514, -36.62384, -36.66256, 
        -36.70122, -36.74002, -36.77938, -36.81972, -36.86115, -36.90337, 
        -36.94578, -36.98806, -37.03001, -37.07208, -37.11356, -37.1565, 
        -37.19989, -37.24343, -37.28677, -37.32969, -37.37214, -37.4144, 
        -37.45685, -37.49976, -37.54314, -37.58682, -37.63054, -37.67383, 
        -37.71627, -37.75748, -37.7972, -37.83444, -37.87125, -37.90719, 
        -37.94292, -37.97889, -38.01524, -38.05188, -38.0888, -38.12587, 
        -38.16312, -38.20039, -38.23726, -38.27313, -38.30692, -38.33837, 
        -38.36744, -38.39471, -38.4208, -38.44546, -38.47092, -38.49617, 
        -38.52116, -38.54573, -38.56985, -38.59336, -38.61599, -38.63731, 
        -38.65691, -38.67477, -38.6907, -38.70523, -38.71845, -38.73098, 
        -38.74318, -38.75558, -38.76866, -38.78265, -38.79742, -38.81145, 
        -38.82613, -38.83993, -38.85271, -38.86472, -38.87674, -38.88951, 
        -38.90371, -38.91982, -38.93832, -38.95908, -38.98141, -39.00484, 
        -39.0289, -39.0534, -39.07825, -39.10342, -39.12875, -39.15416, 
        -39.17935, -39.20408, -39.22707, -39.24952, -39.27008, -39.28878, 
        -39.30547, -39.3208, -39.33553, -39.3505, -39.36596, -39.38221, 
        -39.399, -39.41622, -39.43359, -39.45084, -39.46783, -39.48438, 
        -39.50086, -39.51723, -39.53369, -39.55014, -39.56672, -39.58304, 
        -39.59916, -39.61419, -39.63006, -39.64612, -39.66275, -39.68025, 
        -39.69914, -39.71967, -39.74184, -39.76551, -39.79043, -39.81629, 
        -39.84278, -39.86996, -39.89769, -39.92586, -39.95426, -39.98269, 
        -40.01091, -40.03876, -40.06624, -40.09346, -40.1207, -40.14815, 
        -40.1754, -40.20235, -40.22832, -40.25164, -40.27391, -40.29402, 
        -40.31194, -40.32834, -40.3438, -40.35835, -40.37227, -40.38525, 
        -40.39678, -40.4066, -40.41402, -40.41906, -40.42176, -40.42298, 
        -40.42311, -40.42275, -40.42233, -40.42236, -40.42347, -40.42611, 
        -40.4303, -40.43564, -40.44156, -40.44772, -40.454, -40.46048, 
        -40.46762, -40.47575, -40.4845, -40.49637, -40.51057, -40.52708, 
        -40.54551, -40.5653, -40.58584, -40.60656, -40.62716, -40.64776, 
        -40.6687, -40.69044, -40.71326, -40.73711, -40.76168, -40.78643, 
        -40.81066, -40.83374, -40.85522, -40.87499, -40.89311, -40.91018, 
        -40.9266, -40.94273, -40.9586, -40.97423, -40.98967, -41.00491, 
        -41.01982, -41.03415, -41.04765, -41.06052, -41.07311, -41.08567, 
        -41.09722, -41.10951, -41.12127, -41.13229, -41.14233, -41.1512, 
        -41.15871, -41.16481, -41.16963, -41.17347, -41.17677, -41.17983, 
        -41.18276, -41.18541, -41.18733, -41.1878, -41.18614, -41.18192, 
        -41.17515, -41.16633, -41.15622, -41.14533, -41.13357, -41.12031, 
        -41.1049, -41.08698, -41.06605, -41.04181, -41.01351, -40.98032, 
        -40.94166, -40.89665, -40.84565, -40.78911, -40.72776, -40.6618, 
        -40.59104, -40.51416, -40.42981, -40.33699, -40.23598, -40.1274, 
        -40.01278,
  -34.15664, -34.19833, -34.24053, -34.28241, -34.32571, -34.36897, 
        -34.41166, -34.45353, -34.49467, -34.53532, -34.57557, -34.61578, 
        -34.6553, -34.69452, -34.73272, -34.77069, -34.80803, -34.84425, 
        -34.88147, -34.91925, -34.95812, -34.99821, -35.03962, -35.08214, 
        -35.12536, -35.16972, -35.21442, -35.25949, -35.30391, -35.34706, 
        -35.38859, -35.42846, -35.46568, -35.50301, -35.54021, -35.57808, 
        -35.61699, -35.65692, -35.6977, -35.73907, -35.78093, -35.82312, 
        -35.86552, -35.90757, -35.94901, -35.98969, -36.02985, -36.07008, 
        -36.10963, -36.15107, -36.19298, -36.23521, -36.27695, -36.31742, 
        -36.35683, -36.39568, -36.43454, -36.47385, -36.51336, -36.55299, 
        -36.59252, -36.6321, -36.67209, -36.71283, -36.75347, -36.79576, 
        -36.83811, -36.88026, -36.92227, -36.9649, -37.00804, -37.0518, 
        -37.09601, -37.1404, -37.18426, -37.22779, -37.27068, -37.31344, 
        -37.35662, -37.40033, -37.4445, -37.48789, -37.53212, -37.57578, 
        -37.61843, -37.65972, -37.69946, -37.7377, -37.77473, -37.81108, 
        -37.84747, -37.88429, -37.92181, -37.95947, -37.99701, -38.03476, 
        -38.07224, -38.10965, -38.1464, -38.18089, -38.21433, -38.24527, 
        -38.27397, -38.30095, -38.32714, -38.35308, -38.37869, -38.40409, 
        -38.42946, -38.45465, -38.4794, -38.50383, -38.52724, -38.5493, 
        -38.56937, -38.58755, -38.60388, -38.61843, -38.63089, -38.64351, 
        -38.65593, -38.66883, -38.68253, -38.6973, -38.71268, -38.72831, 
        -38.74348, -38.75759, -38.77077, -38.78335, -38.796, -38.80943, 
        -38.82423, -38.84098, -38.8597, -38.88026, -38.90248, -38.92585, 
        -38.94997, -38.9739, -38.99922, -39.0249, -39.05074, -39.07659, 
        -39.1023, -39.12739, -39.15141, -39.17399, -39.19499, -39.21355, 
        -39.22993, -39.24517, -39.25987, -39.27486, -39.2906, -39.30709, 
        -39.32451, -39.3421, -39.35997, -39.37766, -39.39497, -39.41077, 
        -39.42731, -39.44366, -39.46002, -39.47635, -39.49267, -39.509, 
        -39.52536, -39.54169, -39.55816, -39.57487, -39.59217, -39.61061, 
        -39.63054, -39.65219, -39.67571, -39.7008, -39.72709, -39.75415, 
        -39.78183, -39.80949, -39.83746, -39.86552, -39.89366, -39.92167, 
        -39.94852, -39.97607, -40.00329, -40.03033, -40.05747, -40.08477, 
        -40.11184, -40.13881, -40.16467, -40.18851, -40.21043, -40.23026, 
        -40.24797, -40.26404, -40.27941, -40.29389, -40.30808, -40.32149, 
        -40.33382, -40.34436, -40.35246, -40.3577, -40.36058, -40.36152, 
        -40.36152, -40.36121, -40.36098, -40.36142, -40.36176, -40.36432, 
        -40.36811, -40.37254, -40.37719, -40.38189, -40.38689, -40.39255, 
        -40.39907, -40.40705, -40.41707, -40.4295, -40.44448, -40.46188, 
        -40.4813, -40.50201, -40.52357, -40.54539, -40.5672, -40.5891, 
        -40.61132, -40.63434, -40.65831, -40.68307, -40.70831, -40.73357, 
        -40.75828, -40.78172, -40.80374, -40.82402, -40.84255, -40.85987, 
        -40.87542, -40.89163, -40.90746, -40.92304, -40.93839, -40.95358, 
        -40.96854, -40.983, -40.99667, -41.00965, -41.02208, -41.03437, 
        -41.0466, -41.05871, -41.07044, -41.08148, -41.09158, -41.10035, 
        -41.1078, -41.11378, -41.11866, -41.12283, -41.12669, -41.1309, 
        -41.13531, -41.13954, -41.14301, -41.14489, -41.14442, -41.14121, 
        -41.13533, -41.12733, -41.11795, -41.10799, -41.09724, -41.08522, 
        -41.07114, -41.05451, -41.03484, -41.01163, -40.98415, -40.95061, 
        -40.91202, -40.86674, -40.81611, -40.75951, -40.69818, -40.63256, 
        -40.56222, -40.48645, -40.4039, -40.31344, -40.21516, -40.10999, 
        -39.9997,
  -34.03123, -34.07325, -34.11566, -34.15847, -34.20164, -34.24485, 
        -34.28747, -34.32935, -34.37056, -34.41125, -34.45154, -34.49141, 
        -34.52973, -34.56836, -34.60663, -34.64453, -34.68206, -34.71955, 
        -34.75747, -34.79607, -34.836, -34.87737, -34.9201, -34.96403, 
        -35.00845, -35.05365, -35.09883, -35.14278, -35.18689, -35.22932, 
        -35.2703, -35.30986, -35.3482, -35.38579, -35.42339, -35.46164, 
        -35.5005, -35.5404, -35.58116, -35.62261, -35.66456, -35.70682, 
        -35.74905, -35.78997, -35.83156, -35.87263, -35.91352, -35.95442, 
        -35.99602, -36.03778, -36.07994, -36.12246, -36.16423, -36.20497, 
        -36.24492, -36.28428, -36.32387, -36.36392, -36.40427, -36.44369, 
        -36.48392, -36.52414, -36.56467, -36.60578, -36.64753, -36.6897, 
        -36.73191, -36.77387, -36.81649, -36.86002, -36.9042, -36.94913, 
        -36.99451, -37.03952, -37.0843, -37.12697, -37.17031, -37.21366, 
        -37.25742, -37.30174, -37.34646, -37.3913, -37.43585, -37.47969, 
        -37.5225, -37.56382, -37.6036, -37.64192, -37.67915, -37.71597, 
        -37.75314, -37.79085, -37.82917, -37.86672, -37.90528, -37.94297, 
        -37.98058, -38.01805, -38.0543, -38.08937, -38.12226, -38.15309, 
        -38.18182, -38.20905, -38.23565, -38.2617, -38.28773, -38.31396, 
        -38.33999, -38.36583, -38.39138, -38.41627, -38.43914, -38.46152, 
        -38.48203, -38.50045, -38.51702, -38.53176, -38.54531, -38.55824, 
        -38.57117, -38.58467, -38.59904, -38.61435, -38.63024, -38.64617, 
        -38.66154, -38.67596, -38.68954, -38.70276, -38.71618, -38.73032, 
        -38.74479, -38.76183, -38.78058, -38.80099, -38.82286, -38.84602, 
        -38.87037, -38.8956, -38.92137, -38.9473, -38.97334, -38.99939, 
        -39.02531, -39.0507, -39.075, -39.09818, -39.1193, -39.13817, 
        -39.15499, -39.17048, -39.18536, -39.20055, -39.2155, -39.23236, 
        -39.25006, -39.26802, -39.28592, -39.30387, -39.32129, -39.33841, 
        -39.35529, -39.37177, -39.38809, -39.40425, -39.42057, -39.43705, 
        -39.45367, -39.47054, -39.48764, -39.50506, -39.52317, -39.54233, 
        -39.56303, -39.5856, -39.60992, -39.63589, -39.66217, -39.69012, 
        -39.71864, -39.74712, -39.77549, -39.80358, -39.83167, -39.85961, 
        -39.88741, -39.915, -39.94226, -39.96939, -39.99644, -40.02366, 
        -40.05084, -40.07744, -40.10267, -40.12627, -40.14785, -40.1673, 
        -40.185, -40.20125, -40.21663, -40.23167, -40.24617, -40.26009, 
        -40.2718, -40.28279, -40.291, -40.29644, -40.2993, -40.30028, 
        -40.30017, -40.29999, -40.30011, -40.30087, -40.30252, -40.30509, 
        -40.30806, -40.31137, -40.31475, -40.31807, -40.32178, -40.32627, 
        -40.33209, -40.33983, -40.35025, -40.36358, -40.37975, -40.39841, 
        -40.41902, -40.44098, -40.46349, -40.48629, -40.50904, -40.53197, 
        -40.55519, -40.57817, -40.60304, -40.62847, -40.65417, -40.67998, 
        -40.70533, -40.72964, -40.75242, -40.7734, -40.79253, -40.81027, 
        -40.82708, -40.84312, -40.85884, -40.87421, -40.88934, -40.90441, 
        -40.91927, -40.93382, -40.94762, -40.96067, -40.97312, -40.98521, 
        -40.99712, -41.0089, -41.02032, -41.0311, -41.04079, -41.04926, 
        -41.05643, -41.06242, -41.06754, -41.07233, -41.07701, -41.08237, 
        -41.08834, -41.09419, -41.09817, -41.10126, -41.10182, -41.09947, 
        -41.0944, -41.08718, -41.07862, -41.06939, -41.05953, -41.04862, 
        -41.03582, -41.02057, -41.00196, -40.97945, -40.95247, -40.92017, 
        -40.88174, -40.83682, -40.78555, -40.72915, -40.66826, -40.60299, 
        -40.53318, -40.458, -40.37675, -40.28864, -40.19311, -40.09114, 
        -39.98407,
  -33.90888, -33.95114, -33.99376, -34.03665, -34.0796, -34.12243, 
        -34.16495, -34.20695, -34.2472, -34.28811, -34.32851, -34.36841, 
        -34.40763, -34.44619, -34.48428, -34.52206, -34.5598, -34.59771, 
        -34.6362, -34.67605, -34.71709, -34.7598, -34.80278, -34.84772, 
        -34.89305, -34.93864, -34.98391, -35.02845, -35.0718, -35.11372, 
        -35.15424, -35.19354, -35.23212, -35.27045, -35.30855, -35.34715, 
        -35.38649, -35.42541, -35.46606, -35.50749, -35.54933, -35.59126, 
        -35.63306, -35.67457, -35.71608, -35.75752, -35.79921, -35.84121, 
        -35.88336, -35.92588, -35.96867, -36.01104, -36.05305, -36.09315, 
        -36.13359, -36.1737, -36.21407, -36.25489, -36.29586, -36.33686, 
        -36.37767, -36.41842, -36.45937, -36.50066, -36.54241, -36.58443, 
        -36.62645, -36.66888, -36.71219, -36.75644, -36.80082, -36.84704, 
        -36.89353, -36.93957, -36.98479, -37.02914, -37.07294, -37.11676, 
        -37.16098, -37.20575, -37.2508, -37.29587, -37.34061, -37.3846, 
        -37.4275, -37.46899, -37.509, -37.54654, -37.5841, -37.62147, 
        -37.65924, -37.69768, -37.73686, -37.77614, -37.81486, -37.85294, 
        -37.89028, -37.92707, -37.963, -37.99746, -38.03024, -38.06116, 
        -38.09041, -38.11836, -38.14561, -38.17253, -38.19835, -38.22518, 
        -38.25193, -38.27832, -38.30442, -38.32973, -38.35375, -38.37628, 
        -38.39693, -38.41547, -38.43213, -38.44711, -38.46106, -38.47443, 
        -38.48809, -38.5023, -38.5173, -38.53302, -38.54903, -38.56387, 
        -38.57911, -38.59354, -38.60752, -38.62139, -38.63582, -38.65102, 
        -38.66721, -38.68458, -38.70324, -38.72324, -38.74468, -38.7677, 
        -38.79207, -38.81749, -38.8436, -38.86979, -38.89591, -38.92198, 
        -38.94788, -38.97321, -38.99784, -39.02029, -39.04207, -39.06166, 
        -39.07939, -39.09557, -39.11092, -39.12654, -39.14267, -39.15964, 
        -39.1771, -39.19517, -39.21319, -39.23124, -39.24899, -39.26651, 
        -39.28363, -39.30043, -39.3168, -39.33307, -39.34954, -39.36617, 
        -39.38314, -39.40076, -39.41752, -39.43573, -39.45474, -39.47481, 
        -39.49631, -39.51949, -39.54436, -39.5707, -39.59844, -39.62698, 
        -39.65592, -39.68533, -39.71408, -39.74268, -39.77072, -39.7988, 
        -39.82672, -39.85464, -39.88213, -39.90967, -39.93711, -39.96445, 
        -39.9913, -40.01717, -40.04174, -40.06379, -40.08503, -40.10443, 
        -40.12233, -40.13888, -40.15475, -40.17028, -40.1855, -40.19986, 
        -40.21297, -40.22377, -40.23176, -40.23707, -40.23988, -40.24088, 
        -40.24094, -40.24089, -40.24118, -40.24232, -40.2441, -40.24607, 
        -40.24829, -40.25033, -40.2524, -40.25425, -40.25664, -40.26002, 
        -40.26503, -40.27278, -40.28272, -40.29707, -40.3148, -40.33519, 
        -40.35746, -40.3808, -40.40462, -40.42844, -40.45212, -40.47574, 
        -40.49978, -40.52468, -40.54997, -40.57581, -40.60218, -40.6288, 
        -40.65486, -40.67993, -40.70346, -40.72515, -40.74487, -40.76309, 
        -40.78, -40.79614, -40.81181, -40.82689, -40.84171, -40.85649, 
        -40.87119, -40.88553, -40.89929, -40.91229, -40.92474, -40.93669, 
        -40.94841, -40.9589, -40.96996, -40.98027, -40.98958, -40.9976, 
        -41.0045, -41.01059, -41.01613, -41.02152, -41.0273, -41.03395, 
        -41.04111, -41.04818, -41.0543, -41.0584, -41.05981, -41.05824, 
        -41.05397, -41.04761, -41.0398, -41.03128, -41.02215, -41.01208, 
        -41.00028, -40.9859, -40.96814, -40.94627, -40.91949, -40.88709, 
        -40.84921, -40.80454, -40.75414, -40.6979, -40.6374, -40.57264, 
        -40.50318, -40.42878, -40.34851, -40.26193, -40.16876, -40.06926, 
        -39.96487,
  -33.78872, -33.83133, -33.87417, -33.91606, -33.95895, -34.00154, 
        -34.0437, -34.08556, -34.12708, -34.16822, -34.20888, -34.24883, 
        -34.28806, -34.32651, -34.36445, -34.40222, -34.44016, -34.47755, 
        -34.51701, -34.55772, -34.60003, -34.64392, -34.689, -34.73477, 
        -34.78063, -34.82625, -34.87128, -34.9152, -34.95794, -34.99936, 
        -35.03959, -35.07909, -35.11695, -35.15582, -35.19479, -35.234, 
        -35.27371, -35.31387, -35.35454, -35.39579, -35.43729, -35.47873, 
        -35.52003, -35.5612, -35.60248, -35.64435, -35.68658, -35.72932, 
        -35.77129, -35.8144, -35.85749, -35.90024, -35.94242, -35.98394, 
        -36.02494, -36.06586, -36.10702, -36.14851, -36.19011, -36.23166, 
        -36.27304, -36.31427, -36.35557, -36.39713, -36.43785, -36.47983, 
        -36.52206, -36.56472, -36.60844, -36.65343, -36.69987, -36.74712, 
        -36.79454, -36.84148, -36.88749, -36.93266, -36.97717, -37.0216, 
        -37.0664, -37.11136, -37.15658, -37.20072, -37.24554, -37.2895, 
        -37.33259, -37.37431, -37.41468, -37.45371, -37.49191, -37.52981, 
        -37.56797, -37.60685, -37.64634, -37.68594, -37.72494, -37.76298, 
        -37.80022, -37.83663, -37.87217, -37.90636, -37.93807, -37.96933, 
        -37.99932, -38.02824, -38.05648, -38.0844, -38.11203, -38.13953, 
        -38.1668, -38.19384, -38.22015, -38.24567, -38.26968, -38.29229, 
        -38.31279, -38.33148, -38.34837, -38.36369, -38.37818, -38.39145, 
        -38.40581, -38.42058, -38.43599, -38.45184, -38.46771, -38.4832, 
        -38.4982, -38.51258, -38.52679, -38.54139, -38.55672, -38.57282, 
        -38.58982, -38.6077, -38.62652, -38.64639, -38.6676, -38.69033, 
        -38.71456, -38.7391, -38.76526, -38.7916, -38.81778, -38.84375, 
        -38.86969, -38.8952, -38.92002, -38.9439, -38.96627, -38.98677, 
        -39.00536, -39.02241, -39.03833, -39.0541, -39.07035, -39.0872, 
        -39.10449, -39.12222, -39.14027, -39.15835, -39.17656, -39.19453, 
        -39.21122, -39.22852, -39.24527, -39.2618, -39.27854, -39.29564, 
        -39.31311, -39.3311, -39.34985, -39.36891, -39.38884, -39.40993, 
        -39.43237, -39.45626, -39.48156, -39.50816, -39.5358, -39.56445, 
        -39.59363, -39.62333, -39.65279, -39.68152, -39.71016, -39.73846, 
        -39.76585, -39.79425, -39.8224, -39.85025, -39.878, -39.90538, 
        -39.93174, -39.95687, -39.98071, -40.00319, -40.0243, -40.04389, 
        -40.06216, -40.0794, -40.09606, -40.11224, -40.12799, -40.14285, 
        -40.15572, -40.16627, -40.17405, -40.17911, -40.18187, -40.18299, 
        -40.18311, -40.18319, -40.18356, -40.18457, -40.18477, -40.18612, 
        -40.18707, -40.18792, -40.18874, -40.18929, -40.19037, -40.19271, 
        -40.19724, -40.20467, -40.21603, -40.23173, -40.25112, -40.27357, 
        -40.29788, -40.32315, -40.34867, -40.37388, -40.3986, -40.42325, 
        -40.44819, -40.47338, -40.49929, -40.52603, -40.55281, -40.57973, 
        -40.60637, -40.63198, -40.65606, -40.67818, -40.69831, -40.71684, 
        -40.73402, -40.74933, -40.76496, -40.77997, -40.79459, -40.80906, 
        -40.82336, -40.83734, -40.85079, -40.86361, -40.87577, -40.88764, 
        -40.8993, -40.91064, -40.92151, -40.93158, -40.94043, -40.94819, 
        -40.95503, -40.96127, -40.96728, -40.97332, -40.97996, -40.9874, 
        -40.99549, -41.00342, -41.01025, -41.01506, -41.01723, -41.01641, 
        -41.01302, -41.00741, -41.00033, -40.99228, -40.98367, -40.97413, 
        -40.96299, -40.9493, -40.93225, -40.91083, -40.88449, -40.85258, 
        -40.8136, -40.77001, -40.72041, -40.66533, -40.60556, -40.54107, 
        -40.47206, -40.39794, -40.31837, -40.23314, -40.14187, -40.04467, 
        -39.94227,
  -33.66955, -33.7127, -33.75571, -33.79867, -33.84129, -33.88366, 
        -33.92566, -33.96738, -34.0089, -34.05013, -34.09092, -34.13114, 
        -34.17031, -34.20789, -34.24576, -34.28366, -34.32198, -34.36109, 
        -34.40137, -34.44314, -34.48657, -34.53153, -34.57751, -34.62377, 
        -34.6699, -34.71538, -34.76004, -34.80239, -34.8445, -34.88557, 
        -34.92589, -34.96535, -35.0048, -35.04453, -35.08443, -35.1241, 
        -35.16448, -35.20472, -35.24546, -35.28648, -35.32757, -35.36868, 
        -35.40945, -35.4494, -35.49068, -35.5326, -35.57526, -35.61854, 
        -35.66208, -35.7057, -35.7492, -35.7923, -35.83481, -35.8768, 
        -35.91842, -35.95999, -36.00175, -36.0438, -36.086, -36.12703, 
        -36.1689, -36.21064, -36.25239, -36.29426, -36.33619, -36.37827, 
        -36.42062, -36.4636, -36.50774, -36.55336, -36.60044, -36.64847, 
        -36.6967, -36.7445, -36.79145, -36.8375, -36.88211, -36.92739, 
        -36.97269, -37.01797, -37.06336, -37.10843, -37.15294, -37.19697, 
        -37.23985, -37.28201, -37.32285, -37.36252, -37.40135, -37.43976, 
        -37.47835, -37.51749, -37.55715, -37.59684, -37.63494, -37.67308, 
        -37.71024, -37.7465, -37.78176, -37.81589, -37.84877, -37.88052, 
        -37.91135, -37.9413, -37.97072, -37.99972, -38.02826, -38.05641, 
        -38.08387, -38.11093, -38.13765, -38.16312, -38.18604, -38.20835, 
        -38.22894, -38.24768, -38.26493, -38.28082, -38.29591, -38.31086, 
        -38.32587, -38.34118, -38.35675, -38.37262, -38.38821, -38.40327, 
        -38.41791, -38.43226, -38.44681, -38.46205, -38.47825, -38.49533, 
        -38.51327, -38.53087, -38.55013, -38.5701, -38.59127, -38.61378, 
        -38.63781, -38.66309, -38.68907, -38.71534, -38.7414, -38.76721, 
        -38.79301, -38.81855, -38.84359, -38.86782, -38.89083, -38.91212, 
        -38.93163, -38.94934, -38.96593, -38.98204, -38.99719, -39.01376, 
        -39.03083, -39.04832, -39.06641, -39.08473, -39.10332, -39.12188, 
        -39.14019, -39.15811, -39.17546, -39.19239, -39.20958, -39.22718, 
        -39.24532, -39.26405, -39.28334, -39.30355, -39.32455, -39.34672, 
        -39.37013, -39.39472, -39.42041, -39.44722, -39.47386, -39.50229, 
        -39.53154, -39.56122, -39.59095, -39.62017, -39.64927, -39.67828, 
        -39.70729, -39.73633, -39.76527, -39.79356, -39.82154, -39.84853, 
        -39.8742, -39.89861, -39.92172, -39.94381, -39.96474, -39.98458, 
        -40.00348, -40.02161, -40.03903, -40.05594, -40.07221, -40.08701, 
        -40.09975, -40.10884, -40.11623, -40.12105, -40.12374, -40.12504, 
        -40.12537, -40.12552, -40.12579, -40.12614, -40.12663, -40.12694, 
        -40.12669, -40.12622, -40.12557, -40.12493, -40.12489, -40.12629, 
        -40.13026, -40.13763, -40.14964, -40.16637, -40.18748, -40.2124, 
        -40.23907, -40.26669, -40.29444, -40.32141, -40.34789, -40.37383, 
        -40.39963, -40.42451, -40.45089, -40.47785, -40.50499, -40.5322, 
        -40.55899, -40.58481, -40.60904, -40.63131, -40.65161, -40.67025, 
        -40.68765, -40.70416, -40.72, -40.73514, -40.74977, -40.76395, 
        -40.77789, -40.79126, -40.80419, -40.8166, -40.82865, -40.84029, 
        -40.85195, -40.86337, -40.87426, -40.88433, -40.89302, -40.90089, 
        -40.90786, -40.91439, -40.92073, -40.92735, -40.9346, -40.94243, 
        -40.95086, -40.95914, -40.96631, -40.97054, -40.97313, -40.97301, 
        -40.97027, -40.96548, -40.95903, -40.95152, -40.94318, -40.93396, 
        -40.92307, -40.90984, -40.8932, -40.87234, -40.84676, -40.81554, 
        -40.77849, -40.73567, -40.6872, -40.63315, -40.57422, -40.51013, 
        -40.44122, -40.36777, -40.289, -40.20497, -40.11494, -40.01953, 
        -39.91883,
  -33.55312, -33.5968, -33.6401, -33.683, -33.72548, -33.76754, 
        -33.80931, -33.85101, -33.89145, -33.93285, -33.97366, -34.01397, 
        -34.0533, -34.09193, -34.13011, -34.16832, -34.20705, -34.24688, 
        -34.2881, -34.33087, -34.3753, -34.42096, -34.46753, -34.51334, 
        -34.55936, -34.6047, -34.64877, -34.69167, -34.73348, -34.77454, 
        -34.81488, -34.85493, -34.89497, -34.93534, -34.97571, -35.01629, 
        -35.05702, -35.09766, -35.13743, -35.17831, -35.21912, -35.25987, 
        -35.30054, -35.34136, -35.38271, -35.42477, -35.46767, -35.51121, 
        -35.55514, -35.59917, -35.64306, -35.68653, -35.72945, -35.77184, 
        -35.81297, -35.85502, -35.89727, -35.93972, -35.98228, -36.02473, 
        -36.06709, -36.10935, -36.15165, -36.19407, -36.23642, -36.27888, 
        -36.32146, -36.3648, -36.40931, -36.45532, -36.50164, -36.54996, 
        -36.59866, -36.64717, -36.69522, -36.7426, -36.78944, -36.83575, 
        -36.88169, -36.92729, -36.97269, -37.01765, -37.06217, -37.10584, 
        -37.14896, -37.19117, -37.23254, -37.27288, -37.31151, -37.35059, 
        -37.38954, -37.42873, -37.46828, -37.50795, -37.54723, -37.58576, 
        -37.62313, -37.6595, -37.69477, -37.72897, -37.76219, -37.79449, 
        -37.82606, -37.85699, -37.88739, -37.91716, -37.94492, -37.97352, 
        -38.0012, -38.02872, -38.05515, -38.08061, -38.10434, -38.12648, 
        -38.147, -38.16599, -38.1835, -38.19984, -38.21556, -38.23101, 
        -38.24652, -38.26221, -38.27803, -38.29381, -38.30913, -38.32394, 
        -38.3373, -38.35176, -38.36669, -38.38261, -38.39961, -38.41773, 
        -38.43672, -38.4563, -38.47632, -38.49675, -38.51798, -38.54027, 
        -38.56396, -38.58884, -38.61448, -38.64031, -38.66614, -38.69175, 
        -38.71758, -38.743, -38.76805, -38.79145, -38.81511, -38.83714, 
        -38.85725, -38.87574, -38.8928, -38.90907, -38.92519, -38.94158, 
        -38.95836, -38.97583, -38.99396, -39.0127, -39.03178, -39.05095, 
        -39.06993, -39.08841, -39.10631, -39.12385, -39.14151, -39.1596, 
        -39.17834, -39.19777, -39.21685, -39.2381, -39.26036, -39.28377, 
        -39.30834, -39.33391, -39.36015, -39.38708, -39.41455, -39.44284, 
        -39.4719, -39.50151, -39.53122, -39.56087, -39.59044, -39.62014, 
        -39.64991, -39.67959, -39.70912, -39.73775, -39.76569, -39.79227, 
        -39.81742, -39.8411, -39.86357, -39.8852, -39.9051, -39.9254, 
        -39.94489, -39.9637, -39.98195, -39.99962, -40.01608, -40.03074, 
        -40.0431, -40.0526, -40.05947, -40.06411, -40.06694, -40.06839, 
        -40.06891, -40.06905, -40.06894, -40.06872, -40.06821, -40.06712, 
        -40.0657, -40.06402, -40.06218, -40.06024, -40.05911, -40.05971, 
        -40.06326, -40.07091, -40.08348, -40.10064, -40.12382, -40.15091, 
        -40.18024, -40.21055, -40.24065, -40.26998, -40.29815, -40.32556, 
        -40.35267, -40.37938, -40.40631, -40.4334, -40.46076, -40.48801, 
        -40.51471, -40.54048, -40.56445, -40.58647, -40.60659, -40.62519, 
        -40.64264, -40.65942, -40.6756, -40.69114, -40.70598, -40.72012, 
        -40.73363, -40.7465, -40.75867, -40.7705, -40.78195, -40.79359, 
        -40.80534, -40.8171, -40.82737, -40.83768, -40.84668, -40.85496, 
        -40.86223, -40.86912, -40.8759, -40.88292, -40.89038, -40.89836, 
        -40.90664, -40.91472, -40.92157, -40.92681, -40.92977, -40.93018, 
        -40.92822, -40.92404, -40.918, -40.91084, -40.90268, -40.89357, 
        -40.88274, -40.86967, -40.85349, -40.83337, -40.80849, -40.77837, 
        -40.74245, -40.70078, -40.65329, -40.60033, -40.54206, -40.47874, 
        -40.41025, -40.33734, -40.25942, -40.17647, -40.08802, -39.99384, 
        -39.89442,
  -33.43797, -33.48238, -33.52602, -33.56799, -33.61033, -33.65211, 
        -33.69363, -33.73511, -33.77635, -33.81769, -33.85866, -33.8987, 
        -33.9383, -33.9773, -34.01575, -34.05443, -34.09388, -34.13466, 
        -34.17594, -34.21975, -34.26513, -34.31168, -34.35866, -34.40543, 
        -34.45137, -34.4962, -34.5398, -34.58232, -34.62398, -34.665, 
        -34.70564, -34.74601, -34.78655, -34.8264, -34.86749, -34.90866, 
        -34.94974, -34.9908, -35.03183, -35.0728, -35.11378, -35.15473, 
        -35.19555, -35.23649, -35.278, -35.32018, -35.36317, -35.40695, 
        -35.45011, -35.49442, -35.53854, -35.58232, -35.62558, -35.66826, 
        -35.71062, -35.75292, -35.79543, -35.83807, -35.88078, -35.92359, 
        -35.96635, -36.00915, -36.05206, -36.09505, -36.13817, -36.18002, 
        -36.22331, -36.26718, -36.31186, -36.35794, -36.4054, -36.45383, 
        -36.50294, -36.55218, -36.60132, -36.6502, -36.69841, -36.74583, 
        -36.79253, -36.83855, -36.88401, -36.92892, -36.97231, -37.01607, 
        -37.05912, -37.1016, -37.14328, -37.18417, -37.22451, -37.26419, 
        -37.30361, -37.34306, -37.38276, -37.42255, -37.46193, -37.50069, 
        -37.53834, -37.57495, -37.61051, -37.64505, -37.6777, -37.71055, 
        -37.74284, -37.77458, -37.8056, -37.83565, -37.86488, -37.89334, 
        -37.92137, -37.94836, -37.97499, -38.00007, -38.02373, -38.0457, 
        -38.06617, -38.08527, -38.10303, -38.11983, -38.13604, -38.15095, 
        -38.16693, -38.18298, -38.19884, -38.21441, -38.22956, -38.24417, 
        -38.25853, -38.27317, -38.2886, -38.30513, -38.32298, -38.34219, 
        -38.36233, -38.38309, -38.40411, -38.42528, -38.44669, -38.4689, 
        -38.49215, -38.51649, -38.54052, -38.56586, -38.59132, -38.61665, 
        -38.64167, -38.66676, -38.69182, -38.71662, -38.74073, -38.7633, 
        -38.78424, -38.80342, -38.82096, -38.83755, -38.85379, -38.8699, 
        -38.88695, -38.9044, -38.92273, -38.94171, -38.96111, -38.9807, 
        -38.99919, -39.01832, -39.03688, -39.05507, -39.07333, -39.09195, 
        -39.11119, -39.1313, -39.15238, -39.17458, -39.19813, -39.22279, 
        -39.24844, -39.27488, -39.3018, -39.32889, -39.35635, -39.38458, 
        -39.41354, -39.44299, -39.47269, -39.50255, -39.53258, -39.56287, 
        -39.59351, -39.62298, -39.6529, -39.68169, -39.70937, -39.73546, 
        -39.75998, -39.78297, -39.80515, -39.82648, -39.84734, -39.86779, 
        -39.88775, -39.90721, -39.92608, -39.94399, -39.96064, -39.975, 
        -39.98679, -39.99578, -40.00232, -40.00671, -40.00952, -40.01128, 
        -40.01202, -40.01225, -40.01187, -40.01109, -40.00965, -40.00636, 
        -40.00365, -40.00076, -39.99759, -39.99447, -39.99234, -39.9924, 
        -39.99589, -40.00392, -40.01743, -40.03706, -40.06241, -40.09192, 
        -40.12418, -40.1573, -40.18994, -40.22169, -40.25194, -40.28096, 
        -40.30905, -40.33665, -40.36395, -40.39119, -40.4185, -40.44562, 
        -40.47208, -40.49729, -40.52085, -40.54238, -40.56218, -40.58076, 
        -40.59837, -40.61435, -40.63105, -40.64701, -40.66215, -40.67636, 
        -40.68976, -40.70218, -40.71372, -40.72477, -40.73584, -40.74712, 
        -40.75879, -40.77071, -40.78237, -40.79313, -40.80292, -40.81168, 
        -40.8196, -40.82705, -40.83426, -40.84157, -40.84907, -40.85679, 
        -40.8646, -40.87204, -40.87851, -40.88344, -40.88646, -40.88717, 
        -40.88573, -40.88215, -40.87663, -40.8696, -40.86154, -40.85229, 
        -40.84153, -40.82843, -40.81253, -40.7929, -40.76904, -40.73981, 
        -40.70495, -40.66355, -40.61703, -40.56525, -40.50786, -40.445, 
        -40.37753, -40.30527, -40.22834, -40.1465, -40.05946, -39.96665, 
        -39.86835,
  -33.32293, -33.36816, -33.41234, -33.45556, -33.49782, -33.53948, 
        -33.58085, -33.62188, -33.66295, -33.70397, -33.74474, -33.78504, 
        -33.8249, -33.86303, -33.90199, -33.94128, -33.98156, -34.02328, 
        -34.0666, -34.11161, -34.15786, -34.20486, -34.25195, -34.29847, 
        -34.34401, -34.38852, -34.4318, -34.47414, -34.51481, -34.55602, 
        -34.59692, -34.63768, -34.67858, -34.71974, -34.76136, -34.80285, 
        -34.84402, -34.88559, -34.92723, -34.96874, -35.01031, -35.05182, 
        -35.0931, -35.1336, -35.17529, -35.21766, -35.26068, -35.30441, 
        -35.34858, -35.39299, -35.43742, -35.48135, -35.52469, -35.56752, 
        -35.61002, -35.65245, -35.69497, -35.73764, -35.78046, -35.82244, 
        -35.86552, -35.90891, -35.95246, -35.99611, -36.03979, -36.08347, 
        -36.12745, -36.17182, -36.21735, -36.2633, -36.31067, -36.35917, 
        -36.4086, -36.45873, -36.50911, -36.55926, -36.6077, -36.65619, 
        -36.70369, -36.75019, -36.79591, -36.84097, -36.88544, -36.92931, 
        -36.97252, -37.01511, -37.05707, -37.09843, -37.13924, -37.17943, 
        -37.21928, -37.25888, -37.29892, -37.33898, -37.37779, -37.41697, 
        -37.45509, -37.49207, -37.52805, -37.56296, -37.59711, -37.63059, 
        -37.66345, -37.69569, -37.72702, -37.75727, -37.78627, -37.81461, 
        -37.84218, -37.86911, -37.89527, -37.92019, -37.94359, -37.96448, 
        -37.98497, -38.00415, -38.02219, -38.03919, -38.05569, -38.07215, 
        -38.08853, -38.1048, -38.1209, -38.13648, -38.15151, -38.1661, 
        -38.18068, -38.19577, -38.21165, -38.22866, -38.24741, -38.26766, 
        -38.28901, -38.31002, -38.33219, -38.35414, -38.37601, -38.39819, 
        -38.42105, -38.44484, -38.46924, -38.49402, -38.51886, -38.54361, 
        -38.56839, -38.59291, -38.61789, -38.64317, -38.66734, -38.6904, 
        -38.71194, -38.73167, -38.74978, -38.76683, -38.78337, -38.7988, 
        -38.81588, -38.8335, -38.85209, -38.8713, -38.891, -38.91094, 
        -38.93084, -38.95047, -38.96968, -38.98857, -39.00739, -39.02643, 
        -39.04609, -39.06671, -39.08854, -39.11181, -39.13644, -39.16224, 
        -39.18898, -39.21628, -39.2438, -39.27136, -39.29898, -39.32628, 
        -39.35518, -39.38457, -39.41417, -39.44405, -39.47429, -39.50516, 
        -39.53636, -39.56727, -39.59736, -39.62606, -39.65327, -39.67883, 
        -39.70281, -39.72564, -39.74751, -39.76873, -39.7897, -39.81026, 
        -39.83057, -39.85051, -39.86973, -39.88771, -39.90405, -39.91808, 
        -39.92942, -39.93692, -39.94305, -39.9473, -39.95025, -39.95208, 
        -39.95306, -39.95345, -39.95308, -39.95188, -39.94952, -39.94633, 
        -39.94259, -39.93842, -39.9341, -39.93011, -39.92743, -39.9272, 
        -39.93082, -39.93933, -39.95427, -39.97565, -40.0031, -40.03509, 
        -40.06993, -40.10568, -40.14092, -40.17479, -40.207, -40.23764, 
        -40.26709, -40.29543, -40.32212, -40.34952, -40.37672, -40.40354, 
        -40.42948, -40.4541, -40.47692, -40.49793, -40.51742, -40.53579, 
        -40.55341, -40.57086, -40.58786, -40.6042, -40.61977, -40.63452, 
        -40.64794, -40.66011, -40.67119, -40.68161, -40.69198, -40.70282, 
        -40.71423, -40.72612, -40.73796, -40.74928, -40.75973, -40.76927, 
        -40.77809, -40.78635, -40.79422, -40.80178, -40.80918, -40.81649, 
        -40.82344, -40.82996, -40.83564, -40.8401, -40.84203, -40.84307, 
        -40.84203, -40.83894, -40.83377, -40.8271, -40.81895, -40.80946, 
        -40.79823, -40.78492, -40.76886, -40.74979, -40.72656, -40.69854, 
        -40.66497, -40.62563, -40.58046, -40.52959, -40.47311, -40.41129, 
        -40.34449, -40.27335, -40.19771, -40.11749, -40.03187, -39.94072, 
        -39.8437,
  -33.21018, -33.25612, -33.30104, -33.34457, -33.38703, -33.42864, 
        -33.4697, -33.51054, -33.55037, -33.59118, -33.63181, -33.67211, 
        -33.71198, -33.75146, -33.79091, -33.83092, -33.87209, -33.91483, 
        -33.95927, -34.0052, -34.0521, -34.09938, -34.14638, -34.19164, 
        -34.23685, -34.28096, -34.32408, -34.36645, -34.40831, -34.44982, 
        -34.49106, -34.53217, -34.57333, -34.61464, -34.65616, -34.69777, 
        -34.73933, -34.78147, -34.82268, -34.86505, -34.90747, -34.94982, 
        -34.99201, -35.03411, -35.07628, -35.11877, -35.16174, -35.20533, 
        -35.24942, -35.29386, -35.33816, -35.38195, -35.42533, -35.46816, 
        -35.50972, -35.55222, -35.59478, -35.63747, -35.68034, -35.72345, 
        -35.76687, -35.81065, -35.85472, -35.89898, -35.94329, -35.98768, 
        -36.0323, -36.0774, -36.12323, -36.16986, -36.21746, -36.26517, 
        -36.31499, -36.36584, -36.41723, -36.46851, -36.51905, -36.56848, 
        -36.6167, -36.66379, -36.70995, -36.7554, -36.80025, -36.84445, 
        -36.88794, -36.93077, -36.97297, -37.01465, -37.05481, -37.09541, 
        -37.13553, -37.17552, -37.21575, -37.25619, -37.29651, -37.3362, 
        -37.37484, -37.41232, -37.44869, -37.48413, -37.51885, -37.55295, 
        -37.58641, -37.61903, -37.65046, -37.6805, -37.70906, -37.73569, 
        -37.76272, -37.78923, -37.81501, -37.83977, -37.86295, -37.8848, 
        -37.90541, -37.9246, -37.9427, -37.9599, -37.9767, -37.99339, 
        -38.01009, -38.02681, -38.04313, -38.05885, -38.07395, -38.08868, 
        -38.10248, -38.11788, -38.1343, -38.15218, -38.1718, -38.19293, 
        -38.21541, -38.23864, -38.26194, -38.28484, -38.3073, -38.32963, 
        -38.35227, -38.37553, -38.39931, -38.42337, -38.44746, -38.47151, 
        -38.49567, -38.52013, -38.54514, -38.5691, -38.59377, -38.61752, 
        -38.63955, -38.6599, -38.67867, -38.69629, -38.71326, -38.73029, 
        -38.74757, -38.76551, -38.78426, -38.80364, -38.82363, -38.84386, 
        -38.86409, -38.88428, -38.90414, -38.92368, -38.94302, -38.9624, 
        -38.9823, -39.00322, -39.02558, -39.04858, -39.07412, -39.10088, 
        -39.12849, -39.15655, -39.1847, -39.21285, -39.241, -39.26984, 
        -39.29888, -39.32811, -39.35752, -39.38731, -39.41771, -39.44875, 
        -39.48013, -39.51118, -39.54105, -39.56926, -39.59586, -39.6209, 
        -39.64458, -39.66719, -39.68901, -39.7104, -39.73041, -39.75136, 
        -39.77188, -39.79205, -39.8114, -39.82922, -39.84516, -39.85867, 
        -39.86947, -39.87766, -39.88362, -39.88795, -39.89092, -39.89294, 
        -39.89427, -39.89477, -39.89441, -39.89291, -39.89022, -39.88621, 
        -39.88148, -39.87621, -39.87095, -39.86638, -39.86336, -39.86319, 
        -39.86739, -39.87724, -39.89362, -39.9159, -39.94545, -39.97985, 
        -40.01704, -40.055, -40.09244, -40.12833, -40.16229, -40.19437, 
        -40.22475, -40.25378, -40.28187, -40.3094, -40.33656, -40.36313, 
        -40.38864, -40.41262, -40.43493, -40.45544, -40.47459, -40.49287, 
        -40.51065, -40.52827, -40.54562, -40.5625, -40.57861, -40.59361, 
        -40.60721, -40.61931, -40.63005, -40.63993, -40.64968, -40.65988, 
        -40.6708, -40.68233, -40.69308, -40.70465, -40.71564, -40.72604, 
        -40.73585, -40.74506, -40.75364, -40.76156, -40.76887, -40.77561, 
        -40.78178, -40.78721, -40.79198, -40.79586, -40.79858, -40.79979, 
        -40.79923, -40.79646, -40.79169, -40.78498, -40.77672, -40.76679, 
        -40.75483, -40.74093, -40.72466, -40.70569, -40.68309, -40.65607, 
        -40.62382, -40.58588, -40.54206, -40.49234, -40.43686, -40.37606, 
        -40.31032, -40.24027, -40.16614, -40.08761, -40.00416, -39.91504, 
        -39.82011,
  -33.09865, -33.14545, -33.19104, -33.23515, -33.27693, -33.31854, 
        -33.35942, -33.39997, -33.44064, -33.48134, -33.52191, -33.56219, 
        -33.60213, -33.64189, -33.68178, -33.72252, -33.7646, -33.8083, 
        -33.85273, -33.8994, -33.94667, -33.99393, -34.04068, -34.08667, 
        -34.13155, -34.1757, -34.21896, -34.26168, -34.30389, -34.34576, 
        -34.3873, -34.42858, -34.4698, -34.50976, -34.55095, -34.59251, 
        -34.63456, -34.67738, -34.72048, -34.764, -34.80748, -34.85096, 
        -34.89414, -34.93693, -34.9796, -35.02227, -35.06496, -35.10828, 
        -35.15213, -35.1952, -35.23925, -35.28285, -35.32594, -35.3686, 
        -35.41123, -35.45387, -35.49665, -35.53953, -35.5825, -35.62574, 
        -35.6694, -35.71349, -35.75795, -35.80268, -35.84758, -35.89164, 
        -35.93702, -35.98282, -36.02931, -36.07674, -36.12486, -36.17412, 
        -36.22425, -36.27575, -36.32782, -36.38, -36.43135, -36.48154, 
        -36.53044, -36.57817, -36.62494, -36.67102, -36.71547, -36.76032, 
        -36.80428, -36.84749, -36.89002, -36.93201, -36.97339, -37.01429, 
        -37.05457, -37.09471, -37.13527, -37.17608, -37.21682, -37.25704, 
        -37.29613, -37.33405, -37.37087, -37.40685, -37.44127, -37.47612, 
        -37.51015, -37.543, -37.57433, -37.60381, -37.63172, -37.65868, 
        -37.68513, -37.71099, -37.73635, -37.76077, -37.78394, -37.80569, 
        -37.82647, -37.84572, -37.86381, -37.88109, -37.89794, -37.91481, 
        -37.93093, -37.94799, -37.96464, -37.98058, -37.99597, -38.01101, 
        -38.02615, -38.04207, -38.05906, -38.07757, -38.09771, -38.11963, 
        -38.14307, -38.16742, -38.19183, -38.21572, -38.23894, -38.26165, 
        -38.28429, -38.30713, -38.32935, -38.35268, -38.37606, -38.39943, 
        -38.42307, -38.44725, -38.47213, -38.49733, -38.52226, -38.54642, 
        -38.56909, -38.59013, -38.60968, -38.62813, -38.64585, -38.66341, 
        -38.68106, -38.69928, -38.71823, -38.73778, -38.75798, -38.77842, 
        -38.79917, -38.81886, -38.83955, -38.85972, -38.87954, -38.89917, 
        -38.91916, -38.94016, -38.9627, -38.98712, -39.01334, -39.04071, 
        -39.06897, -39.0976, -39.12633, -39.15519, -39.18425, -39.21356, 
        -39.243, -39.2722, -39.30152, -39.33112, -39.36139, -39.39228, 
        -39.42365, -39.4544, -39.48258, -39.51019, -39.53606, -39.56053, 
        -39.58397, -39.60657, -39.62856, -39.65012, -39.67141, -39.69269, 
        -39.7134, -39.73384, -39.75293, -39.77045, -39.78593, -39.79895, 
        -39.80942, -39.8175, -39.82357, -39.82805, -39.83118, -39.83353, 
        -39.83504, -39.83579, -39.83552, -39.83401, -39.83094, -39.82523, 
        -39.81961, -39.81362, -39.80779, -39.80272, -39.7997, -39.80013, 
        -39.8053, -39.81676, -39.83509, -39.86065, -39.89233, -39.92875, 
        -39.96775, -40.00748, -40.04669, -40.08417, -40.11936, -40.15257, 
        -40.18377, -40.21341, -40.24183, -40.26954, -40.29682, -40.32339, 
        -40.3486, -40.37219, -40.39399, -40.41412, -40.433, -40.45123, 
        -40.46907, -40.48687, -40.50352, -40.5207, -40.5372, -40.5525, 
        -40.56629, -40.57831, -40.58887, -40.59835, -40.60758, -40.61719, 
        -40.62734, -40.63813, -40.64942, -40.66096, -40.67226, -40.68354, 
        -40.69417, -40.70444, -40.71376, -40.72202, -40.72921, -40.73547, 
        -40.74088, -40.74554, -40.74958, -40.75286, -40.7553, -40.75653, 
        -40.75605, -40.75342, -40.74871, -40.74193, -40.73323, -40.72254, 
        -40.7099, -40.69526, -40.67862, -40.65948, -40.63734, -40.61133, 
        -40.58037, -40.54401, -40.50057, -40.45207, -40.39753, -40.33776, 
        -40.2733, -40.20457, -40.13239, -40.05601, -39.97522, -39.88886, 
        -39.79697,
  -32.98809, -33.03534, -33.08141, -33.12599, -33.16906, -33.21082, 
        -33.25164, -33.2921, -33.33253, -33.37309, -33.4137, -33.45417, 
        -33.49441, -33.53359, -33.57411, -33.61557, -33.65841, -33.70293, 
        -33.7489, -33.7959, -33.84301, -33.88994, -33.93641, -33.98207, 
        -34.02715, -34.07139, -34.11518, -34.15877, -34.20037, -34.24289, 
        -34.28502, -34.32668, -34.36794, -34.40892, -34.44982, -34.49143, 
        -34.5335, -34.57664, -34.62059, -34.66489, -34.70936, -34.75356, 
        -34.79755, -34.84116, -34.88344, -34.92608, -34.96876, -35.01178, 
        -35.05518, -35.09882, -35.14238, -35.18559, -35.22836, -35.27088, 
        -35.31348, -35.35626, -35.39925, -35.44239, -35.48565, -35.52916, 
        -35.57203, -35.61637, -35.66112, -35.70633, -35.7518, -35.79755, 
        -35.84368, -35.89033, -35.93771, -35.98581, -36.03461, -36.08442, 
        -36.13516, -36.18692, -36.23962, -36.29239, -36.34446, -36.39431, 
        -36.44392, -36.49239, -36.53988, -36.58669, -36.63286, -36.67809, 
        -36.72258, -36.7664, -36.80935, -36.85184, -36.89385, -36.93491, 
        -36.97548, -37.01579, -37.05633, -37.09737, -37.13717, -37.17766, 
        -37.21712, -37.25551, -37.29293, -37.32958, -37.36574, -37.40123, 
        -37.43578, -37.4688, -37.49992, -37.52885, -37.55605, -37.58221, 
        -37.60809, -37.6333, -37.65812, -37.68224, -37.70533, -37.72618, 
        -37.74693, -37.76645, -37.7847, -37.8021, -37.81898, -37.83601, 
        -37.85324, -37.87053, -37.88737, -37.90346, -37.91899, -37.93435, 
        -37.95004, -37.9666, -37.98422, -38.00322, -38.02404, -38.04671, 
        -38.07102, -38.09526, -38.12062, -38.14543, -38.16941, -38.19267, 
        -38.21551, -38.23825, -38.26095, -38.28366, -38.30648, -38.32919, 
        -38.35226, -38.37599, -38.40065, -38.42594, -38.45121, -38.47581, 
        -38.49923, -38.52127, -38.54193, -38.56144, -38.5801, -38.59735, 
        -38.61551, -38.634, -38.65307, -38.67281, -38.69317, -38.71405, 
        -38.73523, -38.75677, -38.77802, -38.79897, -38.81923, -38.83903, 
        -38.85899, -38.87985, -38.90232, -38.92688, -38.95328, -38.98089, 
        -39.00969, -39.03907, -39.06866, -39.09847, -39.1283, -39.15711, 
        -39.18674, -39.21591, -39.24486, -39.27411, -39.30387, -39.33454, 
        -39.36547, -39.39537, -39.42372, -39.45049, -39.47574, -39.49992, 
        -39.52316, -39.54575, -39.5678, -39.58969, -39.61154, -39.6331, 
        -39.65414, -39.67455, -39.69343, -39.71056, -39.72554, -39.73822, 
        -39.7486, -39.7568, -39.76213, -39.76696, -39.77059, -39.77325, 
        -39.77515, -39.77611, -39.77593, -39.77429, -39.77108, -39.76604, 
        -39.7597, -39.75302, -39.74664, -39.74165, -39.73909, -39.74053, 
        -39.74726, -39.76069, -39.78113, -39.80863, -39.8423, -39.88018, 
        -39.92075, -39.96201, -40.00255, -40.04118, -40.0773, -40.11126, 
        -40.14293, -40.17307, -40.20188, -40.22903, -40.25633, -40.28279, 
        -40.30794, -40.33149, -40.35313, -40.37321, -40.3921, -40.41036, 
        -40.42832, -40.4462, -40.46394, -40.48135, -40.49798, -40.51335, 
        -40.52697, -40.53895, -40.54921, -40.55841, -40.56726, -40.57623, 
        -40.58575, -40.59589, -40.60669, -40.61792, -40.62946, -40.6411, 
        -40.65258, -40.66348, -40.67338, -40.68199, -40.68907, -40.6949, 
        -40.69972, -40.70366, -40.70702, -40.70963, -40.71186, -40.71166, 
        -40.71091, -40.70811, -40.70333, -40.69631, -40.68713, -40.6758, 
        -40.66245, -40.64698, -40.62983, -40.61063, -40.58872, -40.56342, 
        -40.53364, -40.49844, -40.45726, -40.41014, -40.35701, -40.29868, 
        -40.23621, -40.16964, -40.09929, -40.02587, -39.94773, -39.8647, 
        -39.77594,
  -32.88085, -32.9282, -32.97455, -33.01944, -33.0628, -33.10463, 
        -33.1455, -33.18591, -33.22636, -33.26588, -33.30661, -33.34734, 
        -33.38793, -33.42856, -33.46968, -33.51186, -33.55546, -33.60054, 
        -33.64674, -33.69361, -33.74036, -33.78672, -33.83269, -33.87737, 
        -33.92257, -33.96754, -34.01219, -34.05642, -34.10021, -34.14358, 
        -34.18631, -34.22835, -34.26962, -34.3104, -34.35131, -34.39271, 
        -34.43509, -34.47864, -34.52218, -34.56731, -34.61246, -34.65742, 
        -34.70206, -34.74609, -34.78955, -34.83231, -34.87479, -34.91736, 
        -34.96016, -35.00323, -35.04622, -35.08894, -35.13138, -35.17376, 
        -35.21528, -35.2582, -35.30144, -35.34489, -35.38847, -35.4323, 
        -35.47657, -35.5212, -35.56631, -35.61198, -35.65812, -35.70471, 
        -35.75181, -35.79953, -35.84797, -35.89703, -35.94651, -35.99577, 
        -36.04684, -36.099, -36.15208, -36.20523, -36.25774, -36.30924, 
        -36.35958, -36.40882, -36.45716, -36.5048, -36.55169, -36.59737, 
        -36.64243, -36.68671, -36.73044, -36.77349, -36.81598, -36.85666, 
        -36.89752, -36.93783, -36.9782, -37.01881, -37.05952, -37.10008, 
        -37.13985, -37.1787, -37.2167, -37.25402, -37.29082, -37.32685, 
        -37.36175, -37.39477, -37.42566, -37.45424, -37.48085, -37.50542, 
        -37.53049, -37.55517, -37.57943, -37.60324, -37.62631, -37.64838, 
        -37.6694, -37.68911, -37.70756, -37.72507, -37.74212, -37.75914, 
        -37.77642, -37.79377, -37.81062, -37.82677, -37.84244, -37.85813, 
        -37.8743, -37.89043, -37.90878, -37.92849, -37.94992, -37.97323, 
        -37.99816, -38.02406, -38.05009, -38.07568, -38.10043, -38.12438, 
        -38.14769, -38.17056, -38.19307, -38.2154, -38.23765, -38.25957, 
        -38.28225, -38.30566, -38.33025, -38.35545, -38.37995, -38.405, 
        -38.42915, -38.45223, -38.47411, -38.49487, -38.51461, -38.53363, 
        -38.55225, -38.57102, -38.59024, -38.61014, -38.63067, -38.65215, 
        -38.67416, -38.69642, -38.71865, -38.74034, -38.76105, -38.7811, 
        -38.80104, -38.82176, -38.84399, -38.86713, -38.89341, -38.92115, 
        -38.95021, -38.98016, -39.0105, -39.0411, -39.07169, -39.10194, 
        -39.13155, -39.16053, -39.18915, -39.21791, -39.24719, -39.27725, 
        -39.30737, -39.33679, -39.36454, -39.39038, -39.41513, -39.43885, 
        -39.46204, -39.48468, -39.50706, -39.52948, -39.55164, -39.57236, 
        -39.59377, -39.61396, -39.6325, -39.64912, -39.6637, -39.67622, 
        -39.68671, -39.69542, -39.70226, -39.70769, -39.71195, -39.71502, 
        -39.71711, -39.71823, -39.71815, -39.71659, -39.71322, -39.70798, 
        -39.7013, -39.69423, -39.68768, -39.68297, -39.68117, -39.68407, 
        -39.69283, -39.7084, -39.73105, -39.76049, -39.79463, -39.83396, 
        -39.87551, -39.91766, -39.95894, -39.99821, -40.03499, -40.06927, 
        -40.10159, -40.13219, -40.16136, -40.18984, -40.21733, -40.24399, 
        -40.26906, -40.29258, -40.31442, -40.33474, -40.35393, -40.37225, 
        -40.39035, -40.40819, -40.42597, -40.44323, -40.45979, -40.47482, 
        -40.48827, -40.5, -40.51011, -40.51917, -40.52777, -40.53635, 
        -40.54548, -40.55508, -40.56543, -40.5752, -40.5865, -40.59827, 
        -40.61, -40.6212, -40.63135, -40.63995, -40.6468, -40.65237, 
        -40.65665, -40.66005, -40.66275, -40.66496, -40.66646, -40.66692, 
        -40.66574, -40.66269, -40.65743, -40.65, -40.6403, -40.62832, 
        -40.61441, -40.59826, -40.58055, -40.56113, -40.53954, -40.51469, 
        -40.48573, -40.45175, -40.41192, -40.3662, -40.31507, -40.25875, 
        -40.19833, -40.13403, -40.06639, -39.99543, -39.92039, -39.84049, 
        -39.75515,
  -32.77609, -32.82323, -32.86956, -32.91462, -32.95708, -32.99916, 
        -33.04024, -33.08084, -33.12144, -33.16219, -33.20313, -33.24413, 
        -33.2851, -33.32619, -33.36784, -33.41058, -33.45465, -33.49997, 
        -33.54509, -33.59143, -33.63754, -33.68328, -33.72883, -33.77439, 
        -33.82005, -33.8658, -33.91142, -33.95675, -34.00171, -34.04617, 
        -34.0899, -34.13266, -34.17435, -34.21423, -34.25488, -34.29627, 
        -34.33873, -34.3825, -34.42731, -34.47267, -34.51815, -34.56352, 
        -34.60855, -34.65298, -34.69657, -34.73932, -34.78151, -34.82359, 
        -34.86579, -34.90718, -34.94961, -34.99195, -35.03406, -35.07631, 
        -35.11889, -35.16185, -35.20528, -35.24903, -35.29301, -35.33728, 
        -35.38196, -35.42714, -35.47284, -35.51911, -35.56597, -35.6134, 
        -35.66047, -35.70924, -35.75871, -35.80873, -35.85913, -35.90999, 
        -35.96159, -36.01417, -36.06743, -36.12091, -36.17392, -36.22602, 
        -36.27702, -36.327, -36.37606, -36.42427, -36.47157, -36.51686, 
        -36.56228, -36.60702, -36.65126, -36.69505, -36.73819, -36.7804, 
        -36.82156, -36.86194, -36.90207, -36.94235, -36.98288, -37.02335, 
        -37.06339, -37.10272, -37.14132, -37.17927, -37.21655, -37.25188, 
        -37.28678, -37.3197, -37.35028, -37.37848, -37.40472, -37.4297, 
        -37.45404, -37.47821, -37.5021, -37.52572, -37.54884, -37.57116, 
        -37.59253, -37.61265, -37.63149, -37.64922, -37.66638, -37.68343, 
        -37.69969, -37.71688, -37.7337, -37.74991, -37.76575, -37.78177, 
        -37.7985, -37.81627, -37.83527, -37.85565, -37.87766, -37.90144, 
        -37.92677, -37.95307, -37.97955, -38.00562, -38.03098, -38.05555, 
        -38.07953, -38.10283, -38.12554, -38.14676, -38.16863, -38.19046, 
        -38.21278, -38.236, -38.26026, -38.28544, -38.31093, -38.33625, 
        -38.36103, -38.38503, -38.40804, -38.42993, -38.45072, -38.47053, 
        -38.48972, -38.50887, -38.5284, -38.54861, -38.56973, -38.59185, 
        -38.61478, -38.63715, -38.66037, -38.68282, -38.70411, -38.72435, 
        -38.7442, -38.76459, -38.78629, -38.81007, -38.83578, -38.86345, 
        -38.89264, -38.92295, -38.95396, -38.98526, -39.0165, -39.0469, 
        -39.07645, -39.10513, -39.13334, -39.16164, -39.19045, -39.2198, 
        -39.24918, -39.27792, -39.30405, -39.32968, -39.35402, -39.37748, 
        -39.40052, -39.42334, -39.44607, -39.4688, -39.49125, -39.51331, 
        -39.53456, -39.55445, -39.57259, -39.58877, -39.60302, -39.61548, 
        -39.62626, -39.63535, -39.64286, -39.64892, -39.65367, -39.65723, 
        -39.65972, -39.66111, -39.66121, -39.65968, -39.6563, -39.6511, 
        -39.64368, -39.63675, -39.63056, -39.62652, -39.62615, -39.63081, 
        -39.64182, -39.65953, -39.68416, -39.7153, -39.7516, -39.79156, 
        -39.8336, -39.87616, -39.91771, -39.95732, -39.99432, -40.02886, 
        -40.06134, -40.09214, -40.12181, -40.15061, -40.17838, -40.20515, 
        -40.23051, -40.25448, -40.27679, -40.29769, -40.31732, -40.33598, 
        -40.35402, -40.37172, -40.38914, -40.40499, -40.42106, -40.43584, 
        -40.44891, -40.46039, -40.47035, -40.47942, -40.488, -40.49654, 
        -40.50535, -40.51472, -40.52439, -40.53476, -40.54565, -40.55702, 
        -40.56848, -40.57942, -40.58924, -40.59757, -40.60415, -40.60937, 
        -40.61327, -40.61625, -40.61856, -40.62031, -40.62146, -40.62141, 
        -40.61967, -40.616, -40.6102, -40.6022, -40.59185, -40.57939, 
        -40.56482, -40.54827, -40.53026, -40.51068, -40.48914, -40.46473, 
        -40.43659, -40.4037, -40.3654, -40.32053, -40.2713, -40.2174, 
        -40.15936, -40.09769, -40.03267, -39.96416, -39.89165, -39.81435, 
        -39.73204,
  -32.67297, -32.71976, -32.76571, -32.8106, -32.85414, -32.8964, 
        -32.93776, -32.97862, -33.01965, -33.06053, -33.10164, -33.14285, 
        -33.18429, -33.22582, -33.26694, -33.3103, -33.35476, -33.40015, 
        -33.44598, -33.49166, -33.53691, -33.58202, -33.62722, -33.67286, 
        -33.71905, -33.76572, -33.81236, -33.85878, -33.90488, -33.9495, 
        -33.99428, -34.03786, -34.08014, -34.12125, -34.16215, -34.20351, 
        -34.24604, -34.28988, -34.33474, -34.3801, -34.42569, -34.4712, 
        -34.51639, -34.5609, -34.60349, -34.64608, -34.68795, -34.72946, 
        -34.77097, -34.81268, -34.85457, -34.89657, -34.93856, -34.98086, 
        -35.02346, -35.06651, -35.11012, -35.15411, -35.19852, -35.24325, 
        -35.28758, -35.33339, -35.37976, -35.4267, -35.47439, -35.52267, 
        -35.5719, -35.62186, -35.67252, -35.72365, -35.77499, -35.82655, 
        -35.87863, -35.93153, -35.98514, -36.03898, -36.09249, -36.14412, 
        -36.19567, -36.24619, -36.29572, -36.34428, -36.39183, -36.43841, 
        -36.48405, -36.52922, -36.57401, -36.61849, -36.66227, -36.7051, 
        -36.74668, -36.78724, -36.82728, -36.86725, -36.90752, -36.94685, 
        -36.98703, -37.02675, -37.06585, -37.10423, -37.14177, -37.1781, 
        -37.21267, -37.24528, -37.27569, -37.30362, -37.3297, -37.35437, 
        -37.37833, -37.4019, -37.42545, -37.44885, -37.47211, -37.49472, 
        -37.51538, -37.53591, -37.55525, -37.57343, -37.59087, -37.60805, 
        -37.62514, -37.64231, -37.65901, -37.67529, -37.69141, -37.70779, 
        -37.72504, -37.74335, -37.76286, -37.78375, -37.80614, -37.83024, 
        -37.85575, -37.88216, -37.90774, -37.93408, -37.9599, -37.98517, 
        -38.00986, -38.03378, -38.05692, -38.07935, -38.10131, -38.1231, 
        -38.1455, -38.16873, -38.19299, -38.21793, -38.24332, -38.26872, 
        -38.29387, -38.31857, -38.34253, -38.3654, -38.38704, -38.40771, 
        -38.42659, -38.44627, -38.46624, -38.48691, -38.50862, -38.53151, 
        -38.55542, -38.57989, -38.6042, -38.62757, -38.64955, -38.67019, 
        -38.69013, -38.71028, -38.73156, -38.75469, -38.78004, -38.80749, 
        -38.83647, -38.86703, -38.89867, -38.93029, -38.96184, -38.99227, 
        -39.02054, -39.04885, -39.07668, -39.10469, -39.13311, -39.16201, 
        -39.19091, -39.21906, -39.24602, -39.27153, -39.29585, -39.31917, 
        -39.34221, -39.36505, -39.38797, -39.41085, -39.43348, -39.45548, 
        -39.47636, -39.49573, -39.51324, -39.5289, -39.54282, -39.55533, 
        -39.56649, -39.57616, -39.5843, -39.59, -39.59535, -39.59946, 
        -39.60239, -39.60408, -39.6044, -39.60306, -39.59989, -39.59502, 
        -39.58894, -39.5826, -39.57728, -39.57445, -39.57598, -39.58277, 
        -39.59589, -39.61576, -39.64228, -39.6749, -39.71199, -39.75238, 
        -39.79463, -39.83694, -39.8783, -39.91779, -39.95467, -39.98919, 
        -40.02162, -40.05255, -40.08245, -40.11152, -40.13847, -40.16543, 
        -40.1912, -40.21587, -40.23899, -40.26069, -40.28085, -40.2998, 
        -40.31773, -40.33504, -40.35195, -40.36809, -40.38349, -40.39766, 
        -40.41041, -40.42177, -40.4319, -40.44115, -40.44993, -40.45856, 
        -40.46728, -40.47628, -40.48575, -40.49552, -40.50586, -40.51666, 
        -40.52735, -40.53738, -40.54641, -40.554, -40.56012, -40.56492, 
        -40.56859, -40.5715, -40.57351, -40.57496, -40.57558, -40.57491, 
        -40.57145, -40.56707, -40.56057, -40.55182, -40.54103, -40.52818, 
        -40.51339, -40.49659, -40.4784, -40.45877, -40.43722, -40.41322, 
        -40.38566, -40.35385, -40.31702, -40.27501, -40.22813, -40.17676, 
        -40.12135, -40.06236, -39.99967, -39.93318, -39.8624, -39.78709, 
        -39.70698,
  -32.57288, -32.61924, -32.66479, -32.70938, -32.75285, -32.79548, 
        -32.8373, -32.87878, -32.92015, -32.9605, -33.0017, -33.0429, 
        -33.0846, -33.1263, -33.169, -33.21275, -33.25742, -33.3027, 
        -33.34804, -33.39296, -33.43748, -33.48211, -33.52708, -33.57287, 
        -33.6186, -33.66593, -33.71351, -33.76096, -33.80801, -33.85472, 
        -33.90067, -33.9451, -33.98833, -34.03016, -34.07137, -34.11297, 
        -34.15556, -34.1993, -34.2439, -34.28813, -34.33357, -34.37893, 
        -34.42404, -34.46867, -34.51211, -34.55458, -34.59609, -34.63705, 
        -34.67785, -34.71886, -34.76023, -34.80194, -34.84398, -34.88631, 
        -34.92914, -34.97149, -35.01537, -35.05973, -35.10463, -35.15, 
        -35.19604, -35.24262, -35.28979, -35.33758, -35.38597, -35.43516, 
        -35.48528, -35.53624, -35.58804, -35.64021, -35.69241, -35.74369, 
        -35.79646, -35.85006, -35.90427, -35.95877, -36.01284, -36.06592, 
        -36.1177, -36.16835, -36.21795, -36.26649, -36.31419, -36.36087, 
        -36.40675, -36.45239, -36.49771, -36.54253, -36.58714, -36.62952, 
        -36.67149, -36.71241, -36.75251, -36.79238, -36.83243, -36.8727, 
        -36.91288, -36.95286, -36.99228, -37.03092, -37.06845, -37.10464, 
        -37.13884, -37.17093, -37.20106, -37.22901, -37.25492, -37.27938, 
        -37.30197, -37.32517, -37.34842, -37.37169, -37.39508, -37.41784, 
        -37.43995, -37.46091, -37.48054, -37.49908, -37.51684, -37.53419, 
        -37.55144, -37.56861, -37.58551, -37.60208, -37.61861, -37.63553, 
        -37.65326, -37.67102, -37.69089, -37.71198, -37.7345, -37.75861, 
        -37.78409, -37.81036, -37.83694, -37.8634, -37.88958, -37.91552, 
        -37.94088, -37.96545, -37.98928, -38.01226, -38.03472, -38.0571, 
        -38.07986, -38.10336, -38.12757, -38.15236, -38.17746, -38.20174, 
        -38.22696, -38.252, -38.2765, -38.30009, -38.32253, -38.34392, 
        -38.36456, -38.38493, -38.40556, -38.42695, -38.44923, -38.47288, 
        -38.49773, -38.52322, -38.54852, -38.57283, -38.59562, -38.61689, 
        -38.63718, -38.6573, -38.67818, -38.70071, -38.72438, -38.75134, 
        -38.78056, -38.81124, -38.84306, -38.87526, -38.90681, -38.93694, 
        -38.96598, -38.99401, -39.0216, -39.04935, -39.07757, -39.10617, 
        -39.1347, -39.16274, -39.18978, -39.21547, -39.23989, -39.26341, 
        -39.28637, -39.30919, -39.33207, -39.35487, -39.37732, -39.39893, 
        -39.41819, -39.43682, -39.45363, -39.46882, -39.48264, -39.49517, 
        -39.50661, -39.51674, -39.52551, -39.53273, -39.53873, -39.5435, 
        -39.54694, -39.54895, -39.54961, -39.54858, -39.54578, -39.54147, 
        -39.53618, -39.53088, -39.52694, -39.52594, -39.5294, -39.53844, 
        -39.5538, -39.57579, -39.60396, -39.6376, -39.67538, -39.71495, 
        -39.75686, -39.79889, -39.83965, -39.87842, -39.91492, -39.94913, 
        -39.9816, -40.01256, -40.04243, -40.07135, -40.09949, -40.12661, 
        -40.1529, -40.17851, -40.20255, -40.22501, -40.24581, -40.26496, 
        -40.28274, -40.2995, -40.31565, -40.33101, -40.34556, -40.35907, 
        -40.3715, -40.38284, -40.3932, -40.40279, -40.41186, -40.42067, 
        -40.42944, -40.4383, -40.44739, -40.45677, -40.46548, -40.47529, 
        -40.48495, -40.49377, -40.50166, -40.50837, -40.51386, -40.51828, 
        -40.52183, -40.52449, -40.52649, -40.52769, -40.528, -40.52666, 
        -40.5236, -40.51844, -40.51119, -40.50177, -40.49051, -40.47738, 
        -40.46255, -40.44592, -40.42767, -40.40771, -40.38624, -40.3625, 
        -40.33561, -40.30489, -40.26952, -40.22943, -40.18476, -40.13589, 
        -40.08294, -40.02612, -39.96511, -39.90023, -39.8309, -39.75661, 
        -39.6777,
  -32.47506, -32.52074, -32.56576, -32.60994, -32.65227, -32.69514, 
        -32.73773, -32.77998, -32.82198, -32.86374, -32.90525, -32.94659, 
        -32.9882, -33.03022, -33.0731, -33.11694, -33.16159, -33.20653, 
        -33.2513, -33.29458, -33.33854, -33.38268, -33.42768, -33.47367, 
        -33.52077, -33.56862, -33.61689, -33.66497, -33.71291, -33.76061, 
        -33.80748, -33.85323, -33.89724, -33.94009, -33.98107, -34.02307, 
        -34.06577, -34.10938, -34.15368, -34.19849, -34.24352, -34.28867, 
        -34.33371, -34.37794, -34.42135, -34.4637, -34.50504, -34.54555, 
        -34.58576, -34.62614, -34.666, -34.7075, -34.74955, -34.79214, 
        -34.83527, -34.87903, -34.92332, -34.96823, -35.01379, -35.05999, 
        -35.10685, -35.15427, -35.2023, -35.25092, -35.29997, -35.3498, 
        -35.39955, -35.45143, -35.50407, -35.55685, -35.60975, -35.66331, 
        -35.71693, -35.77146, -35.82661, -35.88195, -35.93661, -35.98996, 
        -36.04178, -36.09219, -36.14149, -36.18978, -36.23727, -36.28301, 
        -36.32923, -36.37506, -36.42104, -36.46679, -36.51144, -36.5555, 
        -36.5981, -36.63941, -36.67979, -36.71968, -36.75978, -36.79978, 
        -36.83985, -36.87982, -36.91935, -36.95808, -36.99556, -37.0304, 
        -37.06434, -37.09634, -37.12609, -37.15367, -37.17949, -37.20388, 
        -37.22721, -37.2501, -37.27319, -37.29648, -37.31967, -37.34258, 
        -37.36465, -37.38601, -37.40592, -37.42485, -37.44308, -37.46085, 
        -37.47842, -37.49486, -37.51211, -37.5292, -37.54634, -37.56395, 
        -37.58223, -37.60138, -37.62139, -37.64247, -37.66489, -37.68879, 
        -37.71398, -37.74001, -37.76644, -37.79305, -37.81965, -37.84616, 
        -37.87228, -37.89773, -37.92232, -37.94504, -37.96824, -37.99139, 
        -38.0148, -38.0387, -38.06304, -38.0877, -38.11249, -38.13752, 
        -38.16259, -38.18764, -38.21236, -38.23641, -38.25948, -38.28164, 
        -38.30312, -38.32427, -38.34576, -38.36788, -38.39062, -38.41487, 
        -38.44047, -38.46672, -38.49173, -38.51689, -38.54065, -38.56279, 
        -38.58367, -38.60393, -38.62453, -38.64646, -38.67052, -38.69711, 
        -38.7263, -38.75744, -38.78954, -38.8218, -38.85307, -38.8833, 
        -38.91217, -38.93999, -38.96737, -38.99495, -39.02308, -39.05146, 
        -39.07985, -39.10794, -39.13525, -39.16047, -39.18529, -39.20895, 
        -39.23192, -39.2545, -39.277, -39.29932, -39.3213, -39.34214, 
        -39.3615, -39.37932, -39.39553, -39.4104, -39.42416, -39.43694, 
        -39.44861, -39.45918, -39.4682, -39.47607, -39.48283, -39.48811, 
        -39.49226, -39.49484, -39.4958, -39.49529, -39.49307, -39.48952, 
        -39.48523, -39.48035, -39.47821, -39.4794, -39.48522, -39.49665, 
        -39.5141, -39.53768, -39.56711, -39.60154, -39.63978, -39.68055, 
        -39.72219, -39.76345, -39.80332, -39.84123, -39.87713, -39.91098, 
        -39.9433, -39.97411, -40.00374, -40.03243, -40.06026, -40.08776, 
        -40.11478, -40.14134, -40.1663, -40.18955, -40.21095, -40.2303, 
        -40.24785, -40.26409, -40.27918, -40.29345, -40.30602, -40.3189, 
        -40.33109, -40.34253, -40.35319, -40.36311, -40.37246, -40.38146, 
        -40.39041, -40.39922, -40.4082, -40.41713, -40.42608, -40.43488, 
        -40.44329, -40.45096, -40.45765, -40.46344, -40.46832, -40.47229, 
        -40.47562, -40.47812, -40.47994, -40.48111, -40.48098, -40.47924, 
        -40.47548, -40.46956, -40.46156, -40.4516, -40.43999, -40.42663, 
        -40.41175, -40.39508, -40.37685, -40.35728, -40.33586, -40.31234, 
        -40.28597, -40.25616, -40.22218, -40.18384, -40.14014, -40.09336, 
        -40.04229, -39.98709, -39.92763, -39.8635, -39.79458, -39.72105, 
        -39.64289,
  -32.37815, -32.4233, -32.4677, -32.51148, -32.55478, -32.59781, 
        -32.64093, -32.68401, -32.7268, -32.76917, -32.81103, -32.85262, 
        -32.89428, -32.93644, -32.97832, -33.02216, -33.06645, -33.11097, 
        -33.15514, -33.19894, -33.24252, -33.2865, -33.33133, -33.37775, 
        -33.42515, -33.47329, -33.522, -33.57067, -33.61908, -33.66641, 
        -33.71404, -33.76059, -33.80572, -33.8495, -33.89245, -33.93505, 
        -33.97787, -34.0215, -34.06549, -34.11003, -34.1548, -34.19963, 
        -34.2441, -34.28825, -34.33036, -34.37256, -34.41379, -34.4541, 
        -34.494, -34.53387, -34.57447, -34.61572, -34.65783, -34.70063, 
        -34.74415, -34.78831, -34.83324, -34.8789, -34.92531, -34.97241, 
        -35.02013, -35.06746, -35.11625, -35.16541, -35.21511, -35.2655, 
        -35.31674, -35.36894, -35.42217, -35.47554, -35.52959, -35.58382, 
        -35.63849, -35.69436, -35.7506, -35.80668, -35.86181, -35.91421, 
        -35.96587, -36.016, -36.06493, -36.11287, -36.16018, -36.2071, 
        -36.25361, -36.29987, -36.34628, -36.39267, -36.43822, -36.48245, 
        -36.52599, -36.5677, -36.60835, -36.64839, -36.6883, -36.72694, 
        -36.76701, -36.80678, -36.84604, -36.88454, -36.92192, -36.95748, 
        -36.9913, -37.02298, -37.05259, -37.08019, -37.10593, -37.13012, 
        -37.15326, -37.17596, -37.19883, -37.22195, -37.24506, -37.26794, 
        -37.28908, -37.31024, -37.33059, -37.34996, -37.36868, -37.38702, 
        -37.40509, -37.42298, -37.44075, -37.45848, -37.47641, -37.49477, 
        -37.51369, -37.53328, -37.55339, -37.57438, -37.59654, -37.62012, 
        -37.64495, -37.6707, -37.69707, -37.72278, -37.74971, -37.77681, 
        -37.80368, -37.82994, -37.85536, -37.87986, -37.90384, -37.92767, 
        -37.95171, -37.97608, -38.00067, -38.02536, -38.05009, -38.07491, 
        -38.09991, -38.12489, -38.14972, -38.17408, -38.19772, -38.22059, 
        -38.24188, -38.26385, -38.28595, -38.30869, -38.33208, -38.35643, 
        -38.38239, -38.40885, -38.43537, -38.46142, -38.48623, -38.50944, 
        -38.53114, -38.55185, -38.57243, -38.59385, -38.61744, -38.64399, 
        -38.67312, -38.70424, -38.73659, -38.76889, -38.80024, -38.83041, 
        -38.85818, -38.88591, -38.91325, -38.94067, -38.96856, -38.99692, 
        -39.02567, -39.05391, -39.08165, -39.10814, -39.13348, -39.15741, 
        -39.18023, -39.20237, -39.22435, -39.24578, -39.26667, -39.28656, 
        -39.30521, -39.3222, -39.33799, -39.35258, -39.36623, -39.37906, 
        -39.3909, -39.40177, -39.41154, -39.41912, -39.42653, -39.43259, 
        -39.43738, -39.44069, -39.44229, -39.44228, -39.44078, -39.4383, 
        -39.43536, -39.43324, -39.43321, -39.43673, -39.44494, -39.4586, 
        -39.47789, -39.50282, -39.53315, -39.56812, -39.60659, -39.64717, 
        -39.68839, -39.72896, -39.76796, -39.8051, -39.84042, -39.87394, 
        -39.90584, -39.93638, -39.96574, -39.99414, -40.021, -40.04865, 
        -40.07628, -40.10334, -40.12918, -40.1531, -40.17508, -40.19457, 
        -40.21185, -40.22726, -40.24136, -40.25459, -40.26727, -40.27961, 
        -40.29162, -40.30327, -40.31427, -40.32463, -40.33437, -40.34369, 
        -40.35283, -40.3618, -40.37035, -40.37885, -40.387, -40.39475, 
        -40.4021, -40.40858, -40.41428, -40.41911, -40.42336, -40.42694, 
        -40.42987, -40.43224, -40.43394, -40.43483, -40.43446, -40.43217, 
        -40.42761, -40.41988, -40.41105, -40.40042, -40.38823, -40.37481, 
        -40.35993, -40.34368, -40.326, -40.30664, -40.28545, -40.26204, 
        -40.23614, -40.20705, -40.17421, -40.13714, -40.09595, -40.05061, 
        -40.00101, -39.94681, -39.88799, -39.82421, -39.75556, -39.6821, 
        -39.60418,
  -32.28439, -32.32901, -32.37273, -32.41592, -32.45901, -32.50222, 
        -32.54573, -32.58952, -32.63318, -32.6753, -32.71782, -32.75976, 
        -32.80158, -32.84399, -32.88698, -32.93053, -32.9745, -33.01839, 
        -33.06192, -33.10521, -33.14843, -33.19231, -33.2374, -33.28393, 
        -33.33049, -33.37889, -33.42758, -33.47654, -33.52532, -33.57392, 
        -33.6221, -33.66937, -33.71542, -33.76026, -33.80406, -33.84748, 
        -33.89073, -33.93424, -33.9782, -34.0215, -34.0658, -34.11006, 
        -34.15398, -34.19768, -34.24058, -34.28289, -34.3242, -34.36468, 
        -34.40453, -34.4444, -34.48479, -34.52606, -34.56819, -34.61117, 
        -34.65505, -34.69872, -34.7443, -34.79084, -34.83821, -34.8863, 
        -34.93497, -34.98389, -35.03328, -35.08305, -35.1333, -35.18399, 
        -35.23557, -35.28804, -35.34138, -35.39551, -35.44998, -35.50533, 
        -35.56013, -35.61712, -35.67428, -35.73111, -35.78649, -35.83986, 
        -35.89123, -35.94105, -35.98962, -36.03736, -36.0846, -36.13161, 
        -36.1782, -36.22512, -36.27216, -36.31915, -36.36547, -36.40984, 
        -36.45371, -36.49621, -36.5372, -36.57723, -36.61682, -36.65619, 
        -36.69576, -36.735, -36.77416, -36.81227, -36.8493, -36.88496, 
        -36.91864, -36.95028, -36.97989, -37.00747, -37.03305, -37.05705, 
        -37.07903, -37.10161, -37.12432, -37.14727, -37.17023, -37.19285, 
        -37.21484, -37.23609, -37.25661, -37.27667, -37.29615, -37.31516, 
        -37.33384, -37.35222, -37.37053, -37.38898, -37.40778, -37.42699, 
        -37.44658, -37.4665, -37.48578, -37.50668, -37.52864, -37.55198, 
        -37.57655, -37.60218, -37.6285, -37.6553, -37.68258, -37.71025, 
        -37.73769, -37.76455, -37.79044, -37.81554, -37.84008, -37.86452, 
        -37.88931, -37.91438, -37.93945, -37.96442, -37.98926, -38.01309, 
        -38.03798, -38.063, -38.08797, -38.11266, -38.13683, -38.16045, 
        -38.18353, -38.20619, -38.22895, -38.2518, -38.27534, -38.29956, 
        -38.32512, -38.35168, -38.3787, -38.40555, -38.43148, -38.45589, 
        -38.47855, -38.4999, -38.52064, -38.5422, -38.56425, -38.59045, 
        -38.61963, -38.65101, -38.68357, -38.71577, -38.74712, -38.77723, 
        -38.80601, -38.8338, -38.86104, -38.88831, -38.91599, -38.94425, 
        -38.97325, -39.00199, -39.03014, -39.05706, -39.0826, -39.10661, 
        -39.12908, -39.1508, -39.1719, -39.19242, -39.21188, -39.23064, 
        -39.24714, -39.26377, -39.27914, -39.29365, -39.30723, -39.32005, 
        -39.33202, -39.34307, -39.35327, -39.36263, -39.37101, -39.37822, 
        -39.38406, -39.38818, -39.39066, -39.39142, -39.39103, -39.3897, 
        -39.38847, -39.38828, -39.39056, -39.39661, -39.40716, -39.42263, 
        -39.44352, -39.46966, -39.50058, -39.53575, -39.57418, -39.61448, 
        -39.65429, -39.69418, -39.73241, -39.76882, -39.80345, -39.83662, 
        -39.86832, -39.89855, -39.92756, -39.95545, -39.98316, -40.01084, 
        -40.03871, -40.06627, -40.09257, -40.11713, -40.13949, -40.15919, 
        -40.17626, -40.19106, -40.20428, -40.21661, -40.22861, -40.24055, 
        -40.2525, -40.26423, -40.2755, -40.28633, -40.29665, -40.30648, 
        -40.31585, -40.32472, -40.33293, -40.3407, -40.34805, -40.35415, 
        -40.36036, -40.36589, -40.37086, -40.3751, -40.37873, -40.38168, 
        -40.38421, -40.38623, -40.38768, -40.3882, -40.3873, -40.3845, 
        -40.37946, -40.37209, -40.36254, -40.35112, -40.3384, -40.32476, 
        -40.31006, -40.2943, -40.27708, -40.25807, -40.23717, -40.21405, 
        -40.18841, -40.15989, -40.12776, -40.09164, -40.05154, -40.00721, 
        -39.95829, -39.90463, -39.846, -39.78225, -39.71342, -39.6396, 
        -39.56104,
  -32.19228, -32.23653, -32.27985, -32.32256, -32.36535, -32.40757, 
        -32.45139, -32.49565, -32.53991, -32.58369, -32.62668, -32.66912, 
        -32.71147, -32.75426, -32.79737, -32.84094, -32.88466, -32.92807, 
        -32.97107, -33.01295, -33.0561, -33.10004, -33.1452, -33.19168, 
        -33.23928, -33.28773, -33.33646, -33.38536, -33.4342, -33.48292, 
        -33.53128, -33.57899, -33.62567, -33.67116, -33.71455, -33.75852, 
        -33.80225, -33.84616, -33.89028, -33.93449, -33.97845, -34.02213, 
        -34.06561, -34.10874, -34.1515, -34.19376, -34.23523, -34.27604, 
        -34.31624, -34.35632, -34.39586, -34.4372, -34.47953, -34.52282, 
        -34.56706, -34.61231, -34.65857, -34.70594, -34.75424, -34.80326, 
        -34.85263, -34.90213, -34.95209, -35.00231, -35.05289, -35.10415, 
        -35.15519, -35.20816, -35.26202, -35.31645, -35.37156, -35.42736, 
        -35.48424, -35.54169, -35.59963, -35.65665, -35.71207, -35.76514, 
        -35.81627, -35.86603, -35.91468, -35.96244, -36.00964, -36.05671, 
        -36.10302, -36.15051, -36.19824, -36.24574, -36.29281, -36.33898, 
        -36.38378, -36.42678, -36.4681, -36.50807, -36.54748, -36.5866, 
        -36.62547, -36.66426, -36.7028, -36.74068, -36.77761, -36.81322, 
        -36.84604, -36.87785, -36.9074, -36.93473, -36.96006, -36.98384, 
        -37.00664, -37.02911, -37.05173, -37.07459, -37.09742, -37.11992, 
        -37.14179, -37.1631, -37.18401, -37.20458, -37.2249, -37.24463, 
        -37.26394, -37.28178, -37.30068, -37.31979, -37.33935, -37.35929, 
        -37.37951, -37.39983, -37.42032, -37.44131, -37.46339, -37.48665, 
        -37.51127, -37.53676, -37.5631, -37.59018, -37.61759, -37.64549, 
        -37.67319, -37.70029, -37.72659, -37.75198, -37.77591, -37.80099, 
        -37.82648, -37.85233, -37.87807, -37.90348, -37.92862, -37.95365, 
        -37.97876, -38.00402, -38.0293, -38.05439, -38.07906, -38.10322, 
        -38.12704, -38.15024, -38.17315, -38.19586, -38.21911, -38.24311, 
        -38.26847, -38.29501, -38.32244, -38.34909, -38.37617, -38.40183, 
        -38.42554, -38.44765, -38.46889, -38.49065, -38.51408, -38.54008, 
        -38.56924, -38.60014, -38.63237, -38.66459, -38.69582, -38.72584, 
        -38.75468, -38.78246, -38.80966, -38.83681, -38.86442, -38.89253, 
        -38.92131, -38.95032, -38.97875, -39.00499, -39.03058, -39.05442, 
        -39.07671, -39.09779, -39.11796, -39.13739, -39.15562, -39.17331, 
        -39.18982, -39.20564, -39.22083, -39.23513, -39.24864, -39.26153, 
        -39.27362, -39.28507, -39.29598, -39.30633, -39.31592, -39.32438, 
        -39.33136, -39.33655, -39.3401, -39.34198, -39.34274, -39.34293, 
        -39.34354, -39.34546, -39.34906, -39.35736, -39.37013, -39.38748, 
        -39.40976, -39.43683, -39.46816, -39.50318, -39.54137, -39.58125, 
        -39.62143, -39.66056, -39.69807, -39.73392, -39.76809, -39.80099, 
        -39.8325, -39.86251, -39.89123, -39.91886, -39.94632, -39.9738, 
        -40.00148, -40.02888, -40.05539, -40.08029, -40.10288, -40.12275, 
        -40.13972, -40.15413, -40.16675, -40.17853, -40.19007, -40.20084, 
        -40.21279, -40.22456, -40.23623, -40.24759, -40.25846, -40.26876, 
        -40.27839, -40.28715, -40.29505, -40.30221, -40.30872, -40.31459, 
        -40.32021, -40.32507, -40.3293, -40.33292, -40.33598, -40.33854, 
        -40.34068, -40.34244, -40.34359, -40.34374, -40.34233, -40.33895, 
        -40.33336, -40.32532, -40.31509, -40.30304, -40.28975, -40.2757, 
        -40.26117, -40.24583, -40.22923, -40.21083, -40.19027, -40.16729, 
        -40.14188, -40.1136, -40.08195, -40.04632, -40.00666, -39.96179, 
        -39.91322, -39.85975, -39.8011, -39.73706, -39.66767, -39.59299, 
        -39.51348,
  -32.10053, -32.14467, -32.18787, -32.23042, -32.27299, -32.3161, 
        -32.35997, -32.4044, -32.44897, -32.49317, -32.5367, -32.57969, 
        -32.6226, -32.66585, -32.70942, -32.75206, -32.79564, -32.8389, 
        -32.88169, -32.92451, -32.96772, -33.01167, -33.05686, -33.10323, 
        -33.15073, -33.19899, -33.24761, -33.29635, -33.34508, -33.39285, 
        -33.44119, -33.48872, -33.53561, -33.5813, -33.62615, -33.67059, 
        -33.71475, -33.75903, -33.80354, -33.84766, -33.89136, -33.93469, 
        -33.97769, -34.02045, -34.06294, -34.10419, -34.14603, -34.18718, 
        -34.22783, -34.26837, -34.30923, -34.35096, -34.39368, -34.4374, 
        -34.48215, -34.52798, -34.57491, -34.62305, -34.6721, -34.72183, 
        -34.77181, -34.82078, -34.87098, -34.92165, -34.97284, -35.02475, 
        -35.07756, -35.13125, -35.18576, -35.24085, -35.29652, -35.35288, 
        -35.41001, -35.46785, -35.52562, -35.58245, -35.63739, -35.69014, 
        -35.74017, -35.79007, -35.83896, -35.88708, -35.93469, -35.98218, 
        -36.02993, -36.07805, -36.12621, -36.17432, -36.22199, -36.2688, 
        -36.31419, -36.35777, -36.39948, -36.43963, -36.47882, -36.51754, 
        -36.55499, -36.59342, -36.63151, -36.66913, -36.70592, -36.74168, 
        -36.77559, -36.80739, -36.83665, -36.86388, -36.88896, -36.9124, 
        -36.93503, -36.95746, -36.98007, -37.00293, -37.02571, -37.04816, 
        -37.0701, -37.09066, -37.11203, -37.1332, -37.15413, -37.17456, 
        -37.1945, -37.21391, -37.23333, -37.25299, -37.27313, -37.29373, 
        -37.31451, -37.33536, -37.35626, -37.3777, -37.40008, -37.42366, 
        -37.4483, -37.47396, -37.50035, -37.52636, -37.55401, -37.58166, 
        -37.60923, -37.63638, -37.66277, -37.68845, -37.71383, -37.73953, 
        -37.76577, -37.79234, -37.81879, -37.8448, -37.87046, -37.89586, 
        -37.92134, -37.94697, -37.97264, -37.99814, -38.02324, -38.04783, 
        -38.07196, -38.0945, -38.11742, -38.14004, -38.16286, -38.18665, 
        -38.21181, -38.23846, -38.26646, -38.29488, -38.32315, -38.34983, 
        -38.37466, -38.39767, -38.41955, -38.44171, -38.4654, -38.49146, 
        -38.52034, -38.55103, -38.58274, -38.61456, -38.64548, -38.67529, 
        -38.70403, -38.73079, -38.75795, -38.785, -38.81244, -38.84048, 
        -38.86911, -38.8979, -38.92619, -38.95323, -38.97853, -39.00217, 
        -39.0241, -39.04467, -39.0641, -39.08245, -39.09964, -39.11615, 
        -39.13191, -39.14718, -39.16193, -39.17596, -39.18946, -39.20225, 
        -39.21453, -39.22654, -39.23834, -39.24986, -39.25992, -39.26992, 
        -39.27839, -39.28504, -39.28988, -39.29317, -39.29536, -39.29715, 
        -39.29954, -39.30368, -39.31054, -39.32096, -39.3356, -39.3546, 
        -39.37802, -39.40564, -39.43723, -39.47235, -39.50985, -39.549, 
        -39.58841, -39.62692, -39.66386, -39.69913, -39.73307, -39.7658, 
        -39.79716, -39.82682, -39.85539, -39.88287, -39.90998, -39.93619, 
        -39.96344, -39.99047, -40.01665, -40.04136, -40.064, -40.08388, 
        -40.10087, -40.11528, -40.12786, -40.13953, -40.1509, -40.16261, 
        -40.17462, -40.18655, -40.19852, -40.21021, -40.2216, -40.23241, 
        -40.24215, -40.25083, -40.25832, -40.26466, -40.27054, -40.27575, 
        -40.28048, -40.28468, -40.28822, -40.29132, -40.29387, -40.29599, 
        -40.29783, -40.29937, -40.30026, -40.30006, -40.29823, -40.29436, 
        -40.28827, -40.27979, -40.26809, -40.25536, -40.24154, -40.2273, 
        -40.21291, -40.19796, -40.18203, -40.16414, -40.1437, -40.12077, 
        -40.0952, -40.06681, -40.03512, -39.99966, -39.96016, -39.91638, 
        -39.86796, -39.81449, -39.75571, -39.69123, -39.6211, -39.54529, 
        -39.46463,
  -32.01072, -32.05515, -32.09851, -32.14124, -32.18386, -32.22696, 
        -32.27081, -32.31521, -32.35981, -32.40418, -32.44708, -32.4906, 
        -32.53413, -32.57796, -32.62199, -32.66599, -32.70963, -32.75284, 
        -32.79571, -32.83869, -32.882, -32.92608, -32.97125, -33.01739, 
        -33.06456, -33.11161, -33.16004, -33.20865, -33.25726, -33.30585, 
        -33.35392, -33.40116, -33.44767, -33.49331, -33.53821, -33.58282, 
        -33.62747, -33.67223, -33.71682, -33.76103, -33.80367, -33.84676, 
        -33.8895, -33.93198, -33.97435, -34.01661, -34.0585, -34.10014, 
        -34.1414, -34.1825, -34.22394, -34.26617, -34.30938, -34.35382, 
        -34.3992, -34.44566, -34.49232, -34.5411, -34.5908, -34.64104, 
        -34.69139, -34.74174, -34.79233, -34.84341, -34.89516, -34.94785, 
        -35.00157, -35.0562, -35.11171, -35.16766, -35.2241, -35.28075, 
        -35.33689, -35.39468, -35.45176, -35.50778, -35.562, -35.61445, 
        -35.66556, -35.71573, -35.7651, -35.814, -35.86216, -35.90999, 
        -35.95832, -36.00685, -36.05532, -36.10372, -36.15155, -36.19864, 
        -36.24345, -36.28751, -36.32966, -36.37012, -36.4094, -36.44801, 
        -36.48634, -36.52454, -36.5624, -36.59967, -36.63638, -36.67216, 
        -36.70605, -36.73795, -36.76684, -36.79361, -36.81834, -36.84166, 
        -36.86432, -36.88592, -36.90871, -36.93173, -36.95464, -36.97719, 
        -36.9994, -37.02135, -37.04313, -37.06491, -37.0865, -37.10746, 
        -37.12797, -37.14782, -37.16768, -37.18781, -37.20844, -37.22957, 
        -37.25097, -37.27236, -37.29298, -37.31509, -37.33815, -37.36221, 
        -37.38742, -37.41329, -37.43969, -37.46651, -37.49369, -37.52097, 
        -37.54815, -37.57498, -37.60125, -37.62724, -37.65318, -37.67963, 
        -37.70661, -37.73391, -37.76104, -37.7877, -37.81384, -37.83979, 
        -37.86479, -37.89083, -37.91674, -37.94256, -37.96802, -37.99283, 
        -38.01713, -38.04087, -38.06371, -38.08623, -38.10903, -38.13259, 
        -38.15788, -38.18493, -38.21339, -38.24286, -38.272, -38.29988, 
        -38.32553, -38.34913, -38.37181, -38.39459, -38.41869, -38.44384, 
        -38.47221, -38.50244, -38.5334, -38.56454, -38.59485, -38.62446, 
        -38.65311, -38.68084, -38.70792, -38.73483, -38.76204, -38.78975, 
        -38.81798, -38.84621, -38.87407, -38.90055, -38.92538, -38.94848, 
        -38.96998, -38.99008, -39.0089, -39.02647, -39.04292, -39.05855, 
        -39.07367, -39.08746, -39.10175, -39.11552, -39.12892, -39.14175, 
        -39.15434, -39.16703, -39.17994, -39.19284, -39.20553, -39.2173, 
        -39.22751, -39.2359, -39.24231, -39.24723, -39.25104, -39.25455, 
        -39.25877, -39.26485, -39.27374, -39.28611, -39.30231, -39.32259, 
        -39.34692, -39.37521, -39.40695, -39.44156, -39.47848, -39.51658, 
        -39.55499, -39.59178, -39.62811, -39.66307, -39.69693, -39.72952, 
        -39.76065, -39.79018, -39.81858, -39.84599, -39.87296, -39.89971, 
        -39.92639, -39.95265, -39.97812, -40.00225, -40.02464, -40.04457, 
        -40.06181, -40.07657, -40.08949, -40.10142, -40.11314, -40.12498, 
        -40.13699, -40.14898, -40.16097, -40.17307, -40.18487, -40.1959, 
        -40.20583, -40.21421, -40.22115, -40.22677, -40.2317, -40.23619, 
        -40.23932, -40.24303, -40.24619, -40.24881, -40.25087, -40.25264, 
        -40.25428, -40.25577, -40.25657, -40.25608, -40.25388, -40.24967, 
        -40.24319, -40.23428, -40.22308, -40.20995, -40.19574, -40.18126, 
        -40.16718, -40.15273, -40.13733, -40.11971, -40.09926, -40.07595, 
        -40.05001, -40.0212, -39.98922, -39.95361, -39.91385, -39.86981, 
        -39.82134, -39.76784, -39.70877, -39.64397, -39.57304, -39.49615, 
        -39.41426,
  -31.92213, -31.96709, -32.011, -32.05413, -32.09699, -32.1391, 
        -32.18276, -32.22696, -32.27144, -32.31587, -32.36005, -32.40405, 
        -32.44812, -32.49245, -32.53698, -32.58138, -32.62532, -32.66875, 
        -32.71188, -32.75499, -32.7975, -32.84164, -32.88662, -32.93259, 
        -32.97953, -33.02731, -33.0756, -33.12409, -33.17254, -33.22072, 
        -33.26836, -33.31526, -33.36132, -33.40662, -33.45147, -33.49524, 
        -33.5401, -33.585, -33.62966, -33.67387, -33.71751, -33.76061, 
        -33.80331, -33.84576, -33.88808, -33.93033, -33.97248, -34.01446, 
        -34.05628, -34.09812, -34.13933, -34.1823, -34.22623, -34.27132, 
        -34.31738, -34.36451, -34.41278, -34.46212, -34.51226, -34.56279, 
        -34.6134, -34.66405, -34.71498, -34.76649, -34.81889, -34.8724, 
        -34.92712, -34.98185, -35.0384, -35.09539, -35.15255, -35.20976, 
        -35.26698, -35.32404, -35.38039, -35.43545, -35.48893, -35.541, 
        -35.59214, -35.64269, -35.69275, -35.7421, -35.7908, -35.83921, 
        -35.88666, -35.93531, -35.98392, -36.03221, -36.07993, -36.12691, 
        -36.17288, -36.21739, -36.26016, -36.3012, -36.34089, -36.37974, 
        -36.41816, -36.45623, -36.49386, -36.53095, -36.56734, -36.60274, 
        -36.63556, -36.66718, -36.69622, -36.72277, -36.74736, -36.77071, 
        -36.79363, -36.81657, -36.8397, -36.86297, -36.88614, -36.90901, 
        -36.93155, -36.95394, -36.9762, -36.99851, -37.02056, -37.04208, 
        -37.06295, -37.08333, -37.10262, -37.12325, -37.14446, -37.1662, 
        -37.18827, -37.21048, -37.23287, -37.25574, -37.27944, -37.30417, 
        -37.32974, -37.35585, -37.38228, -37.40891, -37.43567, -37.46239, 
        -37.48897, -37.51535, -37.54152, -37.56771, -37.59424, -37.62041, 
        -37.64819, -37.6762, -37.70398, -37.73128, -37.75808, -37.78471, 
        -37.81114, -37.83743, -37.86356, -37.88945, -37.91499, -37.94007, 
        -37.96448, -37.98815, -38.01115, -38.03378, -38.0567, -38.08061, 
        -38.10625, -38.13371, -38.16278, -38.19176, -38.22152, -38.24992, 
        -38.27631, -38.30083, -38.32434, -38.34795, -38.37267, -38.39897, 
        -38.42691, -38.45625, -38.48639, -38.51661, -38.54642, -38.57555, 
        -38.60395, -38.63149, -38.65845, -38.68508, -38.71195, -38.73926, 
        -38.76689, -38.79445, -38.82134, -38.84703, -38.87022, -38.89284, 
        -38.91389, -38.93364, -38.95206, -38.96917, -38.98508, -39.0001, 
        -39.01463, -39.0289, -39.04277, -39.05625, -39.06938, -39.08235, 
        -39.09549, -39.10902, -39.12307, -39.13748, -39.15177, -39.16534, 
        -39.17752, -39.18788, -39.19628, -39.20302, -39.20865, -39.21397, 
        -39.22002, -39.22793, -39.23755, -39.25147, -39.26898, -39.29019, 
        -39.3152, -39.34373, -39.3754, -39.40968, -39.44584, -39.48307, 
        -39.52052, -39.55745, -39.59338, -39.62815, -39.66182, -39.69423, 
        -39.72522, -39.75473, -39.78298, -39.8103, -39.83701, -39.86333, 
        -39.88919, -39.91446, -39.93892, -39.96226, -39.98413, -40.00405, 
        -40.02168, -40.03704, -40.05072, -40.06332, -40.07546, -40.08755, 
        -40.09857, -40.1105, -40.12246, -40.13454, -40.14645, -40.15763, 
        -40.16756, -40.17585, -40.18248, -40.18778, -40.19218, -40.19607, 
        -40.19958, -40.20266, -40.20521, -40.20724, -40.20889, -40.21041, 
        -40.21196, -40.21339, -40.21413, -40.21353, -40.21108, -40.2065, 
        -40.19965, -40.19042, -40.17886, -40.16543, -40.151, -40.13671, 
        -40.12282, -40.10883, -40.09355, -40.07577, -40.05489, -40.03098, 
        -40.00428, -39.97482, -39.94222, -39.90603, -39.86589, -39.82161, 
        -39.7729, -39.7183, -39.65918, -39.59399, -39.52234, -39.44452, 
        -39.36173,
  -31.83461, -31.8791, -31.92387, -31.96771, -32.01107, -32.05443, 
        -32.09789, -32.14183, -32.18613, -32.23055, -32.27486, -32.31923, 
        -32.36377, -32.40849, -32.45343, -32.49726, -32.54155, -32.58531, 
        -32.62875, -32.67219, -32.716, -32.76009, -32.80483, -32.85056, 
        -32.89724, -32.94485, -32.99314, -33.0416, -33.09001, -33.13804, 
        -33.1842, -33.2306, -33.2762, -33.32118, -33.36589, -33.41059, 
        -33.45539, -33.5001, -33.54443, -33.5885, -33.63224, -33.67551, 
        -33.71848, -33.76108, -33.80356, -33.84488, -33.88707, -33.92933, 
        -33.97165, -34.01434, -34.05754, -34.10141, -34.14619, -34.19192, 
        -34.23868, -34.28648, -34.33537, -34.3852, -34.43565, -34.48638, 
        -34.53714, -34.58796, -34.63821, -34.69025, -34.74333, -34.79776, 
        -34.85352, -34.91052, -34.96825, -35.02626, -35.08427, -35.14207, 
        -35.19906, -35.25549, -35.31105, -35.36496, -35.41764, -35.46943, 
        -35.51967, -35.57056, -35.62148, -35.67134, -35.72044, -35.76954, 
        -35.8177, -35.86611, -35.91433, -35.96227, -36.00933, -36.05589, 
        -36.1018, -36.14668, -36.19013, -36.23196, -36.27238, -36.31178, 
        -36.34954, -36.38786, -36.42527, -36.46218, -36.49797, -36.53282, 
        -36.56627, -36.59753, -36.62651, -36.65306, -36.67781, -36.70167, 
        -36.72513, -36.74865, -36.77235, -36.79618, -36.81982, -36.84324, 
        -36.86625, -36.8879, -36.91056, -36.93314, -36.95546, -36.97725, 
        -36.99854, -37.01939, -37.04019, -37.06134, -37.08312, -37.1055, 
        -37.1284, -37.15164, -37.17503, -37.19883, -37.2233, -37.24859, 
        -37.27456, -37.30089, -37.32731, -37.35377, -37.37907, -37.40508, 
        -37.43085, -37.45662, -37.48255, -37.50898, -37.53612, -37.564, 
        -37.59244, -37.62107, -37.64948, -37.67744, -37.70493, -37.73209, 
        -37.75888, -37.78529, -37.81144, -37.83723, -37.86282, -37.88792, 
        -37.91222, -37.93584, -37.95831, -37.98139, -38.00492, -38.02958, 
        -38.05587, -38.08393, -38.11351, -38.14384, -38.1739, -38.20251, 
        -38.22929, -38.25447, -38.27888, -38.30341, -38.32883, -38.35526, 
        -38.38287, -38.41138, -38.44043, -38.46967, -38.49878, -38.52743, 
        -38.55552, -38.58289, -38.60868, -38.63512, -38.66156, -38.68832, 
        -38.71518, -38.7419, -38.76775, -38.79244, -38.81606, -38.83801, 
        -38.85876, -38.87828, -38.89649, -38.91341, -38.92901, -38.94359, 
        -38.95766, -38.97141, -38.98485, -38.99798, -39.01097, -39.02414, 
        -39.038, -39.05225, -39.06747, -39.08349, -39.09918, -39.11342, 
        -39.12745, -39.14, -39.15041, -39.15922, -39.16685, -39.17404, 
        -39.18183, -39.19138, -39.20354, -39.2188, -39.2373, -39.25924, 
        -39.28465, -39.31326, -39.34467, -39.37862, -39.41412, -39.45041, 
        -39.48693, -39.5231, -39.55855, -39.59321, -39.62674, -39.65902, 
        -39.68985, -39.71923, -39.74742, -39.77472, -39.80132, -39.8273, 
        -39.85139, -39.87547, -39.89888, -39.92107, -39.94223, -39.96194, 
        -39.97996, -39.9961, -40.01064, -40.02407, -40.03683, -40.04922, 
        -40.06126, -40.07307, -40.08475, -40.0966, -40.10833, -40.11945, 
        -40.12941, -40.13771, -40.14426, -40.14942, -40.1534, -40.15679, 
        -40.15968, -40.16212, -40.16406, -40.16557, -40.1669, -40.1683, 
        -40.16993, -40.17166, -40.17224, -40.1715, -40.16882, -40.16374, 
        -40.15642, -40.14674, -40.13479, -40.12025, -40.10588, -40.09168, 
        -40.07786, -40.064, -40.04853, -40.03027, -40.00866, -39.98386, 
        -39.95623, -39.92587, -39.89247, -39.85558, -39.81484, -39.77015, 
        -39.72114, -39.66725, -39.60806, -39.54253, -39.47036, -39.39192, 
        -39.30868,
  -31.74743, -31.7936, -31.83904, -31.88368, -31.9276, -31.97112, 
        -32.01455, -32.05834, -32.10243, -32.14685, -32.19043, -32.23515, 
        -32.28007, -32.32519, -32.37043, -32.41558, -32.46013, -32.50426, 
        -32.54808, -32.59177, -32.63556, -32.67963, -32.72425, -32.76973, 
        -32.81623, -32.86275, -32.91101, -32.95958, -33.008, -33.05582, 
        -33.10278, -33.14888, -33.19429, -33.23924, -33.28397, -33.32857, 
        -33.37299, -33.41711, -33.46089, -33.50451, -33.54718, -33.59065, 
        -33.63406, -33.67717, -33.71994, -33.76246, -33.80492, -33.84754, 
        -33.89043, -33.93381, -33.97785, -34.02264, -34.06825, -34.11474, 
        -34.16218, -34.21068, -34.25919, -34.30946, -34.36015, -34.41095, 
        -34.46177, -34.5128, -34.56441, -34.61688, -34.6707, -34.72606, 
        -34.78291, -34.84094, -34.89966, -34.95853, -35.01707, -35.07484, 
        -35.13198, -35.18689, -35.24152, -35.29479, -35.34702, -35.39862, 
        -35.44991, -35.50136, -35.55247, -35.60298, -35.65271, -35.70172, 
        -35.75011, -35.79803, -35.84544, -35.89233, -35.93871, -35.98488, 
        -36.02972, -36.07496, -36.11906, -36.16182, -36.20314, -36.24337, 
        -36.28263, -36.32103, -36.35847, -36.39489, -36.43017, -36.46424, 
        -36.49688, -36.52777, -36.55679, -36.58375, -36.60912, -36.63374, 
        -36.65812, -36.68146, -36.70597, -36.73052, -36.75488, -36.7788, 
        -36.80217, -36.82524, -36.84797, -36.87048, -36.89281, -36.91468, 
        -36.93633, -36.95779, -36.97927, -37.00111, -37.02361, -37.04686, 
        -37.07074, -37.09498, -37.11938, -37.14302, -37.16816, -37.19386, 
        -37.22015, -37.24674, -37.2734, -37.29974, -37.32578, -37.35121, 
        -37.37628, -37.40134, -37.42685, -37.45328, -37.48073, -37.5091, 
        -37.53806, -37.5672, -37.59618, -37.62483, -37.65294, -37.68053, 
        -37.70652, -37.73298, -37.75895, -37.78466, -37.81003, -37.83491, 
        -37.8592, -37.88311, -37.90659, -37.93043, -37.95503, -37.98088, 
        -38.00811, -38.03694, -38.0669, -38.09731, -38.12713, -38.15563, 
        -38.18251, -38.20823, -38.23351, -38.25907, -38.28528, -38.31213, 
        -38.33847, -38.36615, -38.39414, -38.42241, -38.4508, -38.47894, 
        -38.50662, -38.53367, -38.5602, -38.58644, -38.61264, -38.63887, 
        -38.66494, -38.69058, -38.71549, -38.73945, -38.76234, -38.78404, 
        -38.80452, -38.82398, -38.84203, -38.85886, -38.87435, -38.8887, 
        -38.90244, -38.91573, -38.92762, -38.94035, -38.95322, -38.96658, 
        -38.9808, -38.99603, -39.01226, -39.02918, -39.04627, -39.063, 
        -39.07883, -39.0933, -39.10606, -39.1171, -39.1268, -39.13592, 
        -39.14558, -39.15675, -39.17035, -39.18677, -39.20616, -39.22859, 
        -39.25413, -39.28274, -39.31414, -39.3477, -39.38258, -39.41805, 
        -39.45362, -39.48899, -39.52298, -39.55735, -39.59079, -39.62294, 
        -39.65357, -39.68277, -39.71087, -39.73814, -39.76461, -39.79017, 
        -39.81463, -39.83782, -39.85994, -39.88107, -39.90158, -39.92112, 
        -39.93944, -39.9563, -39.97171, -39.98588, -39.99926, -40.01197, 
        -40.02405, -40.03566, -40.04691, -40.05805, -40.06921, -40.08012, 
        -40.08998, -40.09844, -40.10524, -40.11057, -40.11457, -40.11757, 
        -40.11979, -40.12046, -40.12173, -40.12278, -40.12386, -40.12529, 
        -40.12719, -40.12881, -40.12973, -40.12878, -40.12554, -40.11991, 
        -40.11195, -40.10176, -40.08954, -40.07584, -40.06149, -40.04732, 
        -40.03345, -40.01915, -40.00308, -39.98406, -39.96159, -39.93585, 
        -39.90714, -39.87569, -39.84129, -39.80357, -39.76222, -39.71696, 
        -39.66752, -39.61337, -39.55375, -39.48781, -39.41522, -39.33671, 
        -39.25365,
  -31.66302, -31.70973, -31.75566, -31.80071, -31.8449, -31.8885, 
        -31.93096, -31.97466, -32.01881, -32.06341, -32.10836, -32.15356, 
        -32.19899, -32.24458, -32.29018, -32.33552, -32.38036, -32.42465, 
        -32.46852, -32.51221, -32.55492, -32.59888, -32.64342, -32.68883, 
        -32.73532, -32.78284, -32.83112, -32.8797, -32.92809, -32.97586, 
        -33.02278, -33.06892, -33.11447, -33.15963, -33.2045, -33.24805, 
        -33.29215, -33.33572, -33.37887, -33.42192, -33.46517, -33.50871, 
        -33.55238, -33.59595, -33.63914, -33.68214, -33.72511, -33.76823, 
        -33.8117, -33.85573, -33.90047, -33.945, -33.99136, -34.03858, 
        -34.08676, -34.13597, -34.18609, -34.23686, -34.28791, -34.33897, 
        -34.39, -34.44126, -34.49314, -34.54606, -34.60043, -34.65644, 
        -34.71402, -34.77177, -34.83113, -34.8905, -34.94934, -35.00727, 
        -35.06407, -35.11955, -35.17364, -35.22646, -35.27841, -35.32995, 
        -35.38145, -35.43305, -35.48449, -35.53539, -35.58546, -35.6346, 
        -35.68287, -35.72931, -35.77602, -35.82211, -35.86789, -35.91365, 
        -35.9594, -36.00488, -36.04956, -36.09305, -36.13519, -36.17603, 
        -36.21568, -36.25418, -36.29147, -36.32751, -36.36229, -36.39585, 
        -36.42812, -36.45792, -36.48709, -36.51467, -36.54092, -36.56656, 
        -36.59186, -36.61715, -36.64249, -36.66782, -36.69286, -36.71734, 
        -36.74113, -36.7643, -36.78699, -36.80938, -36.83158, -36.85366, 
        -36.87569, -36.89775, -36.91901, -36.9417, -36.96508, -36.98927, 
        -37.01413, -37.03936, -37.06467, -37.0901, -37.11583, -37.14202, 
        -37.16865, -37.19545, -37.22216, -37.24852, -37.27433, -37.29944, 
        -37.32402, -37.34854, -37.3736, -37.3997, -37.42706, -37.45464, 
        -37.48389, -37.51353, -37.54307, -37.57221, -37.60069, -37.62859, 
        -37.65561, -37.6819, -37.7077, -37.73318, -37.75833, -37.78305, 
        -37.80739, -37.83151, -37.8556, -37.88042, -37.90631, -37.93325, 
        -37.96144, -37.99084, -38.021, -38.05125, -38.07978, -38.10806, 
        -38.13503, -38.16116, -38.18711, -38.21346, -38.24029, -38.26751, 
        -38.29477, -38.322, -38.34932, -38.37683, -38.40449, -38.43202, 
        -38.45916, -38.48573, -38.51186, -38.53773, -38.5635, -38.58915, 
        -38.61449, -38.63931, -38.66344, -38.68677, -38.70925, -38.72966, 
        -38.7501, -38.76946, -38.7876, -38.80444, -38.81999, -38.83439, 
        -38.84789, -38.86074, -38.8732, -38.88554, -38.89819, -38.91155, 
        -38.92602, -38.94175, -38.95865, -38.97643, -38.99463, -39.01271, 
        -39.03019, -39.04667, -39.06163, -39.07495, -39.08687, -39.09812, 
        -39.10969, -39.12262, -39.13769, -39.15427, -39.17448, -39.19746, 
        -39.22326, -39.25191, -39.28315, -39.31629, -39.35051, -39.38514, 
        -39.4197, -39.45418, -39.48846, -39.52235, -39.55551, -39.58752, 
        -39.61808, -39.64727, -39.67526, -39.70242, -39.72869, -39.75383, 
        -39.7776, -39.79998, -39.82132, -39.84167, -39.86159, -39.881, 
        -39.89963, -39.91708, -39.93322, -39.94814, -39.96204, -39.97501, 
        -39.98722, -39.9975, -40.00808, -40.01833, -40.02868, -40.0389, 
        -40.04853, -40.05704, -40.06407, -40.06957, -40.07361, -40.07637, 
        -40.0781, -40.07915, -40.07985, -40.08051, -40.08141, -40.08288, 
        -40.08482, -40.08664, -40.08744, -40.0863, -40.08269, -40.07659, 
        -40.06819, -40.05764, -40.04515, -40.03124, -40.01665, -40.00211, 
        -39.98764, -39.97264, -39.95573, -39.93581, -39.91239, -39.88563, 
        -39.8559, -39.82343, -39.7881, -39.74962, -39.7076, -39.66175, 
        -39.6117, -39.55692, -39.49562, -39.42912, -39.35631, -39.27805, 
        -39.19635,
  -31.58008, -31.62618, -31.67245, -31.7177, -31.76197, -31.80557, 
        -31.84902, -31.89276, -31.9371, -31.98199, -32.02736, -32.07308, 
        -32.11904, -32.16509, -32.21102, -32.25558, -32.30053, -32.34486, 
        -32.3887, -32.43228, -32.47586, -32.51974, -32.56427, -32.60972, 
        -32.65626, -32.70383, -32.75212, -32.80056, -32.849, -32.89672, 
        -32.94268, -32.98901, -33.03494, -33.08056, -33.12579, -33.17043, 
        -33.21429, -33.25736, -33.29986, -33.3423, -33.38517, -33.42862, 
        -33.47264, -33.5167, -33.56057, -33.6042, -33.64675, -33.6904, 
        -33.73438, -33.77891, -33.82418, -33.87032, -33.91736, -33.96534, 
        -34.01435, -34.06436, -34.11521, -34.16656, -34.21804, -34.26945, 
        -34.3208, -34.37236, -34.42353, -34.47676, -34.53143, -34.58785, 
        -34.64582, -34.70496, -34.76467, -34.82431, -34.88331, -34.94124, 
        -34.99785, -35.053, -35.10673, -35.15927, -35.21117, -35.26273, 
        -35.31432, -35.36502, -35.41665, -35.46783, -35.51823, -35.56759, 
        -35.61578, -35.66279, -35.70878, -35.75413, -35.7993, -35.84466, 
        -35.8903, -35.93592, -35.98102, -36.02515, -36.06799, -36.10944, 
        -36.14944, -36.18697, -36.22404, -36.25971, -36.29408, -36.32724, 
        -36.35933, -36.3902, -36.41982, -36.44818, -36.47548, -36.50204, 
        -36.52823, -36.5543, -36.58039, -36.60646, -36.63222, -36.6573, 
        -36.68144, -36.70469, -36.72626, -36.74843, -36.77049, -36.79269, 
        -36.81517, -36.83798, -36.86117, -36.88486, -36.90921, -36.93433, 
        -36.96009, -36.98618, -37.01233, -37.03844, -37.06469, -37.09123, 
        -37.11809, -37.14504, -37.17184, -37.19826, -37.22307, -37.24813, 
        -37.27254, -37.29678, -37.32148, -37.34718, -37.37421, -37.40256, 
        -37.43192, -37.46178, -37.49161, -37.52097, -37.54958, -37.57743, 
        -37.60432, -37.63046, -37.65606, -37.68142, -37.70639, -37.73094, 
        -37.75535, -37.77983, -37.80385, -37.8298, -37.85686, -37.88501, 
        -37.91416, -37.94409, -37.97433, -38.00428, -38.03334, -38.06124, 
        -38.08818, -38.11465, -38.14116, -38.16833, -38.19584, -38.22341, 
        -38.25072, -38.2777, -38.30455, -38.3315, -38.35854, -38.38543, 
        -38.41191, -38.43792, -38.46356, -38.48802, -38.51338, -38.53853, 
        -38.56326, -38.58739, -38.6109, -38.63378, -38.65594, -38.67727, 
        -38.69766, -38.71701, -38.73524, -38.75224, -38.76798, -38.78255, 
        -38.79598, -38.80858, -38.82066, -38.83265, -38.84506, -38.85836, 
        -38.87291, -38.88889, -38.90618, -38.92451, -38.9435, -38.96269, 
        -38.98056, -38.99895, -39.01603, -39.03157, -39.04573, -39.05912, 
        -39.07266, -39.08733, -39.10386, -39.12257, -39.14365, -39.16719, 
        -39.19334, -39.22216, -39.25333, -39.28612, -39.3197, -39.35345, 
        -39.38707, -39.4206, -39.45407, -39.48736, -39.52013, -39.55191, 
        -39.58234, -39.6114, -39.6393, -39.66631, -39.69239, -39.71728, 
        -39.74069, -39.76163, -39.78235, -39.80228, -39.8218, -39.84104, 
        -39.85979, -39.87767, -39.89436, -39.90978, -39.92408, -39.93726, 
        -39.94926, -39.96004, -39.96983, -39.97912, -39.98844, -39.99789, 
        -40.00713, -40.01567, -40.023, -40.02884, -40.03302, -40.03561, 
        -40.03689, -40.03733, -40.03746, -40.03774, -40.03851, -40.03998, 
        -40.042, -40.0439, -40.04462, -40.04325, -40.03926, -40.03267, 
        -40.02375, -40.01276, -39.99997, -39.98574, -39.97061, -39.95435, 
        -39.93885, -39.92266, -39.90465, -39.88376, -39.85947, -39.8318, 
        -39.80114, -39.76759, -39.73134, -39.69225, -39.64959, -39.60306, 
        -39.5522, -39.49646, -39.43515, -39.3678, -39.29486, -39.21738, 
        -39.13761,
  -31.49746, -31.54485, -31.5913, -31.63661, -31.68083, -31.72438, 
        -31.76788, -31.81176, -31.85625, -31.90144, -31.94723, -31.99251, 
        -32.03905, -32.08556, -32.13179, -32.17743, -32.22231, -32.26649, 
        -32.31017, -32.35358, -32.39712, -32.44108, -32.48577, -32.53139, 
        -32.57808, -32.62469, -32.67303, -32.72146, -32.76956, -32.81725, 
        -32.86404, -32.91055, -32.95691, -33.00314, -33.04877, -33.09364, 
        -33.13746, -33.18034, -33.2226, -33.26474, -33.30741, -33.34986, 
        -33.39406, -33.43858, -33.48309, -33.52745, -33.57165, -33.61592, 
        -33.66042, -33.70538, -33.75107, -33.79766, -33.84534, -33.89413, 
        -33.944, -33.99487, -34.04644, -34.09739, -34.1494, -34.20131, 
        -34.25313, -34.3051, -34.35756, -34.41094, -34.46575, -34.5221, 
        -34.58005, -34.63928, -34.69889, -34.75862, -34.81781, -34.8757, 
        -34.93228, -34.98613, -35.0396, -35.09214, -35.14399, -35.19555, 
        -35.24714, -35.29883, -35.35048, -35.40179, -35.45233, -35.50203, 
        -35.55025, -35.597, -35.64247, -35.68735, -35.73207, -35.77718, 
        -35.82277, -35.86747, -35.91282, -35.95737, -36.00071, -36.04254, 
        -36.08274, -36.12111, -36.15802, -36.19331, -36.22754, -36.26065, 
        -36.2928, -36.32407, -36.35439, -36.38365, -36.41186, -36.43916, 
        -36.46604, -36.49254, -36.51809, -36.5447, -36.57112, -36.5968, 
        -36.62138, -36.64482, -36.6675, -36.68964, -36.7117, -36.73419, 
        -36.75717, -36.78078, -36.80498, -36.82965, -36.85495, -36.8808, 
        -36.90726, -36.93395, -36.96074, -36.98753, -37.01322, -37.0401, 
        -37.0672, -37.09423, -37.12116, -37.14754, -37.1734, -37.19863, 
        -37.22317, -37.24754, -37.27206, -37.29739, -37.32387, -37.35189, 
        -37.38113, -37.41092, -37.44075, -37.47005, -37.49849, -37.52612, 
        -37.55278, -37.57793, -37.60343, -37.62875, -37.65366, -37.67831, 
        -37.70286, -37.72781, -37.75366, -37.78067, -37.8089, -37.83802, 
        -37.86787, -37.89813, -37.92821, -37.95779, -37.98643, -38.01406, 
        -38.04104, -38.06797, -38.09507, -38.12273, -38.1507, -38.17852, 
        -38.20494, -38.23182, -38.25834, -38.28487, -38.31142, -38.33766, 
        -38.36344, -38.38883, -38.41396, -38.43887, -38.46376, -38.48851, 
        -38.51271, -38.53623, -38.55929, -38.58183, -38.60382, -38.62513, 
        -38.64554, -38.66491, -38.68325, -38.70044, -38.71648, -38.7313, 
        -38.74488, -38.75742, -38.76929, -38.7801, -38.79232, -38.8055, 
        -38.81995, -38.83593, -38.85328, -38.87192, -38.89153, -38.91162, 
        -38.93181, -38.95191, -38.97104, -38.98866, -39.00511, -39.02063, 
        -39.03619, -39.0526, -39.0705, -39.09052, -39.1125, -39.13673, 
        -39.16333, -39.19248, -39.22355, -39.25591, -39.2888, -39.32169, 
        -39.35438, -39.38698, -39.41859, -39.45116, -39.48339, -39.51482, 
        -39.54506, -39.57399, -39.60174, -39.62848, -39.65442, -39.6792, 
        -39.7025, -39.72438, -39.74494, -39.76459, -39.78379, -39.80281, 
        -39.82158, -39.83978, -39.85688, -39.8727, -39.88717, -39.90019, 
        -39.91163, -39.92169, -39.93066, -39.93913, -39.94767, -39.95645, 
        -39.9653, -39.97369, -39.98117, -39.98715, -39.9914, -39.99398, 
        -39.995, -39.9949, -39.99442, -39.99331, -39.99383, -39.99512, 
        -39.99711, -39.99896, -39.99966, -39.9982, -39.99404, -39.98708, 
        -39.9777, -39.96623, -39.953, -39.93819, -39.92222, -39.90575, 
        -39.88891, -39.87122, -39.85197, -39.83015, -39.80509, -39.77663, 
        -39.74516, -39.7109, -39.67381, -39.63406, -39.59078, -39.5435, 
        -39.49158, -39.43472, -39.37208, -39.30375, -39.23064, -39.15432, 
        -39.07724,
  -31.41645, -31.46424, -31.51095, -31.55639, -31.6007, -31.64433, 
        -31.68689, -31.73085, -31.77548, -31.82093, -31.86713, -31.91391, 
        -31.96093, -32.00789, -32.05422, -32.09975, -32.14437, -32.18826, 
        -32.23167, -32.27507, -32.31867, -32.36196, -32.40707, -32.45309, 
        -32.49999, -32.54776, -32.59604, -32.6444, -32.69242, -32.73984, 
        -32.78668, -32.83315, -32.87967, -32.92604, -32.97195, -33.01694, 
        -33.05994, -33.10301, -33.1454, -33.18774, -33.23058, -33.27415, 
        -33.31858, -33.3635, -33.4085, -33.45345, -33.49836, -33.54332, 
        -33.58849, -33.63393, -33.68009, -33.72628, -33.77452, -33.82404, 
        -33.87472, -33.92625, -33.97849, -34.03107, -34.08368, -34.1362, 
        -34.18857, -34.241, -34.29377, -34.3473, -34.4021, -34.45844, 
        -34.51631, -34.5752, -34.63379, -34.69357, -34.75256, -34.81018, 
        -34.86675, -34.92149, -34.97497, -35.02727, -35.0791, -35.13056, 
        -35.18203, -35.23373, -35.28517, -35.33648, -35.38694, -35.43663, 
        -35.48478, -35.53036, -35.57564, -35.62027, -35.66492, -35.71006, 
        -35.75574, -35.80149, -35.84699, -35.89172, -35.93532, -35.97736, 
        -36.01758, -36.05581, -36.09249, -36.12756, -36.16175, -36.19493, 
        -36.2276, -36.25946, -36.28949, -36.3196, -36.3485, -36.37644, 
        -36.40372, -36.43045, -36.45722, -36.48418, -36.51107, -36.53731, 
        -36.56247, -36.58646, -36.60955, -36.63201, -36.65446, -36.67738, 
        -36.70095, -36.7254, -36.75038, -36.77502, -36.80094, -36.82747, 
        -36.85442, -36.88174, -36.9091, -36.9364, -36.96358, -36.99082, 
        -37.01798, -37.04505, -37.07186, -37.09826, -37.12431, -37.14965, 
        -37.17434, -37.19862, -37.22297, -37.24814, -37.27445, -37.30221, 
        -37.33018, -37.35993, -37.38965, -37.41879, -37.44712, -37.47455, 
        -37.50112, -37.52712, -37.55273, -37.57809, -37.60312, -37.62794, 
        -37.65285, -37.67838, -37.70504, -37.73285, -37.76177, -37.79153, 
        -37.82171, -37.85204, -37.88205, -37.91154, -37.94, -37.96668, 
        -37.99381, -38.02085, -38.04819, -38.07597, -38.10398, -38.13187, 
        -38.1592, -38.18591, -38.21218, -38.23826, -38.26417, -38.28984, 
        -38.31511, -38.33997, -38.36463, -38.38917, -38.41377, -38.43801, 
        -38.46175, -38.48532, -38.50812, -38.53028, -38.55194, -38.57325, 
        -38.59271, -38.61201, -38.6302, -38.64749, -38.66372, -38.67882, 
        -38.69257, -38.70517, -38.71706, -38.72885, -38.74105, -38.75414, 
        -38.7685, -38.78434, -38.80182, -38.82062, -38.84087, -38.86178, 
        -38.88332, -38.9049, -38.92594, -38.94553, -38.96401, -38.98159, 
        -38.999, -39.01722, -39.03643, -39.05759, -39.07953, -39.10452, 
        -39.1316, -39.16104, -39.19199, -39.22392, -39.25619, -39.28832, 
        -39.32018, -39.35189, -39.38371, -39.41555, -39.44715, -39.47813, 
        -39.5081, -39.53685, -39.56445, -39.59106, -39.61671, -39.64149, 
        -39.66484, -39.68663, -39.70721, -39.72675, -39.74577, -39.76474, 
        -39.7837, -39.80211, -39.81951, -39.83548, -39.84977, -39.86224, 
        -39.87294, -39.88207, -39.88935, -39.89719, -39.9052, -39.91357, 
        -39.92213, -39.93023, -39.93744, -39.94344, -39.94773, -39.95015, 
        -39.95092, -39.95049, -39.94965, -39.94913, -39.94934, -39.9505, 
        -39.95222, -39.9542, -39.95481, -39.9534, -39.94907, -39.94185, 
        -39.93206, -39.92013, -39.90598, -39.89017, -39.87296, -39.85512, 
        -39.83667, -39.8176, -39.79715, -39.77439, -39.74866, -39.7197, 
        -39.68761, -39.65275, -39.61517, -39.57457, -39.53058, -39.48235, 
        -39.42911, -39.3707, -39.30664, -39.23746, -39.16335, -39.0886, 
        -39.01445,
  -31.33638, -31.38442, -31.43037, -31.47602, -31.52064, -31.56452, 
        -31.60822, -31.65224, -31.69695, -31.74257, -31.78909, -31.83628, 
        -31.88373, -31.93086, -31.97716, -32.02237, -32.06555, -32.10904, 
        -32.1523, -32.19574, -32.23976, -32.28458, -32.33028, -32.3768, 
        -32.42406, -32.4719, -32.52008, -32.56822, -32.61596, -32.6631, 
        -32.70977, -32.75525, -32.80172, -32.84806, -32.89396, -32.9391, 
        -32.98335, -33.02676, -33.06975, -33.11265, -33.15599, -33.20005, 
        -33.24486, -33.29018, -33.33571, -33.38129, -33.42589, -33.47156, 
        -33.5174, -33.56357, -33.61037, -33.65813, -33.70707, -33.75727, 
        -33.80859, -33.86065, -33.91336, -33.9664, -34.01959, -34.07269, 
        -34.12567, -34.17859, -34.2317, -34.28444, -34.33928, -34.3955, 
        -34.45309, -34.51176, -34.57109, -34.63051, -34.68927, -34.74712, 
        -34.80342, -34.85812, -34.91142, -34.96371, -35.01543, -35.06691, 
        -35.11832, -35.16968, -35.21983, -35.2706, -35.32071, -35.36987, 
        -35.41777, -35.46424, -35.50952, -35.55437, -35.59931, -35.64473, 
        -35.69059, -35.73652, -35.78209, -35.82689, -35.87046, -35.91259, 
        -35.95282, -35.99112, -36.02663, -36.06174, -36.09591, -36.12946, 
        -36.16251, -36.19496, -36.22665, -36.25735, -36.28685, -36.31513, 
        -36.34245, -36.36929, -36.39618, -36.42334, -36.45061, -36.47746, 
        -36.5034, -36.52822, -36.55206, -36.57428, -36.5974, -36.62095, 
        -36.6453, -36.67063, -36.69639, -36.72267, -36.74928, -36.77622, 
        -36.80352, -36.83112, -36.8589, -36.88667, -36.91432, -36.9418, 
        -36.96904, -36.99603, -37.02275, -37.04918, -37.07523, -37.0998, 
        -37.12473, -37.14921, -37.17367, -37.19875, -37.22492, -37.25248, 
        -37.28128, -37.31079, -37.34034, -37.36938, -37.39763, -37.42503, 
        -37.45172, -37.47792, -37.50375, -37.52929, -37.55458, -37.57972, 
        -37.60506, -37.63113, -37.65829, -37.68565, -37.71498, -37.74493, 
        -37.7751, -37.80524, -37.83509, -37.86442, -37.89301, -37.92087, 
        -37.94825, -37.97547, -38.00285, -38.03045, -38.05814, -38.08564, 
        -38.1126, -38.13899, -38.16488, -38.19044, -38.21577, -38.24081, 
        -38.2655, -38.28989, -38.31414, -38.33739, -38.36166, -38.38576, 
        -38.40949, -38.43266, -38.45539, -38.47754, -38.49917, -38.52018, 
        -38.54034, -38.55952, -38.57773, -38.59503, -38.61134, -38.62647, 
        -38.64034, -38.65308, -38.66514, -38.67707, -38.68941, -38.70258, 
        -38.71695, -38.73279, -38.7502, -38.76945, -38.79014, -38.81194, 
        -38.83486, -38.8569, -38.87946, -38.90099, -38.92134, -38.94077, 
        -38.95996, -38.97963, -39.00034, -39.0225, -39.04647, -39.07211, 
        -39.09985, -39.12942, -39.1603, -39.1919, -39.22364, -39.25519, 
        -39.28644, -39.31754, -39.34863, -39.37973, -39.41066, -39.44109, 
        -39.47064, -39.49914, -39.5265, -39.55288, -39.57839, -39.60294, 
        -39.6263, -39.64828, -39.6679, -39.68749, -39.7065, -39.72553, 
        -39.74445, -39.76297, -39.78047, -39.79633, -39.81015, -39.82183, 
        -39.83158, -39.83989, -39.84748, -39.85497, -39.86281, -39.87111, 
        -39.87929, -39.88717, -39.89425, -39.90011, -39.90434, -39.90662, 
        -39.90717, -39.9065, -39.90538, -39.90449, -39.90434, -39.90515, 
        -39.90663, -39.90846, -39.90913, -39.90767, -39.90327, -39.89585, 
        -39.88558, -39.87276, -39.85766, -39.84061, -39.82206, -39.80259, 
        -39.78162, -39.76107, -39.73949, -39.71598, -39.68972, -39.66031, 
        -39.62779, -39.59237, -39.55423, -39.51296, -39.46798, -39.4185, 
        -39.3639, -39.30383, -39.23832, -39.16817, -39.09542, -39.02225, 
        -38.95133,
  -31.25661, -31.30474, -31.35184, -31.39783, -31.44279, -31.48701, 
        -31.53091, -31.57499, -31.61975, -31.66551, -31.71231, -31.75884, 
        -31.80651, -31.85362, -31.89968, -31.94441, -31.9881, -32.03123, 
        -32.07444, -32.11803, -32.16268, -32.20825, -32.25474, -32.30178, 
        -32.34946, -32.3971, -32.44413, -32.49186, -32.5393, -32.58614, 
        -32.6326, -32.67897, -32.7253, -32.77134, -32.81708, -32.86222, 
        -32.90676, -32.95079, -32.99453, -33.03823, -33.08235, -33.12617, 
        -33.17154, -33.21745, -33.26363, -33.30979, -33.35606, -33.40245, 
        -33.44911, -33.49615, -33.54383, -33.59236, -33.64193, -33.69275, 
        -33.74447, -33.79695, -33.84995, -33.90234, -33.95591, -34.00944, 
        -34.063, -34.11644, -34.16997, -34.22394, -34.27884, -34.33501, 
        -34.39238, -34.45065, -34.50946, -34.56852, -34.62714, -34.68483, 
        -34.74107, -34.79568, -34.84789, -34.9002, -34.95198, -35.00349, 
        -35.05477, -35.10579, -35.15637, -35.20627, -35.25552, -35.30367, 
        -35.3513, -35.3976, -35.44303, -35.48824, -35.53368, -35.57951, 
        -35.62565, -35.67173, -35.71635, -35.76117, -35.80484, -35.847, 
        -35.88723, -35.92585, -35.96254, -35.9978, -36.03209, -36.06598, 
        -36.09939, -36.13226, -36.16435, -36.19537, -36.2251, -36.2535, 
        -36.28085, -36.30771, -36.33365, -36.36096, -36.38865, -36.41626, 
        -36.44311, -36.46898, -36.49385, -36.51814, -36.54232, -36.56661, 
        -36.59181, -36.61788, -36.64463, -36.67154, -36.69867, -36.72598, 
        -36.7534, -36.78115, -36.80922, -36.83736, -36.86442, -36.89206, 
        -36.91933, -36.94625, -36.97282, -36.99923, -37.02542, -37.05123, 
        -37.07652, -37.10135, -37.12607, -37.15128, -37.17747, -37.20491, 
        -37.23349, -37.26275, -37.29206, -37.32107, -37.3494, -37.37718, 
        -37.40419, -37.43088, -37.45597, -37.48181, -37.5076, -37.53314, 
        -37.55875, -37.58537, -37.61293, -37.64151, -37.67089, -37.70068, 
        -37.73057, -37.76033, -37.78992, -37.81918, -37.848, -37.87619, 
        -37.90403, -37.93121, -37.9585, -37.98547, -38.01231, -38.03905, 
        -38.06537, -38.09019, -38.11552, -38.14046, -38.16507, -38.1894, 
        -38.21347, -38.23736, -38.26128, -38.28525, -38.30933, -38.33332, 
        -38.35715, -38.38045, -38.40312, -38.42521, -38.44665, -38.46736, 
        -38.4873, -38.50631, -38.52441, -38.54165, -38.55791, -38.57302, 
        -38.58692, -38.59982, -38.61207, -38.62331, -38.63594, -38.64937, 
        -38.664, -38.68, -38.69762, -38.71719, -38.7384, -38.76118, 
        -38.78535, -38.80977, -38.83374, -38.8569, -38.879, -38.9001, 
        -38.92086, -38.94192, -38.96388, -38.98713, -39.01183, -39.03825, 
        -39.06662, -39.09641, -39.12727, -39.15858, -39.18996, -39.22128, 
        -39.25225, -39.28299, -39.31361, -39.34309, -39.37331, -39.40306, 
        -39.43206, -39.46014, -39.48719, -39.51322, -39.53837, -39.5626, 
        -39.58579, -39.60787, -39.62864, -39.64842, -39.66763, -39.68665, 
        -39.70542, -39.72402, -39.7414, -39.75689, -39.77005, -39.78085, 
        -39.78965, -39.79715, -39.80421, -39.81153, -39.8193, -39.8276, 
        -39.83579, -39.84359, -39.8506, -39.85627, -39.86032, -39.86261, 
        -39.86312, -39.86226, -39.86087, -39.85959, -39.85807, -39.85849, 
        -39.8598, -39.86108, -39.86144, -39.86005, -39.85547, -39.84778, 
        -39.83693, -39.82315, -39.80687, -39.78846, -39.76843, -39.74733, 
        -39.72591, -39.70404, -39.68148, -39.65734, -39.6307, -39.60105, 
        -39.56818, -39.53232, -39.49342, -39.45116, -39.40502, -39.35407, 
        -39.29787, -39.23614, -39.16933, -39.09858, -39.02622, -38.95472, 
        -38.88694,
  -31.17971, -31.22773, -31.27486, -31.321, -31.36625, -31.41078, 
        -31.45489, -31.49807, -31.54292, -31.58886, -31.63595, -31.68368, 
        -31.73139, -31.77831, -31.82402, -31.86837, -31.91183, -31.95483, 
        -31.99806, -32.04204, -32.08716, -32.13245, -32.17947, -32.22705, 
        -32.27473, -32.3223, -32.36997, -32.41739, -32.46447, -32.51108, 
        -32.55743, -32.60342, -32.64943, -32.69535, -32.74085, -32.78605, 
        -32.82987, -32.87443, -32.91892, -32.9635, -33.00846, -33.05408, 
        -33.10037, -33.14706, -33.19392, -33.24077, -33.28771, -33.3349, 
        -33.3824, -33.43049, -33.47912, -33.52848, -33.57782, -33.62912, 
        -33.68129, -33.73411, -33.78736, -33.84098, -33.89479, -33.94869, 
        -34.00256, -34.05646, -34.11042, -34.16472, -34.21984, -34.27592, 
        -34.33295, -34.39071, -34.4491, -34.50669, -34.56493, -34.62231, 
        -34.67843, -34.73302, -34.78631, -34.83871, -34.89064, -34.9422, 
        -34.9934, -35.04422, -35.09415, -35.14313, -35.19125, -35.2385, 
        -35.28503, -35.33088, -35.37547, -35.42095, -35.46677, -35.51294, 
        -35.5593, -35.60548, -35.65113, -35.69599, -35.73986, -35.7823, 
        -35.82304, -35.86203, -35.89914, -35.93479, -35.96948, -36.00358, 
        -36.03719, -36.07021, -36.10131, -36.13236, -36.16196, -36.19038, 
        -36.21771, -36.24475, -36.27189, -36.29956, -36.32785, -36.35614, 
        -36.38391, -36.41078, -36.43678, -36.46219, -36.48746, -36.51297, 
        -36.53916, -36.56602, -36.5935, -36.62117, -36.64783, -36.67545, 
        -36.70305, -36.73092, -36.7591, -36.78745, -36.81567, -36.8435, 
        -36.87079, -36.89772, -36.92418, -36.95065, -36.97706, -37.00322, 
        -37.02887, -37.05415, -37.07935, -37.10489, -37.13113, -37.15852, 
        -37.18687, -37.21484, -37.24404, -37.27302, -37.30167, -37.33003, 
        -37.35748, -37.38485, -37.41131, -37.43742, -37.46332, -37.48936, 
        -37.51565, -37.54249, -37.57038, -37.59897, -37.62823, -37.65776, 
        -37.68729, -37.71676, -37.74612, -37.77538, -37.80436, -37.83186, 
        -37.85987, -37.88703, -37.9138, -37.93969, -37.96575, -37.99133, 
        -38.01676, -38.04179, -38.06636, -38.09047, -38.11418, -38.1377, 
        -38.16116, -38.18461, -38.20819, -38.23195, -38.25592, -38.28001, 
        -38.30404, -38.32755, -38.35029, -38.37239, -38.39355, -38.414, 
        -38.43355, -38.45137, -38.4693, -38.48635, -38.50251, -38.51759, 
        -38.53156, -38.54459, -38.55715, -38.56971, -38.58275, -38.59664, 
        -38.61165, -38.62807, -38.64615, -38.66614, -38.68818, -38.71206, 
        -38.7373, -38.76302, -38.78845, -38.81296, -38.83625, -38.85864, 
        -38.88059, -38.90284, -38.92571, -38.94984, -38.97539, -39.00161, 
        -39.03046, -39.06062, -39.09159, -39.12296, -39.15432, -39.18562, 
        -39.21668, -39.24743, -39.27781, -39.30788, -39.33741, -39.36637, 
        -39.39467, -39.42213, -39.44865, -39.47428, -39.49908, -39.52283, 
        -39.5457, -39.56755, -39.58833, -39.60831, -39.62778, -39.64706, 
        -39.66596, -39.6842, -39.70135, -39.71634, -39.72876, -39.73867, 
        -39.74661, -39.75343, -39.75993, -39.76595, -39.7738, -39.78203, 
        -39.7904, -39.79834, -39.80515, -39.81072, -39.81478, -39.81711, 
        -39.81769, -39.81684, -39.81532, -39.81384, -39.81296, -39.81305, 
        -39.81385, -39.81465, -39.81464, -39.81267, -39.80771, -39.79942, 
        -39.78775, -39.77294, -39.75549, -39.73579, -39.71441, -39.69189, 
        -39.66924, -39.64633, -39.62282, -39.59798, -39.57107, -39.54124, 
        -39.50815, -39.47179, -39.43206, -39.38863, -39.34086, -39.28819, 
        -39.2301, -39.16667, -39.09863, -39.02735, -38.95554, -38.88492, 
        -38.82056,
  -31.10466, -31.15263, -31.1987, -31.24489, -31.29023, -31.33486, 
        -31.37909, -31.42342, -31.4685, -31.51467, -31.56193, -31.60978, 
        -31.65742, -31.70416, -31.74964, -31.79387, -31.83627, -31.87939, 
        -31.92288, -31.96728, -32.01284, -32.05955, -32.10703, -32.15475, 
        -32.20239, -32.24982, -32.29707, -32.34409, -32.39085, -32.43726, 
        -32.48334, -32.52829, -32.57395, -32.61957, -32.66503, -32.71031, 
        -32.75554, -32.80063, -32.84581, -32.89121, -32.937, -32.98345, 
        -33.03059, -33.07811, -33.1257, -33.17319, -33.22087, -33.26796, 
        -33.31646, -33.36559, -33.41523, -33.46545, -33.51646, -33.56831, 
        -33.6209, -33.67408, -33.72768, -33.78149, -33.83551, -33.88959, 
        -33.9437, -33.99788, -34.05218, -34.1058, -34.16102, -34.21695, 
        -34.27369, -34.33102, -34.38892, -34.4469, -34.50457, -34.5615, 
        -34.61728, -34.67189, -34.72537, -34.77801, -34.83009, -34.88179, 
        -34.9331, -34.9836, -35.03212, -35.08039, -35.12749, -35.17341, 
        -35.21883, -35.26402, -35.30924, -35.35476, -35.40078, -35.44718, 
        -35.4936, -35.53983, -35.58545, -35.63049, -35.67457, -35.71743, 
        -35.75875, -35.79832, -35.83514, -35.87144, -35.90665, -35.94107, 
        -35.97483, -36.00779, -36.03978, -36.07058, -36.10001, -36.12837, 
        -36.15572, -36.18312, -36.21065, -36.23899, -36.26786, -36.29683, 
        -36.32535, -36.35309, -36.38011, -36.40567, -36.4321, -36.45876, 
        -36.48592, -36.51367, -36.5419, -36.57026, -36.59858, -36.62659, 
        -36.65443, -36.68235, -36.71054, -36.73888, -36.76716, -36.7951, 
        -36.82232, -36.84928, -36.87588, -36.90262, -36.92939, -36.956, 
        -36.98125, -37.00704, -37.03269, -37.05856, -37.08496, -37.11219, 
        -37.14032, -37.16911, -37.19818, -37.22731, -37.25639, -37.28493, 
        -37.31311, -37.34083, -37.36776, -37.39437, -37.42072, -37.44717, 
        -37.47393, -37.50128, -37.52928, -37.55789, -37.5859, -37.61509, 
        -37.64429, -37.67352, -37.70279, -37.73206, -37.76127, -37.7899, 
        -37.81739, -37.8439, -37.86977, -37.89511, -37.91987, -37.94452, 
        -37.96894, -37.99306, -38.01672, -38.03984, -38.06266, -38.08532, 
        -38.1081, -38.13106, -38.15434, -38.17798, -38.20084, -38.22496, 
        -38.24911, -38.27306, -38.29579, -38.31777, -38.33894, -38.35889, 
        -38.37808, -38.39664, -38.41447, -38.4314, -38.44759, -38.46263, 
        -38.47664, -38.48991, -38.50283, -38.51585, -38.52933, -38.54369, 
        -38.55921, -38.57615, -38.5949, -38.61568, -38.63863, -38.66359, 
        -38.69004, -38.71701, -38.74264, -38.76821, -38.79255, -38.81567, 
        -38.83851, -38.86155, -38.88546, -38.91034, -38.9366, -38.96444, 
        -38.99383, -39.02437, -39.05564, -39.0873, -39.11897, -39.15052, 
        -39.18184, -39.2127, -39.24305, -39.27274, -39.30174, -39.33002, 
        -39.3576, -39.38441, -39.41035, -39.43541, -39.45966, -39.48281, 
        -39.50499, -39.52652, -39.54725, -39.56652, -39.5864, -39.60572, 
        -39.62479, -39.64297, -39.65965, -39.67406, -39.68578, -39.69482, 
        -39.70197, -39.70803, -39.71407, -39.72065, -39.72834, -39.73672, 
        -39.74533, -39.7533, -39.7603, -39.7658, -39.76983, -39.7722, 
        -39.77288, -39.77214, -39.77061, -39.76903, -39.76805, -39.76781, 
        -39.7681, -39.76826, -39.76742, -39.76458, -39.75885, -39.74971, 
        -39.73714, -39.72137, -39.70277, -39.68212, -39.65966, -39.63635, 
        -39.61267, -39.58758, -39.56313, -39.53771, -39.51035, -39.48027, 
        -39.44692, -39.41004, -39.36941, -39.32449, -39.27497, -39.22023, 
        -39.16029, -39.09523, -39.02603, -38.95455, -38.8835, -38.81589, 
        -38.75497,
  -31.03041, -31.07843, -31.12536, -31.17141, -31.21666, -31.26128, 
        -31.30564, -31.35012, -31.39553, -31.442, -31.48944, -31.53732, 
        -31.58388, -31.63043, -31.67577, -31.72008, -31.76373, -31.80727, 
        -31.85126, -31.89611, -31.94214, -31.98915, -32.03681, -32.08457, 
        -32.13209, -32.17926, -32.22506, -32.27163, -32.31804, -32.36423, 
        -32.41014, -32.45583, -32.50146, -32.54691, -32.59247, -32.63791, 
        -32.68356, -32.72914, -32.77493, -32.82089, -32.86742, -32.91476, 
        -32.96172, -33.01, -33.05833, -33.10657, -33.15502, -33.20394, 
        -33.25345, -33.30358, -33.35421, -33.40529, -33.45696, -33.50931, 
        -33.56234, -33.61592, -33.66985, -33.72397, -33.77721, -33.83132, 
        -33.88548, -33.93991, -33.99446, -34.0493, -34.1046, -34.16044, 
        -34.21688, -34.27377, -34.33094, -34.38814, -34.44502, -34.5013, 
        -34.55676, -34.61128, -34.66499, -34.71692, -34.76925, -34.82106, 
        -34.87244, -34.92306, -34.97257, -35.02042, -35.06662, -35.11125, 
        -35.15539, -35.19948, -35.24404, -35.28927, -35.33529, -35.38186, 
        -35.42825, -35.47432, -35.51875, -35.56375, -35.60791, -35.65113, 
        -35.69304, -35.73343, -35.77212, -35.80933, -35.84527, -35.88013, 
        -35.91405, -35.94698, -35.97882, -36.00946, -36.03893, -36.06732, 
        -36.09503, -36.12283, -36.151, -36.17902, -36.20848, -36.23796, 
        -36.267, -36.29541, -36.32328, -36.35088, -36.37848, -36.40617, 
        -36.4342, -36.46264, -36.49154, -36.52074, -36.54974, -36.57829, 
        -36.60649, -36.63445, -36.66246, -36.69065, -36.71882, -36.74559, 
        -36.77296, -36.79988, -36.82697, -36.85427, -36.8815, -36.90853, 
        -36.93521, -36.96156, -36.9879, -37.01405, -37.04063, -37.06785, 
        -37.09575, -37.12437, -37.15347, -37.18273, -37.21199, -37.24099, 
        -37.26962, -37.29776, -37.32521, -37.35117, -37.37803, -37.40493, 
        -37.43214, -37.4598, -37.48795, -37.51648, -37.54526, -37.57414, 
        -37.6031, -37.63229, -37.66162, -37.69093, -37.71988, -37.74804, 
        -37.77508, -37.80088, -37.82583, -37.85002, -37.8739, -37.89756, 
        -37.92107, -37.94433, -37.9661, -37.98834, -38.01021, -38.03202, 
        -38.05408, -38.07653, -38.09948, -38.12283, -38.14662, -38.1706, 
        -38.19486, -38.21867, -38.24177, -38.26367, -38.28436, -38.30416, 
        -38.32308, -38.34132, -38.35906, -38.37605, -38.39222, -38.40738, 
        -38.42171, -38.43533, -38.44879, -38.4623, -38.47529, -38.49012, 
        -38.5061, -38.52358, -38.543, -38.56477, -38.58886, -38.61511, 
        -38.64291, -38.67097, -38.69841, -38.7248, -38.74985, -38.77372, 
        -38.79712, -38.8208, -38.84543, -38.87117, -38.89794, -38.92624, 
        -38.95617, -38.98731, -39.01898, -39.05096, -39.08302, -39.11483, 
        -39.14655, -39.17777, -39.20811, -39.23754, -39.26607, -39.29279, 
        -39.31975, -39.34605, -39.37127, -39.39572, -39.41902, -39.44123, 
        -39.46289, -39.48393, -39.50459, -39.52501, -39.54521, -39.56483, 
        -39.58397, -39.60201, -39.61826, -39.63213, -39.6432, -39.65162, 
        -39.65783, -39.66323, -39.66867, -39.67493, -39.68252, -39.69102, 
        -39.6998, -39.70805, -39.71512, -39.72067, -39.7246, -39.72691, 
        -39.72762, -39.72693, -39.72551, -39.72401, -39.72305, -39.72166, 
        -39.72149, -39.72082, -39.71886, -39.71478, -39.70795, -39.69788, 
        -39.68428, -39.66761, -39.64843, -39.62704, -39.60435, -39.58024, 
        -39.55565, -39.53064, -39.50499, -39.4786, -39.45063, -39.42019, 
        -39.38648, -39.34924, -39.30742, -39.26108, -39.20966, -39.15298, 
        -39.09105, -39.02463, -38.95456, -38.88332, -38.8131, -38.74774, 
        -38.69093,
  -30.95835, -31.00634, -31.05335, -31.09928, -31.14445, -31.18904, 
        -31.23357, -31.27742, -31.32314, -31.36989, -31.41757, -31.46552, 
        -31.513, -31.55955, -31.6049, -31.64928, -31.69332, -31.73744, 
        -31.7821, -31.82762, -31.87414, -31.92135, -31.96807, -32.01579, 
        -32.06314, -32.10992, -32.15627, -32.20241, -32.24839, -32.29427, 
        -32.33998, -32.38544, -32.43094, -32.4766, -32.52227, -32.56805, 
        -32.6141, -32.65909, -32.70531, -32.7519, -32.7991, -32.84718, 
        -32.89597, -32.9451, -32.99429, -33.04343, -33.09275, -33.14253, 
        -33.19291, -33.2439, -33.29547, -33.34734, -33.39959, -33.45135, 
        -33.50471, -33.55859, -33.61277, -33.66698, -33.72121, -33.77544, 
        -33.82981, -33.88441, -33.93925, -33.99435, -34.04978, -34.10564, 
        -34.16176, -34.21818, -34.27451, -34.32975, -34.3857, -34.44111, 
        -34.496, -34.55035, -34.60407, -34.6572, -34.70971, -34.76177, 
        -34.81332, -34.86417, -34.91376, -34.96139, -35.00694, -35.05077, 
        -35.09383, -35.13691, -35.17969, -35.22451, -35.27036, -35.31667, 
        -35.36289, -35.40874, -35.45375, -35.49847, -35.54263, -35.58608, 
        -35.62844, -35.66942, -35.70903, -35.74712, -35.78381, -35.81924, 
        -35.85351, -35.88665, -35.9187, -35.94851, -35.97818, -36.0069, 
        -36.03509, -36.06339, -36.09222, -36.1218, -36.15175, -36.18164, 
        -36.21104, -36.23991, -36.26844, -36.29694, -36.32549, -36.35411, 
        -36.38287, -36.41215, -36.44176, -36.47148, -36.50011, -36.52925, 
        -36.5578, -36.5858, -36.61371, -36.64151, -36.66932, -36.69697, 
        -36.72437, -36.75169, -36.77929, -36.80718, -36.83499, -36.86263, 
        -36.88992, -36.91677, -36.94348, -36.97024, -36.99707, -37.02425, 
        -37.05203, -37.07944, -37.10836, -37.1376, -37.16692, -37.19612, 
        -37.22509, -37.25361, -37.2816, -37.30917, -37.33658, -37.36397, 
        -37.39161, -37.41947, -37.44775, -37.47612, -37.50473, -37.53336, 
        -37.56214, -37.59122, -37.62045, -37.64955, -37.67812, -37.70568, 
        -37.73097, -37.75602, -37.78004, -37.80339, -37.82644, -37.84938, 
        -37.87222, -37.8948, -37.91692, -37.93841, -37.95951, -37.98057, 
        -38.00188, -38.02352, -38.04586, -38.06887, -38.09231, -38.11617, 
        -38.14014, -38.16381, -38.18679, -38.20854, -38.22916, -38.24878, 
        -38.26752, -38.28574, -38.30243, -38.31949, -38.33577, -38.35121, 
        -38.36596, -38.38021, -38.39428, -38.40844, -38.42301, -38.43827, 
        -38.45467, -38.47263, -38.49269, -38.51531, -38.54075, -38.56808, 
        -38.59688, -38.6259, -38.65446, -38.68182, -38.70762, -38.7323, 
        -38.7565, -38.78075, -38.80601, -38.83215, -38.8594, -38.88821, 
        -38.91754, -38.9491, -38.98122, -39.01355, -39.04588, -39.07808, 
        -39.11003, -39.14147, -39.17189, -39.20103, -39.22921, -39.25641, 
        -39.28273, -39.30824, -39.33262, -39.35594, -39.37836, -39.39983, 
        -39.42083, -39.44159, -39.46222, -39.48282, -39.50331, -39.5233, 
        -39.54247, -39.5603, -39.57615, -39.58944, -39.59993, -39.60775, 
        -39.61343, -39.61823, -39.62325, -39.62925, -39.6357, -39.64429, 
        -39.65323, -39.66162, -39.66876, -39.67433, -39.67817, -39.68042, 
        -39.68107, -39.68047, -39.67912, -39.6776, -39.67675, -39.67616, 
        -39.67554, -39.67387, -39.6706, -39.66522, -39.65715, -39.64603, 
        -39.63175, -39.61452, -39.59497, -39.57364, -39.55058, -39.52628, 
        -39.50092, -39.47469, -39.44765, -39.41998, -39.39094, -39.35981, 
        -39.32574, -39.28774, -39.24492, -39.19726, -39.14426, -39.08591, 
        -39.02254, -38.95477, -38.88464, -38.81368, -38.74546, -38.68307, 
        -38.63079,
  -30.88737, -30.93547, -30.98248, -31.02746, -31.07261, -31.11732, 
        -31.162, -31.20726, -31.25344, -31.3005, -31.34835, -31.39634, 
        -31.44386, -31.49038, -31.53584, -31.58041, -31.62492, -31.66884, 
        -31.71432, -31.76062, -31.80765, -31.85515, -31.90289, -31.95049, 
        -31.99758, -32.04409, -32.09002, -32.13565, -32.18118, -32.22668, 
        -32.27211, -32.31749, -32.36201, -32.40782, -32.45387, -32.5001, 
        -32.54644, -32.59284, -32.63937, -32.68641, -32.73418, -32.78286, 
        -32.83257, -32.88263, -32.93283, -32.98292, -33.03316, -33.08286, 
        -33.13412, -33.18597, -33.2382, -33.2907, -33.34338, -33.39642, 
        -33.44995, -33.50398, -33.55825, -33.61251, -33.66668, -33.72096, 
        -33.77554, -33.83041, -33.88567, -33.94111, -33.99572, -34.05167, 
        -34.10769, -34.16335, -34.21896, -34.27414, -34.32891, -34.38336, 
        -34.43745, -34.49133, -34.5449, -34.59803, -34.65061, -34.70269, 
        -34.75426, -34.80531, -34.85524, -34.90189, -34.9473, -34.99069, 
        -35.03316, -35.07558, -35.11882, -35.16327, -35.20894, -35.25475, 
        -35.30046, -35.3457, -35.39004, -35.43421, -35.4781, -35.52151, 
        -35.56405, -35.60552, -35.64575, -35.68367, -35.72117, -35.7573, 
        -35.79206, -35.82563, -35.85808, -35.8894, -35.91961, -35.94891, 
        -35.97773, -36.00665, -36.03612, -36.06624, -36.09667, -36.12675, 
        -36.1563, -36.1854, -36.21439, -36.2435, -36.27187, -36.30127, 
        -36.33076, -36.36038, -36.39066, -36.42121, -36.45146, -36.48104, 
        -36.5099, -36.53797, -36.56561, -36.59314, -36.62061, -36.64814, 
        -36.6757, -36.70352, -36.7318, -36.76024, -36.78871, -36.81691, 
        -36.84365, -36.87107, -36.89832, -36.92543, -36.95267, -36.98001, 
        -37.00776, -37.03598, -37.0647, -37.09381, -37.12299, -37.15218, 
        -37.18128, -37.2102, -37.2388, -37.267, -37.29494, -37.3228, 
        -37.3507, -37.37878, -37.40704, -37.43532, -37.4636, -37.49092, 
        -37.51962, -37.5486, -37.57767, -37.60657, -37.63464, -37.66146, 
        -37.68698, -37.71113, -37.73422, -37.75691, -37.77945, -37.80199, 
        -37.8244, -37.84651, -37.86814, -37.88916, -37.90966, -37.9301, 
        -37.95056, -37.97153, -37.99309, -38.01543, -38.03847, -38.06093, 
        -38.08459, -38.10803, -38.13079, -38.15251, -38.17302, -38.19246, 
        -38.21107, -38.22923, -38.24695, -38.26406, -38.28062, -38.29646, 
        -38.31168, -38.32671, -38.34149, -38.35648, -38.37167, -38.38745, 
        -38.40435, -38.42284, -38.44355, -38.46693, -38.49317, -38.52151, 
        -38.55143, -38.58151, -38.61106, -38.63832, -38.6651, -38.69064, 
        -38.71557, -38.74068, -38.76635, -38.79288, -38.82051, -38.84964, 
        -38.88017, -38.91197, -38.94439, -38.97706, -39.0097, -39.04216, 
        -39.07423, -39.10564, -39.13612, -39.16527, -39.19299, -39.21965, 
        -39.24531, -39.26987, -39.2933, -39.31558, -39.33692, -39.35766, 
        -39.37807, -39.39859, -39.41928, -39.44012, -39.46082, -39.48002, 
        -39.49918, -39.51672, -39.53215, -39.54496, -39.55502, -39.56249, 
        -39.56792, -39.5725, -39.57716, -39.58298, -39.59022, -39.59883, 
        -39.60777, -39.61619, -39.62325, -39.62887, -39.63266, -39.6347, 
        -39.63523, -39.63475, -39.63345, -39.63193, -39.63102, -39.63012, 
        -39.62873, -39.62608, -39.62157, -39.61483, -39.60554, -39.59345, 
        -39.57855, -39.56113, -39.54164, -39.52033, -39.49757, -39.47311, 
        -39.44708, -39.41956, -39.39099, -39.36066, -39.3303, -39.29824, 
        -39.26344, -39.22494, -39.18151, -39.13263, -39.07841, -39.0187, 
        -38.95422, -38.88593, -38.81573, -38.7459, -38.67991, -38.62149, 
        -38.57344,
  -30.81649, -30.86468, -30.91181, -30.95787, -31.00318, -31.04811, 
        -31.09325, -31.13898, -31.18552, -31.23286, -31.28079, -31.32879, 
        -31.3754, -31.42206, -31.46774, -31.51278, -31.55785, -31.60346, 
        -31.64989, -31.69693, -31.74434, -31.79209, -31.83983, -31.88726, 
        -31.93423, -31.98054, -32.02606, -32.07017, -32.11519, -32.16026, 
        -32.2054, -32.25066, -32.29644, -32.34265, -32.38914, -32.43593, 
        -32.48269, -32.52943, -32.57626, -32.62352, -32.67186, -32.72123, 
        -32.77065, -32.82179, -32.87298, -32.9241, -32.97531, -33.02691, 
        -33.079, -33.13162, -33.18452, -33.23747, -33.29044, -33.34358, 
        -33.39705, -33.45096, -33.50512, -33.55931, -33.61248, -33.66678, 
        -33.72155, -33.77684, -33.8324, -33.88828, -33.94424, -34.00029, 
        -34.05596, -34.11135, -34.16645, -34.22036, -34.27394, -34.32729, 
        -34.38037, -34.43354, -34.48659, -34.53851, -34.59094, -34.6427, 
        -34.69466, -34.74579, -34.79548, -34.84347, -34.88924, -34.9327, 
        -34.97519, -35.01764, -35.06071, -35.10479, -35.1498, -35.19509, 
        -35.24007, -35.28421, -35.32792, -35.37056, -35.41392, -35.45702, 
        -35.49952, -35.54103, -35.58164, -35.62109, -35.65927, -35.69605, 
        -35.73151, -35.76571, -35.79882, -35.83089, -35.86179, -35.89178, 
        -35.9213, -35.95097, -35.98114, -36.01172, -36.04142, -36.07164, 
        -36.10122, -36.13029, -36.15954, -36.18914, -36.21904, -36.24901, 
        -36.27914, -36.30941, -36.34028, -36.37133, -36.40213, -36.4322, 
        -36.46124, -36.48933, -36.51675, -36.54396, -36.57136, -36.59886, 
        -36.62568, -36.65405, -36.683, -36.71218, -36.74118, -36.76982, 
        -36.798, -36.82583, -36.85356, -36.88123, -36.90887, -36.93655, 
        -36.96443, -36.99259, -37.02113, -37.04996, -37.07889, -37.10798, 
        -37.13719, -37.16639, -37.19551, -37.22325, -37.25171, -37.27993, 
        -37.30807, -37.33619, -37.36431, -37.39233, -37.42031, -37.44836, 
        -37.4768, -37.50563, -37.53456, -37.56303, -37.59064, -37.6169, 
        -37.6416, -37.66497, -37.68752, -37.70964, -37.73189, -37.75418, 
        -37.77636, -37.79818, -37.81944, -37.8391, -37.85925, -37.87916, 
        -37.89899, -37.91916, -37.93993, -37.96151, -37.98391, -38.00688, 
        -38.03022, -38.05343, -38.07608, -38.0978, -38.11827, -38.13764, 
        -38.15619, -38.17421, -38.19194, -38.20908, -38.2258, -38.24215, 
        -38.25805, -38.27357, -38.28949, -38.30516, -38.32116, -38.3367, 
        -38.35431, -38.37347, -38.39491, -38.4189, -38.44578, -38.47509, 
        -38.50572, -38.5369, -38.56739, -38.59669, -38.62456, -38.65127, 
        -38.67722, -38.70284, -38.72893, -38.7557, -38.78349, -38.81264, 
        -38.84324, -38.87514, -38.90778, -38.94065, -38.97347, -39.00604, 
        -39.03816, -39.0695, -39.09982, -39.12878, -39.15634, -39.18246, 
        -39.20616, -39.22992, -39.25222, -39.27328, -39.29379, -39.31381, 
        -39.33379, -39.35427, -39.37508, -39.39613, -39.41712, -39.43742, 
        -39.45635, -39.47352, -39.48848, -39.5009, -39.51073, -39.51816, 
        -39.52358, -39.52815, -39.53282, -39.53849, -39.54568, -39.55396, 
        -39.56254, -39.57086, -39.57787, -39.58329, -39.58704, -39.58915, 
        -39.58979, -39.58924, -39.58789, -39.58636, -39.58508, -39.58354, 
        -39.58136, -39.5766, -39.57089, -39.56291, -39.55255, -39.53962, 
        -39.52419, -39.50661, -39.48718, -39.46634, -39.44397, -39.41951, 
        -39.39289, -39.36411, -39.33381, -39.30283, -39.27087, -39.23774, 
        -39.20211, -39.16292, -39.11914, -39.06974, -39.01464, -38.95408, 
        -38.88895, -38.82038, -38.75061, -38.68235, -38.61911, -38.56446, 
        -38.52071,
  -30.74783, -30.79609, -30.84331, -30.88962, -30.93523, -30.98065, 
        -31.02634, -31.07253, -31.11839, -31.16588, -31.21386, -31.26194, 
        -31.30961, -31.35653, -31.40255, -31.44817, -31.49387, -31.54035, 
        -31.58746, -31.63509, -31.68292, -31.73065, -31.77728, -31.82489, 
        -31.87177, -31.91772, -31.96286, -32.00749, -32.05194, -32.09655, 
        -32.1414, -32.18677, -32.23273, -32.27965, -32.32691, -32.37442, 
        -32.4217, -32.46785, -32.51495, -32.56263, -32.6115, -32.66167, 
        -32.71287, -32.76479, -32.8169, -32.86898, -32.92107, -32.97356, 
        -33.02639, -33.07964, -33.13306, -33.18639, -33.23952, -33.29166, 
        -33.345, -33.3986, -33.45247, -33.50647, -33.56054, -33.61496, 
        -33.67, -33.72562, -33.78163, -33.83795, -33.89416, -33.95026, 
        -34.00573, -34.06062, -34.11463, -34.16808, -34.21956, -34.27179, 
        -34.32401, -34.37626, -34.4286, -34.48097, -34.53303, -34.58501, 
        -34.6362, -34.68705, -34.73709, -34.78556, -34.83147, -34.87573, 
        -34.9189, -34.96183, -35.00502, -35.04779, -35.09202, -35.13623, 
        -35.17997, -35.22322, -35.26608, -35.3091, -35.35231, -35.39504, 
        -35.43706, -35.47842, -35.51905, -35.55878, -35.59739, -35.63481, 
        -35.67089, -35.70581, -35.73967, -35.7725, -35.80309, -35.83387, 
        -35.86418, -35.89453, -35.92525, -35.95633, -35.98721, -36.01745, 
        -36.04692, -36.07601, -36.10531, -36.13512, -36.16545, -36.196, 
        -36.22651, -36.2575, -36.28886, -36.3205, -36.35176, -36.38121, 
        -36.4104, -36.43844, -36.46577, -36.49298, -36.52011, -36.54778, 
        -36.57605, -36.60509, -36.63464, -36.66443, -36.69401, -36.72306, 
        -36.75154, -36.77978, -36.80783, -36.83591, -36.86404, -36.89221, 
        -36.92046, -36.94879, -36.97632, -37.00491, -37.03362, -37.06257, 
        -37.09185, -37.12123, -37.15069, -37.17988, -37.20871, -37.23718, 
        -37.26541, -37.29345, -37.3213, -37.34895, -37.37654, -37.40418, 
        -37.4322, -37.46068, -37.4894, -37.51754, -37.5448, -37.5704, 
        -37.59465, -37.61641, -37.63857, -37.66056, -37.68269, -37.70484, 
        -37.72671, -37.74828, -37.76929, -37.7897, -37.80956, -37.82905, 
        -37.84838, -37.86791, -37.88794, -37.9087, -37.93048, -37.95291, 
        -37.97594, -37.99892, -38.02161, -38.04348, -38.06415, -38.08361, 
        -38.10215, -38.1201, -38.13662, -38.15375, -38.17055, -38.18712, 
        -38.20368, -38.22005, -38.23684, -38.25325, -38.27029, -38.28777, 
        -38.30634, -38.3264, -38.3486, -38.37354, -38.40112, -38.43103, 
        -38.46231, -38.49431, -38.5258, -38.55619, -38.58531, -38.61316, 
        -38.63986, -38.66636, -38.69272, -38.71947, -38.74728, -38.77629, 
        -38.80672, -38.83764, -38.87037, -38.90334, -38.93621, -38.96873, 
        -39.00064, -39.0318, -39.06201, -39.09079, -39.11792, -39.14357, 
        -39.16772, -39.19033, -39.21137, -39.23146, -39.25119, -39.27061, 
        -39.29065, -39.3111, -39.33212, -39.35332, -39.37426, -39.39452, 
        -39.41321, -39.42979, -39.44436, -39.45665, -39.46641, -39.47391, 
        -39.47966, -39.48445, -39.4893, -39.49507, -39.50196, -39.50994, 
        -39.5172, -39.52492, -39.53154, -39.53664, -39.54041, -39.54271, 
        -39.54357, -39.5432, -39.54189, -39.54023, -39.5384, -39.53609, 
        -39.53283, -39.52801, -39.52111, -39.51213, -39.50085, -39.48715, 
        -39.47116, -39.45342, -39.43419, -39.41367, -39.39151, -39.3671, 
        -39.33986, -39.30983, -39.27792, -39.24531, -39.21185, -39.17731, 
        -39.14115, -39.1015, -39.05739, -39.00783, -38.95243, -38.89147, 
        -38.82599, -38.75746, -38.6882, -38.62151, -38.56087, -38.50986, 
        -38.47039,
  -30.68072, -30.72887, -30.77631, -30.82193, -30.86803, -30.91403, 
        -30.96027, -31.00693, -31.05407, -31.10169, -31.14966, -31.19772, 
        -31.24547, -31.29261, -31.3391, -31.38523, -31.43181, -31.47897, 
        -31.52565, -31.57373, -31.62179, -31.66961, -31.7175, -31.76487, 
        -31.81173, -31.85746, -31.90216, -31.94628, -31.99021, -32.03439, 
        -32.07911, -32.12473, -32.17042, -32.21802, -32.26619, -32.31442, 
        -32.36234, -32.40997, -32.4577, -32.50607, -32.55555, -32.60636, 
        -32.65831, -32.71072, -32.76351, -32.8163, -32.86911, -32.92234, 
        -32.9748, -33.02861, -33.08244, -33.1361, -33.18945, -33.2426, 
        -33.29573, -33.34901, -33.40243, -33.45614, -33.5101, -33.5646, 
        -33.61988, -33.67587, -33.73231, -33.78876, -33.84392, -33.89971, 
        -33.95493, -34.00921, -34.06257, -34.1151, -34.16693, -34.21849, 
        -34.26979, -34.32137, -34.37321, -34.42508, -34.47687, -34.52837, 
        -34.57943, -34.63004, -34.67949, -34.72714, -34.77369, -34.81885, 
        -34.86296, -34.90636, -34.94958, -34.99286, -35.03615, -35.07916, 
        -35.12165, -35.16381, -35.20602, -35.24858, -35.2914, -35.33386, 
        -35.37555, -35.41669, -35.45724, -35.49598, -35.53476, -35.57257, 
        -35.60909, -35.64462, -35.67923, -35.7126, -35.74503, -35.77659, 
        -35.8076, -35.83858, -35.86978, -35.90105, -35.93208, -35.96241, 
        -35.99192, -36.02111, -36.05054, -36.08052, -36.11106, -36.14093, 
        -36.17204, -36.20357, -36.2355, -36.26756, -36.29921, -36.32988, 
        -36.35934, -36.38752, -36.41494, -36.44204, -36.46933, -36.49717, 
        -36.526, -36.55554, -36.58562, -36.61586, -36.64582, -36.67521, 
        -36.70402, -36.73148, -36.75999, -36.78839, -36.81686, -36.84549, 
        -36.87417, -36.90294, -36.93169, -36.96042, -36.98922, -37.01819, 
        -37.04744, -37.07693, -37.10662, -37.13604, -37.16507, -37.19366, 
        -37.22177, -37.24951, -37.27694, -37.30407, -37.33107, -37.35713, 
        -37.38463, -37.41268, -37.44101, -37.46908, -37.49591, -37.52156, 
        -37.5456, -37.56841, -37.59032, -37.6121, -37.63387, -37.65567, 
        -37.67722, -37.69853, -37.71931, -37.73948, -37.75909, -37.77825, 
        -37.79726, -37.81634, -37.83591, -37.85616, -37.87721, -37.89936, 
        -37.92099, -37.94389, -37.9666, -37.98857, -38.00944, -38.029, 
        -38.0476, -38.06557, -38.08294, -38.10003, -38.11696, -38.13375, 
        -38.15076, -38.16803, -38.18539, -38.20308, -38.22106, -38.23966, 
        -38.25927, -38.28034, -38.3036, -38.32938, -38.3577, -38.38843, 
        -38.42047, -38.45296, -38.48526, -38.5166, -38.54573, -38.57447, 
        -38.60192, -38.62896, -38.65551, -38.68244, -38.71021, -38.73898, 
        -38.76933, -38.80117, -38.8338, -38.86692, -38.89964, -38.93197, 
        -38.96373, -38.99469, -39.02463, -39.05334, -39.08038, -39.10567, 
        -39.12914, -39.15097, -39.17123, -39.19041, -39.20956, -39.22876, 
        -39.24848, -39.26897, -39.28989, -39.31087, -39.33152, -39.35131, 
        -39.36844, -39.38473, -39.39897, -39.41093, -39.42082, -39.42877, 
        -39.43505, -39.44041, -39.44566, -39.45169, -39.45863, -39.46618, 
        -39.474, -39.48106, -39.48717, -39.49182, -39.49547, -39.49788, 
        -39.49892, -39.49873, -39.49755, -39.49574, -39.49341, -39.49033, 
        -39.48603, -39.48002, -39.47203, -39.46209, -39.44984, -39.43555, 
        -39.41908, -39.40106, -39.38187, -39.36139, -39.33916, -39.31433, 
        -39.2863, -39.2552, -39.22203, -39.18768, -39.15289, -39.11649, 
        -39.07967, -39.04001, -38.99583, -38.94628, -38.89086, -38.82976, 
        -38.76402, -38.69541, -38.62659, -38.56103, -38.50242, -38.45415, 
        -38.41802,
  -30.61428, -30.66241, -30.70996, -30.75695, -30.8036, -30.85018, 
        -30.89697, -30.94406, -30.99138, -31.03904, -31.08694, -31.13489, 
        -31.1826, -31.22888, -31.27588, -31.32268, -31.36993, -31.41765, 
        -31.46604, -31.5144, -31.56267, -31.61063, -31.65865, -31.70604, 
        -31.75272, -31.79824, -31.84266, -31.88635, -31.92894, -31.97293, 
        -32.01761, -32.06367, -32.11091, -32.15936, -32.20848, -32.25758, 
        -32.30627, -32.3546, -32.40305, -32.45223, -32.50252, -32.554, 
        -32.60653, -32.65841, -32.71157, -32.76482, -32.81829, -32.8721, 
        -32.92607, -32.98026, -33.03443, -33.08837, -33.14194, -33.19516, 
        -33.24813, -33.30098, -33.35392, -33.40722, -33.46092, -33.51448, 
        -33.57001, -33.62619, -33.68269, -33.73908, -33.7951, -33.85045, 
        -33.90506, -33.95879, -34.01164, -34.06368, -34.11507, -34.16608, 
        -34.21696, -34.26799, -34.31938, -34.37067, -34.42109, -34.47236, 
        -34.52293, -34.57308, -34.62246, -34.67078, -34.71793, -34.76384, 
        -34.80868, -34.85259, -34.89577, -34.93834, -34.98047, -35.02213, 
        -35.0633, -35.10451, -35.14624, -35.18857, -35.23014, -35.27241, 
        -35.31414, -35.35511, -35.39512, -35.43469, -35.4736, -35.51139, 
        -35.54818, -35.58409, -35.61904, -35.65304, -35.68611, -35.71835, 
        -35.75005, -35.7816, -35.81316, -35.84459, -35.87463, -35.90512, 
        -35.93483, -35.96422, -35.99383, -36.02396, -36.05466, -36.08584, 
        -36.11746, -36.1495, -36.18188, -36.21429, -36.24623, -36.27722, 
        -36.307, -36.33554, -36.36319, -36.39044, -36.41796, -36.44627, 
        -36.4744, -36.50441, -36.53493, -36.56553, -36.59578, -36.62547, 
        -36.65467, -36.68322, -36.71181, -36.74049, -36.76933, -36.79837, 
        -36.82754, -36.85688, -36.88614, -36.9153, -36.94443, -36.97363, 
        -37.00305, -37.03267, -37.06236, -37.09187, -37.11995, -37.14844, 
        -37.17622, -37.20345, -37.23021, -37.25665, -37.2828, -37.30921, 
        -37.33604, -37.36356, -37.39147, -37.41925, -37.44626, -37.472, 
        -37.49623, -37.51921, -37.54119, -37.56273, -37.58409, -37.6055, 
        -37.62688, -37.64776, -37.66822, -37.68811, -37.70653, -37.72556, 
        -37.74448, -37.76335, -37.78251, -37.80231, -37.82308, -37.84467, 
        -37.86686, -37.8897, -37.91241, -37.93446, -37.95549, -37.97524, 
        -37.99394, -38.01168, -38.02894, -38.046, -38.06302, -38.0803, 
        -38.09797, -38.11597, -38.13421, -38.15276, -38.17178, -38.19157, 
        -38.21151, -38.23391, -38.25833, -38.28531, -38.31467, -38.34601, 
        -38.37878, -38.41187, -38.44477, -38.47686, -38.50762, -38.53701, 
        -38.56519, -38.59239, -38.61927, -38.64633, -38.67401, -38.70256, 
        -38.73271, -38.76434, -38.79704, -38.82996, -38.86273, -38.89482, 
        -38.92627, -38.95697, -38.98677, -39.01535, -39.04232, -39.06738, 
        -39.09046, -39.11065, -39.13015, -39.1489, -39.16784, -39.18696, 
        -39.20671, -39.22703, -39.24755, -39.26806, -39.28806, -39.30709, 
        -39.32457, -39.34035, -39.35414, -39.36598, -39.37614, -39.38464, 
        -39.39171, -39.39785, -39.40377, -39.41005, -39.41713, -39.42458, 
        -39.4317, -39.43818, -39.44353, -39.44778, -39.451, -39.45335, 
        -39.45454, -39.45461, -39.45367, -39.4518, -39.44907, -39.44526, 
        -39.44, -39.43298, -39.423, -39.41204, -39.39917, -39.38407, 
        -39.36723, -39.34896, -39.32956, -39.30878, -39.28611, -39.26068, 
        -39.23173, -39.19953, -39.16513, -39.12971, -39.09406, -39.05796, 
        -39.02088, -38.98123, -38.93732, -38.88792, -38.83239, -38.77084, 
        -38.7045, -38.63532, -38.56623, -38.50109, -38.44379, -38.3975, 
        -38.36415,
  -30.55063, -30.59861, -30.64628, -30.69366, -30.74087, -30.78801, 
        -30.83531, -30.88271, -30.92922, -30.97686, -31.0246, -31.0723, 
        -31.11982, -31.1671, -31.21434, -31.26172, -31.30962, -31.35816, 
        -31.40693, -31.4558, -31.50444, -31.5528, -31.60088, -31.64744, 
        -31.694, -31.7393, -31.78345, -31.8269, -31.87033, -31.91433, 
        -31.95942, -32.00585, -32.05389, -32.10321, -32.15322, -32.20314, 
        -32.25257, -32.30165, -32.34991, -32.3999, -32.45095, -32.50301, 
        -32.55587, -32.60904, -32.66251, -32.71622, -32.77024, -32.82451, 
        -32.87893, -32.93342, -32.98786, -33.04209, -33.09588, -33.14916, 
        -33.20095, -33.2534, -33.30577, -33.35856, -33.41193, -33.46649, 
        -33.52198, -33.57818, -33.63456, -33.69068, -33.74621, -33.80101, 
        -33.85495, -33.90815, -33.96061, -34.01234, -34.06252, -34.1134, 
        -34.16409, -34.21484, -34.26568, -34.31675, -34.36781, -34.41878, 
        -34.46896, -34.51835, -34.56743, -34.6155, -34.66294, -34.70926, 
        -34.7547, -34.79873, -34.84166, -34.88348, -34.92337, -34.96362, 
        -35.00346, -35.04386, -35.0856, -35.1279, -35.17041, -35.21258, 
        -35.25404, -35.29472, -35.3347, -35.37413, -35.41269, -35.45039, 
        -35.48718, -35.52314, -35.55824, -35.59264, -35.62523, -35.6581, 
        -35.69046, -35.72251, -35.75436, -35.78588, -35.81713, -35.84771, 
        -35.8777, -35.90746, -35.9374, -35.9677, -35.99856, -36.03005, 
        -36.06215, -36.09466, -36.12735, -36.15998, -36.19205, -36.22334, 
        -36.25259, -36.28172, -36.3099, -36.33757, -36.36546, -36.39407, 
        -36.42358, -36.45387, -36.48465, -36.51555, -36.54591, -36.57584, 
        -36.60533, -36.63413, -36.66304, -36.69182, -36.72076, -36.75011, 
        -36.77979, -36.80965, -36.83953, -36.86827, -36.89804, -36.92773, 
        -36.95741, -36.98715, -37.01683, -37.04636, -37.07537, -37.10365, 
        -37.131, -37.15753, -37.1834, -37.20886, -37.23407, -37.25959, 
        -37.28571, -37.3126, -37.34009, -37.36766, -37.39479, -37.42088, 
        -37.44565, -37.46904, -37.49024, -37.51167, -37.53276, -37.55373, 
        -37.57455, -37.59506, -37.61525, -37.63496, -37.6543, -37.67333, 
        -37.69225, -37.71112, -37.73016, -37.74969, -37.76994, -37.7911, 
        -37.81291, -37.83531, -37.85782, -37.87975, -37.90071, -37.92052, 
        -37.93897, -37.95672, -37.97367, -37.98963, -38.00695, -38.0248, 
        -38.04336, -38.06242, -38.08184, -38.10151, -38.12171, -38.14267, 
        -38.16479, -38.18854, -38.21432, -38.24256, -38.27322, -38.30552, 
        -38.33888, -38.37256, -38.40586, -38.43826, -38.46944, -38.49923, 
        -38.5278, -38.55544, -38.58249, -38.60947, -38.63708, -38.66569, 
        -38.69568, -38.72717, -38.75872, -38.79168, -38.82433, -38.85631, 
        -38.88757, -38.91797, -38.94759, -38.97608, -39.00296, -39.02793, 
        -39.0508, -39.07169, -39.09108, -39.10966, -39.12837, -39.14757, 
        -39.16733, -39.18723, -39.20716, -39.22673, -39.24577, -39.26389, 
        -39.28061, -39.2957, -39.30909, -39.32096, -39.33145, -39.34058, 
        -39.34853, -39.35562, -39.36233, -39.36917, -39.37627, -39.3835, 
        -39.39019, -39.39493, -39.39957, -39.40323, -39.40612, -39.4082, 
        -39.40941, -39.40968, -39.40895, -39.4072, -39.40417, -39.39972, 
        -39.39362, -39.38568, -39.37581, -39.36414, -39.35053, -39.33496, 
        -39.31793, -39.29939, -39.27956, -39.25836, -39.23503, -39.20863, 
        -39.17873, -39.14565, -39.1104, -39.07428, -39.03795, -39.00157, 
        -38.96447, -38.92495, -38.88138, -38.83197, -38.77594, -38.71361, 
        -38.64601, -38.57547, -38.50527, -38.43954, -38.38247, -38.33745, 
        -38.30629,
  -30.48868, -30.53646, -30.58419, -30.63188, -30.67859, -30.72624, 
        -30.77404, -30.82185, -30.86956, -30.91716, -30.96463, -31.01193, 
        -31.05907, -31.10623, -31.15364, -31.20148, -31.24995, -31.29899, 
        -31.34742, -31.39689, -31.44614, -31.49506, -31.54345, -31.59101, 
        -31.63747, -31.68268, -31.72677, -31.77019, -31.81389, -31.85815, 
        -31.9038, -31.95081, -31.99954, -32.04866, -32.09948, -32.1501, 
        -32.2003, -32.25017, -32.30022, -32.3508, -32.40241, -32.45478, 
        -32.50774, -32.56112, -32.61485, -32.66895, -32.72348, -32.77826, 
        -32.83311, -32.88693, -32.94156, -32.99595, -33.04992, -33.1032, 
        -33.15578, -33.20783, -33.25974, -33.31193, -33.36487, -33.41916, 
        -33.47432, -33.53043, -33.58639, -33.64208, -33.69716, -33.7503, 
        -33.80358, -33.85618, -33.90826, -33.95977, -34.01084, -34.06171, 
        -34.11244, -34.16325, -34.21416, -34.26507, -34.31556, -34.36595, 
        -34.41557, -34.46479, -34.51297, -34.56086, -34.60729, -34.65368, 
        -34.69919, -34.74318, -34.78554, -34.82656, -34.86617, -34.90551, 
        -34.94463, -34.98477, -35.02614, -35.06847, -35.11094, -35.15302, 
        -35.19439, -35.235, -35.2748, -35.31398, -35.35123, -35.38869, 
        -35.42533, -35.4611, -35.49622, -35.53071, -35.56474, -35.59818, 
        -35.63116, -35.66366, -35.69582, -35.72753, -35.75891, -35.78971, 
        -35.82015, -35.85036, -35.88062, -35.91117, -35.94226, -35.97308, 
        -36.00561, -36.03857, -36.0715, -36.10405, -36.13622, -36.16771, 
        -36.19844, -36.22826, -36.25721, -36.28549, -36.31374, -36.34271, 
        -36.37243, -36.40288, -36.43368, -36.46463, -36.49521, -36.52537, 
        -36.55516, -36.58429, -36.6124, -36.64124, -36.67052, -36.70024, 
        -36.73033, -36.7607, -36.79121, -36.82162, -36.85199, -36.88223, 
        -36.91227, -36.94218, -36.97193, -37.00138, -37.03026, -37.05825, 
        -37.0851, -37.11087, -37.1357, -37.16002, -37.18424, -37.20892, 
        -37.23329, -37.25937, -37.28637, -37.3137, -37.34094, -37.36749, 
        -37.3929, -37.41692, -37.43948, -37.46103, -37.48178, -37.50219, 
        -37.52248, -37.54268, -37.56258, -37.58221, -37.6016, -37.62081, 
        -37.6399, -37.6588, -37.67793, -37.69732, -37.7172, -37.73775, 
        -37.75904, -37.77981, -37.80168, -37.82311, -37.84363, -37.86298, 
        -37.8813, -37.89858, -37.91549, -37.93251, -37.95024, -37.96893, 
        -37.98869, -38.00909, -38.02986, -38.05079, -38.07235, -38.09452, 
        -38.11788, -38.14293, -38.17006, -38.19976, -38.23173, -38.26515, 
        -38.29927, -38.33344, -38.36705, -38.39958, -38.4309, -38.46001, 
        -38.48887, -38.51671, -38.5439, -38.57102, -38.59865, -38.62727, 
        -38.65727, -38.68867, -38.72116, -38.75409, -38.78677, -38.81874, 
        -38.84986, -38.88013, -38.90953, -38.93781, -38.96445, -38.98927, 
        -39.01208, -39.033, -39.05249, -39.07128, -39.09015, -39.10939, 
        -39.12884, -39.14832, -39.16736, -39.18592, -39.2039, -39.22104, 
        -39.237, -39.25051, -39.26359, -39.27544, -39.28634, -39.29604, 
        -39.30479, -39.3127, -39.32021, -39.32755, -39.33481, -39.34174, 
        -39.34793, -39.35308, -39.35715, -39.36029, -39.36283, -39.36465, 
        -39.36568, -39.36604, -39.36544, -39.36361, -39.36036, -39.35539, 
        -39.34859, -39.3399, -39.32932, -39.3169, -39.30283, -39.28705, 
        -39.26981, -39.25119, -39.23137, -39.20956, -39.18554, -39.15825, 
        -39.12748, -39.09367, -39.0578, -39.02127, -38.98464, -38.9482, 
        -38.91026, -38.87096, -38.82698, -38.77731, -38.72068, -38.65696, 
        -38.58724, -38.5145, -38.44219, -38.37486, -38.31701, -38.2723, 
        -38.24287,
  -30.42707, -30.47463, -30.52241, -30.57037, -30.61837, -30.66657, 
        -30.71488, -30.76318, -30.81123, -30.85891, -30.90615, -30.95305, 
        -30.99978, -31.04568, -31.09311, -31.14118, -31.19006, -31.23968, 
        -31.28979, -31.34006, -31.39011, -31.43962, -31.48833, -31.536, 
        -31.58237, -31.62748, -31.67162, -31.71541, -31.75848, -31.80335, 
        -31.84988, -31.89773, -31.94694, -31.99782, -32.0492, -32.10055, 
        -32.15144, -32.20207, -32.2527, -32.30378, -32.35565, -32.40817, 
        -32.46111, -32.51465, -32.56761, -32.62201, -32.67697, -32.73219, 
        -32.78735, -32.84238, -32.89713, -32.95158, -33.00554, -33.05879, 
        -33.1112, -33.16297, -33.21468, -33.26653, -33.31908, -33.37291, 
        -33.42648, -33.48204, -33.5375, -33.59254, -33.64685, -33.70043, 
        -33.75314, -33.80519, -33.85677, -33.90803, -33.95905, -34.00989, 
        -34.06077, -34.11171, -34.16267, -34.21339, -34.26358, -34.31208, 
        -34.3609, -34.40938, -34.45721, -34.50473, -34.55172, -34.59821, 
        -34.64367, -34.68748, -34.72941, -34.76959, -34.80863, -34.84711, 
        -34.88586, -34.92598, -34.96726, -35.00939, -35.05069, -35.09261, 
        -35.13385, -35.17437, -35.21416, -35.25317, -35.29132, -35.32861, 
        -35.36507, -35.40072, -35.43574, -35.47032, -35.50451, -35.53841, 
        -35.57193, -35.60495, -35.63742, -35.66935, -35.70085, -35.73093, 
        -35.76178, -35.79245, -35.82313, -35.85395, -35.88531, -35.91747, 
        -35.95034, -35.98351, -36.01654, -36.04914, -36.08124, -36.11288, 
        -36.14401, -36.17446, -36.20408, -36.23308, -36.26179, -36.29102, 
        -36.32087, -36.3503, -36.38103, -36.41183, -36.44247, -36.4728, 
        -36.50272, -36.53236, -36.56173, -36.59121, -36.621, -36.65119, 
        -36.68182, -36.71279, -36.7439, -36.77486, -36.80561, -36.83612, 
        -36.86639, -36.89648, -36.9263, -36.95569, -36.98445, -37.0111, 
        -37.03741, -37.06244, -37.08629, -37.10954, -37.13272, -37.1564, 
        -37.18095, -37.20642, -37.23277, -37.25983, -37.28711, -37.31403, 
        -37.34004, -37.36467, -37.38776, -37.40951, -37.43022, -37.45026, 
        -37.47015, -37.48996, -37.50965, -37.52922, -37.5487, -37.56725, 
        -37.58646, -37.60557, -37.62474, -37.6441, -37.66357, -37.68358, 
        -37.70417, -37.72502, -37.74594, -37.76647, -37.78621, -37.80492, 
        -37.82265, -37.83967, -37.85641, -37.87368, -37.89207, -37.91169, 
        -37.93261, -37.95446, -37.9767, -37.99932, -38.0224, -38.04606, 
        -38.0708, -38.09622, -38.12491, -38.15605, -38.18921, -38.22363, 
        -38.25866, -38.29329, -38.3269, -38.35971, -38.39119, -38.42149, 
        -38.45041, -38.47844, -38.5058, -38.53312, -38.56094, -38.58969, 
        -38.61975, -38.65112, -38.68359, -38.7165, -38.7492, -38.78119, 
        -38.81229, -38.84245, -38.87157, -38.89945, -38.92583, -38.95052, 
        -38.9735, -38.99469, -39.01351, -39.03264, -39.05173, -39.0708, 
        -39.08993, -39.10874, -39.12699, -39.14462, -39.16166, -39.17802, 
        -39.19333, -39.20742, -39.22029, -39.23223, -39.24339, -39.25372, 
        -39.26316, -39.27174, -39.2796, -39.28726, -39.29436, -39.30093, 
        -39.30666, -39.31128, -39.31488, -39.31769, -39.31997, -39.3216, 
        -39.32251, -39.32288, -39.32216, -39.3202, -39.31663, -39.31116, 
        -39.30374, -39.29442, -39.28325, -39.27037, -39.25496, -39.23912, 
        -39.22198, -39.20344, -39.18343, -39.16135, -39.13666, -39.10872, 
        -39.07745, -39.04325, -39.0072, -38.97051, -38.93392, -38.89754, 
        -38.86058, -38.82132, -38.77752, -38.72705, -38.66912, -38.60311, 
        -38.53061, -38.4545, -38.37897, -38.30911, -38.24963, -38.20487, 
        -38.17691,
  -30.3677, -30.41512, -30.46283, -30.51089, -30.55916, -30.60778, 
        -30.65672, -30.70561, -30.75421, -30.80116, -30.84836, -30.89502, 
        -30.94153, -30.98824, -31.03557, -31.08378, -31.13294, -31.18301, 
        -31.23382, -31.28489, -31.33584, -31.38596, -31.43507, -31.48169, 
        -31.528, -31.5731, -31.61741, -31.66161, -31.70635, -31.75223, 
        -31.79961, -31.84827, -31.89843, -31.94994, -32.00183, -32.05371, 
        -32.10519, -32.15637, -32.20757, -32.25792, -32.30991, -32.3623, 
        -32.4152, -32.46865, -32.52262, -32.57737, -32.63271, -32.68814, 
        -32.7435, -32.79854, -32.85325, -32.90757, -32.96146, -33.01468, 
        -33.06613, -33.11791, -33.16944, -33.22104, -33.27328, -33.32662, 
        -33.38074, -33.4352, -33.48994, -33.54417, -33.59768, -33.65044, 
        -33.70245, -33.75393, -33.80511, -33.85604, -33.90705, -33.95687, 
        -34.00785, -34.05904, -34.11016, -34.16072, -34.21043, -34.25921, 
        -34.30715, -34.35451, -34.40189, -34.44908, -34.49614, -34.54248, 
        -34.58764, -34.63116, -34.67266, -34.71232, -34.74981, -34.78791, 
        -34.82682, -34.86685, -34.90808, -34.95005, -34.99216, -35.03387, 
        -35.07501, -35.11552, -35.15522, -35.19416, -35.23226, -35.26948, 
        -35.30597, -35.34167, -35.37671, -35.41127, -35.44563, -35.47879, 
        -35.51269, -35.54608, -35.57882, -35.61097, -35.64262, -35.67398, 
        -35.70518, -35.73628, -35.76733, -35.79856, -35.83029, -35.8628, 
        -35.89608, -35.92943, -35.96255, -35.99495, -36.02684, -36.05836, 
        -36.08968, -36.11954, -36.14977, -36.17939, -36.20864, -36.2381, 
        -36.268, -36.29825, -36.32878, -36.3594, -36.3901, -36.42064, 
        -36.45081, -36.4809, -36.51081, -36.54095, -36.57153, -36.60247, 
        -36.63382, -36.66532, -36.69674, -36.72789, -36.75768, -36.78816, 
        -36.81844, -36.84857, -36.8785, -36.9079, -36.9365, -36.96385, 
        -36.98983, -37.01429, -37.03733, -37.05965, -37.08186, -37.10465, 
        -37.12832, -37.15311, -37.17887, -37.20561, -37.23283, -37.25999, 
        -37.28646, -37.31165, -37.33523, -37.35622, -37.37696, -37.39692, 
        -37.41651, -37.43604, -37.45559, -37.47518, -37.49493, -37.51448, 
        -37.53399, -37.55341, -37.57274, -37.59182, -37.61084, -37.63033, 
        -37.65007, -37.6699, -37.68968, -37.7091, -37.72784, -37.74577, 
        -37.76299, -37.77966, -37.79643, -37.81413, -37.83225, -37.85298, 
        -37.87506, -37.8983, -37.92206, -37.94637, -37.97099, -37.99627, 
        -38.02258, -38.05051, -38.08061, -38.11317, -38.14761, -38.18281, 
        -38.21846, -38.25362, -38.28778, -38.32073, -38.35235, -38.38273, 
        -38.41174, -38.43991, -38.46766, -38.4953, -38.52332, -38.55231, 
        -38.5825, -38.61388, -38.64628, -38.67914, -38.71086, -38.74299, 
        -38.77425, -38.80439, -38.83318, -38.86067, -38.88676, -38.91131, 
        -38.93459, -38.95617, -38.97687, -38.9962, -39.01532, -39.03405, 
        -39.05254, -39.07067, -39.08823, -39.10515, -39.12151, -39.13729, 
        -39.15218, -39.16603, -39.17881, -39.19075, -39.20203, -39.21265, 
        -39.22242, -39.23147, -39.23964, -39.24721, -39.25391, -39.26004, 
        -39.26528, -39.26951, -39.27286, -39.27458, -39.27666, -39.27809, 
        -39.27902, -39.27927, -39.27854, -39.27628, -39.27235, -39.26638, 
        -39.25841, -39.24858, -39.23694, -39.22379, -39.20929, -39.19359, 
        -39.17667, -39.15832, -39.13821, -39.11586, -39.09073, -39.06252, 
        -39.03112, -38.99704, -38.96125, -38.92467, -38.88812, -38.85168, 
        -38.81477, -38.77514, -38.7308, -38.67963, -38.61985, -38.55115, 
        -38.4752, -38.39495, -38.31525, -38.24204, -38.18031, -38.13494, 
        -38.10841,
  -30.30914, -30.35642, -30.40416, -30.45236, -30.49993, -30.54898, 
        -30.59842, -30.64807, -30.69732, -30.74583, -30.79338, -30.84011, 
        -30.88665, -30.93326, -30.98062, -31.02894, -31.07815, -31.1286, 
        -31.17999, -31.23084, -31.28259, -31.33325, -31.38255, -31.43039, 
        -31.47661, -31.52173, -31.56629, -31.61105, -31.65664, -31.70354, 
        -31.75201, -31.8017, -31.85269, -31.90457, -31.95617, -32.00844, 
        -32.06034, -32.11216, -32.16356, -32.21529, -32.26726, -32.31967, 
        -32.37247, -32.42581, -32.47988, -32.53452, -32.58974, -32.64518, 
        -32.70039, -32.75428, -32.8088, -32.86298, -32.91679, -32.97009, 
        -33.02271, -33.07465, -33.12619, -33.17778, -33.22984, -33.28261, 
        -33.33593, -33.3895, -33.44302, -33.49624, -33.54885, -33.60077, 
        -33.65108, -33.702, -33.75273, -33.80337, -33.85412, -33.90485, 
        -33.95601, -34.00707, -34.05802, -34.10837, -34.15761, -34.20569, 
        -34.2529, -34.29968, -34.34646, -34.39339, -34.44023, -34.4855, 
        -34.53067, -34.57409, -34.61539, -34.65485, -34.69318, -34.73131, 
        -34.77015, -34.81015, -34.85121, -34.89299, -34.935, -34.97667, 
        -35.01772, -35.05807, -35.09766, -35.13665, -35.17472, -35.21116, 
        -35.24784, -35.28382, -35.31907, -35.35378, -35.38819, -35.42244, 
        -35.45642, -35.48997, -35.52285, -35.55511, -35.58687, -35.61841, 
        -35.64986, -35.6813, -35.71271, -35.74434, -35.77649, -35.80945, 
        -35.84205, -35.87565, -35.90857, -35.9407, -35.97227, -36.00348, 
        -36.03471, -36.06581, -36.09642, -36.12652, -36.15628, -36.18605, 
        -36.21598, -36.24609, -36.27639, -36.30692, -36.33767, -36.36823, 
        -36.39891, -36.42955, -36.46011, -36.49015, -36.52156, -36.55337, 
        -36.58535, -36.61726, -36.64871, -36.67965, -36.71006, -36.7402, 
        -36.77026, -36.80029, -36.8302, -36.85966, -36.88822, -36.91548, 
        -36.94127, -36.96533, -36.98782, -37.00954, -37.03099, -37.05288, 
        -37.0758, -37.09883, -37.12406, -37.1504, -37.17745, -37.20469, 
        -37.23129, -37.25681, -37.28078, -37.30312, -37.32407, -37.34402, 
        -37.36348, -37.38282, -37.4023, -37.42197, -37.44169, -37.46159, 
        -37.48119, -37.50062, -37.51988, -37.53888, -37.5577, -37.57662, 
        -37.5956, -37.61449, -37.63212, -37.65036, -37.66811, -37.68531, 
        -37.70209, -37.71864, -37.73563, -37.75375, -37.7737, -37.79549, 
        -37.81871, -37.84313, -37.86834, -37.89404, -37.92037, -37.9473, 
        -37.97524, -38.0048, -38.03637, -38.07016, -38.10575, -38.14212, 
        -38.17843, -38.21417, -38.24883, -38.2822, -38.31389, -38.34431, 
        -38.37258, -38.40089, -38.42894, -38.45702, -38.48537, -38.51463, 
        -38.54505, -38.57645, -38.60879, -38.64157, -38.67413, -38.70621, 
        -38.73736, -38.76738, -38.79602, -38.82336, -38.84931, -38.87401, 
        -38.89761, -38.92015, -38.94095, -38.96078, -38.97936, -38.99775, 
        -39.01565, -39.03323, -39.05028, -39.06682, -39.0828, -39.09821, 
        -39.11287, -39.12659, -39.1393, -39.15023, -39.16151, -39.17218, 
        -39.18218, -39.19133, -39.19949, -39.20667, -39.21296, -39.21842, 
        -39.22315, -39.22693, -39.22998, -39.23244, -39.23444, -39.23591, 
        -39.23689, -39.23716, -39.23641, -39.23406, -39.22974, -39.22338, 
        -39.21494, -39.20465, -39.19273, -39.17947, -39.16498, -39.14941, 
        -39.13266, -39.11446, -39.09444, -39.07206, -39.04696, -39.0188, 
        -38.98763, -38.95397, -38.9187, -38.88263, -38.84639, -38.81001, 
        -38.77283, -38.73283, -38.68697, -38.63433, -38.57203, -38.50005, 
        -38.41983, -38.33495, -38.25071, -38.1732, -38.10891, -38.06298, 
        -38.03777,
  -30.25071, -30.2979, -30.34571, -30.39402, -30.44284, -30.4923, 
        -30.54235, -30.59253, -30.64247, -30.69157, -30.73967, -30.78695, 
        -30.83386, -30.88071, -30.92737, -30.9758, -31.02533, -31.07599, 
        -31.12769, -31.18009, -31.23224, -31.28333, -31.33294, -31.3809, 
        -31.42727, -31.47255, -31.51748, -31.56284, -31.60941, -31.65649, 
        -31.70609, -31.75691, -31.80863, -31.86107, -31.91382, -31.96651, 
        -32.01892, -32.07098, -32.1227, -32.17467, -32.22681, -32.27929, 
        -32.33214, -32.38538, -32.43819, -32.49257, -32.54737, -32.60223, 
        -32.65706, -32.71154, -32.76587, -32.81996, -32.87381, -32.92725, 
        -32.98013, -33.03231, -33.08406, -33.13562, -33.1875, -33.23971, 
        -33.29123, -33.34357, -33.39586, -33.44786, -33.49942, -33.55042, 
        -33.60101, -33.65139, -33.7017, -33.75205, -33.80261, -33.85324, 
        -33.90405, -33.95505, -34.00586, -34.05585, -34.10468, -34.15131, 
        -34.19793, -34.24418, -34.2906, -34.33733, -34.38412, -34.43048, 
        -34.47571, -34.51915, -34.5605, -34.60002, -34.63842, -34.67657, 
        -34.71541, -34.7552, -34.79623, -34.83791, -34.87985, -34.92062, 
        -34.96169, -35.00188, -35.04128, -35.08003, -35.11825, -35.15599, 
        -35.19311, -35.22945, -35.26505, -35.29996, -35.3345, -35.36877, 
        -35.40271, -35.43623, -35.46914, -35.50146, -35.53325, -35.56483, 
        -35.59537, -35.62708, -35.65885, -35.69075, -35.72338, -35.75669, 
        -35.79055, -35.8242, -35.857, -35.88878, -35.91979, -35.95062, 
        -35.98158, -36.01259, -36.04342, -36.07389, -36.10403, -36.13409, 
        -36.16417, -36.19432, -36.22369, -36.25415, -36.28476, -36.31575, 
        -36.34674, -36.37792, -36.40905, -36.44093, -36.47321, -36.50585, 
        -36.53838, -36.57037, -36.60156, -36.63196, -36.6617, -36.6912, 
        -36.72073, -36.75047, -36.78025, -36.80975, -36.83851, -36.86585, 
        -36.89065, -36.91476, -36.93715, -36.95834, -36.9793, -37.00055, 
        -37.02264, -37.04606, -37.07071, -37.09663, -37.12346, -37.15055, 
        -37.1772, -37.20279, -37.22692, -37.24949, -37.27061, -37.2906, 
        -37.30997, -37.32916, -37.34861, -37.36831, -37.38817, -37.40806, 
        -37.42675, -37.44615, -37.46531, -37.48433, -37.50304, -37.52161, 
        -37.53999, -37.55798, -37.57553, -37.59273, -37.60955, -37.62617, 
        -37.64268, -37.65936, -37.67677, -37.69561, -37.7164, -37.73911, 
        -37.76335, -37.78883, -37.8152, -37.8421, -37.86976, -37.8982, 
        -37.9278, -37.95897, -37.99099, -38.02599, -38.06242, -38.09954, 
        -38.13685, -38.17325, -38.2086, -38.24247, -38.2747, -38.30541, 
        -38.33484, -38.36347, -38.39181, -38.4203, -38.44928, -38.4789, 
        -38.50948, -38.54098, -38.57318, -38.60578, -38.63818, -38.6701, 
        -38.70112, -38.73096, -38.75946, -38.78668, -38.81268, -38.83768, 
        -38.8618, -38.88475, -38.906, -38.92463, -38.94287, -38.96084, 
        -38.97837, -38.99561, -39.01244, -39.02877, -39.04457, -39.05976, 
        -39.07424, -39.08781, -39.10048, -39.11226, -39.12346, -39.13415, 
        -39.14415, -39.15328, -39.16123, -39.16805, -39.17376, -39.17868, 
        -39.18279, -39.18605, -39.18867, -39.19077, -39.19257, -39.19407, 
        -39.19518, -39.19554, -39.19483, -39.19249, -39.18808, -39.18133, 
        -39.17241, -39.16175, -39.14964, -39.13628, -39.12191, -39.10549, 
        -39.08891, -39.07091, -39.05117, -39.02912, -39.00438, -38.97663, 
        -38.94601, -38.91308, -38.8785, -38.84308, -38.80729, -38.77095, 
        -38.7334, -38.69284, -38.64668, -38.59193, -38.52689, -38.45115, 
        -38.36627, -38.27679, -38.18786, -38.10612, -38.03913, -37.99255, 
        -37.96877,
  -30.19505, -30.24205, -30.28983, -30.33828, -30.38739, -30.4372, 
        -30.4876, -30.53822, -30.58855, -30.63716, -30.68588, -30.73393, 
        -30.78161, -30.82936, -30.87749, -30.92629, -30.97607, -31.02701, 
        -31.07902, -31.1316, -31.18394, -31.23528, -31.2851, -31.33324, 
        -31.37888, -31.42459, -31.47011, -31.51623, -31.5638, -31.61298, 
        -31.66362, -31.71532, -31.76773, -31.82055, -31.87355, -31.92646, 
        -31.97906, -32.03133, -32.08345, -32.13468, -32.18712, -32.2398, 
        -32.29274, -32.34591, -32.3994, -32.45327, -32.50737, -32.56153, 
        -32.61564, -32.66965, -32.72364, -32.77759, -32.83153, -32.88516, 
        -32.93827, -32.98964, -33.04164, -33.09332, -33.14499, -33.19667, 
        -33.24818, -33.29936, -33.35024, -33.40086, -33.45127, -33.5014, 
        -33.55133, -33.60122, -33.65117, -33.70124, -33.75155, -33.8021, 
        -33.85185, -33.90264, -33.95309, -34.00271, -34.05114, -34.09838, 
        -34.14476, -34.19086, -34.23713, -34.28376, -34.33059, -34.37701, 
        -34.42231, -34.46583, -34.50732, -34.54704, -34.58565, -34.62299, 
        -34.66179, -34.70152, -34.74234, -34.78408, -34.82624, -34.86819, 
        -34.90929, -34.9493, -34.98836, -35.02692, -35.06523, -35.10328, 
        -35.14083, -35.1776, -35.21357, -35.24877, -35.28348, -35.31774, 
        -35.35064, -35.38414, -35.41709, -35.44942, -35.48122, -35.51276, 
        -35.54433, -35.57609, -35.6081, -35.64048, -35.67341, -35.70698, 
        -35.74083, -35.77429, -35.80678, -35.83813, -35.86872, -35.89917, 
        -35.92978, -35.95958, -35.99037, -36.02098, -36.05144, -36.08179, 
        -36.11209, -36.14238, -36.17276, -36.20334, -36.23421, -36.26549, 
        -36.29688, -36.32843, -36.36043, -36.39289, -36.42575, -36.45877, 
        -36.49146, -36.52331, -36.55407, -36.58378, -36.61272, -36.64045, 
        -36.66929, -36.6985, -36.728, -36.75743, -36.78636, -36.81404, 
        -36.84023, -36.86465, -36.88722, -36.9084, -36.92902, -36.94978, 
        -36.97131, -36.99412, -37.0182, -37.04371, -37.07023, -37.09706, 
        -37.12356, -37.14902, -37.17313, -37.19576, -37.21593, -37.23587, 
        -37.25508, -37.27407, -37.29337, -37.31312, -37.33294, -37.35277, 
        -37.37247, -37.39174, -37.4109, -37.42997, -37.44882, -37.46735, 
        -37.48534, -37.50266, -37.51936, -37.53563, -37.55169, -37.5678, 
        -37.58414, -37.60102, -37.61902, -37.63871, -37.66044, -37.68406, 
        -37.7083, -37.73456, -37.76168, -37.78952, -37.81825, -37.84806, 
        -37.8792, -37.91196, -37.94637, -37.98244, -38.01976, -38.05775, 
        -38.09581, -38.13326, -38.16936, -38.20384, -38.23656, -38.26759, 
        -38.29734, -38.32636, -38.35525, -38.3842, -38.4137, -38.44392, 
        -38.47483, -38.50652, -38.53873, -38.57117, -38.60339, -38.63406, 
        -38.66481, -38.69439, -38.72272, -38.74988, -38.77605, -38.80135, 
        -38.82565, -38.84852, -38.86988, -38.88943, -38.9077, -38.92532, 
        -38.94265, -38.95977, -38.97655, -38.99281, -39.00846, -39.02349, 
        -39.03775, -39.05114, -39.06364, -39.07531, -39.08635, -39.09689, 
        -39.10683, -39.11583, -39.1237, -39.13021, -39.13547, -39.13997, 
        -39.14355, -39.14631, -39.14837, -39.15002, -39.15048, -39.15188, 
        -39.153, -39.15349, -39.15291, -39.15062, -39.14608, -39.13906, 
        -39.12976, -39.11869, -39.10629, -39.09285, -39.07856, -39.06338, 
        -39.04712, -39.02956, -39.01031, -38.9889, -38.96483, -38.93782, 
        -38.90799, -38.87588, -38.84215, -38.80738, -38.77191, -38.73558, 
        -38.69747, -38.65588, -38.60792, -38.55083, -38.48267, -38.40324, 
        -38.3143, -38.21994, -38.12643, -38.04136, -37.97204, -37.92453, 
        -37.90193,
  -30.14174, -30.18853, -30.23619, -30.28469, -30.33398, -30.38298, 
        -30.43354, -30.48432, -30.53488, -30.5849, -30.63409, -30.68283, 
        -30.73149, -30.78025, -30.8292, -30.87867, -30.92896, -30.9803, 
        -31.03251, -31.08423, -31.13663, -31.18802, -31.238, -31.28642, 
        -31.33344, -31.37981, -31.42602, -31.47304, -31.52165, -31.57174, 
        -31.62321, -31.67554, -31.72833, -31.78129, -31.8334, -31.88645, 
        -31.93912, -31.99162, -32.04409, -32.09673, -32.14959, -32.20264, 
        -32.2558, -32.30896, -32.36207, -32.41539, -32.46869, -32.52197, 
        -32.57531, -32.6287, -32.68122, -32.73487, -32.78866, -32.84228, 
        -32.89549, -32.94821, -33.00034, -33.05197, -33.10339, -33.15447, 
        -33.20504, -33.2551, -33.30465, -33.35394, -33.40325, -33.45253, 
        -33.50087, -33.5504, -33.60017, -33.65018, -33.70047, -33.751, 
        -33.80168, -33.85224, -33.90238, -33.95192, -33.99997, -34.04699, 
        -34.09335, -34.1395, -34.18575, -34.23228, -34.27918, -34.32557, 
        -34.36977, -34.41338, -34.45501, -34.49499, -34.53382, -34.57234, 
        -34.61118, -34.65097, -34.69188, -34.73382, -34.7762, -34.81832, 
        -34.8595, -34.89948, -34.93828, -34.97668, -35.01499, -35.05316, 
        -35.08999, -35.1271, -35.16338, -35.19888, -35.23373, -35.26805, 
        -35.30193, -35.33544, -35.36842, -35.40079, -35.43269, -35.46439, 
        -35.49606, -35.52803, -35.56028, -35.59286, -35.62596, -35.65946, 
        -35.69301, -35.72509, -35.75708, -35.78796, -35.81823, -35.84835, 
        -35.87862, -35.90919, -35.93983, -35.97046, -36.00109, -36.03172, 
        -36.06232, -36.0929, -36.12347, -36.15422, -36.18528, -36.21672, 
        -36.2485, -36.28063, -36.31316, -36.34596, -36.37801, -36.41093, 
        -36.44336, -36.47486, -36.50507, -36.53423, -36.56254, -36.59052, 
        -36.61861, -36.64715, -36.67614, -36.70534, -36.73424, -36.76242, 
        -36.78916, -36.81411, -36.83718, -36.8587, -36.87937, -36.89991, 
        -36.92094, -36.94318, -36.96577, -36.99081, -37.01684, -37.0433, 
        -37.06946, -37.09464, -37.11864, -37.14118, -37.16224, -37.18209, 
        -37.20109, -37.21985, -37.23898, -37.25851, -37.27816, -37.29787, 
        -37.31755, -37.33692, -37.35621, -37.37544, -37.39442, -37.41307, 
        -37.43089, -37.44774, -37.46381, -37.47835, -37.49373, -37.50935, 
        -37.52572, -37.54276, -37.5613, -37.58194, -37.60466, -37.62919, 
        -37.65509, -37.68194, -37.70959, -37.73817, -37.76788, -37.79906, 
        -37.83167, -37.86586, -37.90173, -37.93893, -37.97708, -38.01589, 
        -38.05486, -38.09301, -38.12996, -38.16516, -38.19843, -38.23, 
        -38.26026, -38.28884, -38.31831, -38.34798, -38.37799, -38.40873, 
        -38.44012, -38.47207, -38.50432, -38.53658, -38.56868, -38.60007, 
        -38.63052, -38.6598, -38.68791, -38.71493, -38.74105, -38.76633, 
        -38.79056, -38.81341, -38.83458, -38.85411, -38.87235, -38.89009, 
        -38.90746, -38.92466, -38.94144, -38.9576, -38.97313, -38.98783, 
        -39.00178, -39.01511, -39.02735, -39.03877, -39.04858, -39.05889, 
        -39.06864, -39.07754, -39.08528, -39.09168, -39.09674, -39.101, 
        -39.10426, -39.10661, -39.10831, -39.10956, -39.11063, -39.11169, 
        -39.11273, -39.11312, -39.11253, -39.11019, -39.10558, -39.09837, 
        -39.08876, -39.0774, -39.06481, -39.05112, -39.03682, -39.02206, 
        -39.00618, -38.98918, -38.9707, -38.95014, -38.92695, -38.90088, 
        -38.87195, -38.84075, -38.80784, -38.77362, -38.7384, -38.70182, 
        -38.66294, -38.61996, -38.56995, -38.51027, -38.43808, -38.35521, 
        -38.26251, -38.16424, -38.06702, -37.97906, -37.90816, -37.86021, 
        -37.83838,
  -30.0902, -30.13681, -30.18427, -30.23269, -30.28192, -30.33187, 
        -30.38237, -30.43307, -30.48361, -30.53374, -30.58345, -30.63301, 
        -30.68263, -30.73234, -30.78228, -30.83154, -30.88252, -30.93434, 
        -30.98682, -31.03962, -31.0921, -31.14357, -31.1937, -31.24241, 
        -31.29001, -31.33688, -31.38396, -31.43202, -31.48127, -31.53097, 
        -31.58318, -31.63589, -31.68876, -31.74184, -31.79494, -31.84805, 
        -31.90085, -31.95357, -32.00637, -32.05943, -32.11277, -32.16623, 
        -32.21965, -32.27282, -32.32573, -32.37717, -32.42968, -32.48222, 
        -32.53482, -32.58762, -32.64053, -32.69364, -32.74701, -32.8004, 
        -32.85357, -32.90639, -32.95866, -33.01037, -33.06147, -33.11193, 
        -33.16159, -33.20945, -33.25784, -33.30601, -33.35431, -33.40287, 
        -33.45181, -33.50116, -33.5509, -33.60098, -33.65142, -33.70199, 
        -33.75264, -33.80308, -33.85302, -33.90189, -33.95, -33.99689, 
        -34.04238, -34.08906, -34.13551, -34.18204, -34.22881, -34.27502, 
        -34.32041, -34.36392, -34.40575, -34.44601, -34.48519, -34.52405, 
        -34.56323, -34.60321, -34.64423, -34.68628, -34.72884, -34.77113, 
        -34.81136, -34.85128, -34.89003, -34.92817, -34.96634, -35.00456, 
        -35.04247, -35.07981, -35.11639, -35.15213, -35.18716, -35.22158, 
        -35.25552, -35.28902, -35.32201, -35.35454, -35.38665, -35.41861, 
        -35.4506, -35.48175, -35.51429, -35.547, -35.57991, -35.61304, 
        -35.64607, -35.67855, -35.70997, -35.74038, -35.77036, -35.80019, 
        -35.83025, -35.86047, -35.89089, -35.92145, -35.95222, -35.9831, 
        -36.01404, -36.04497, -36.07575, -36.10571, -36.13696, -36.16857, 
        -36.20056, -36.23293, -36.26564, -36.29851, -36.33138, -36.36397, 
        -36.39594, -36.42686, -36.45665, -36.48551, -36.5134, -36.54085, 
        -36.56835, -36.59613, -36.62448, -36.65322, -36.68201, -36.71034, 
        -36.73761, -36.76223, -36.786, -36.80809, -36.82907, -36.84965, 
        -36.87053, -36.8923, -36.91542, -36.93986, -36.96531, -36.99118, 
        -37.01679, -37.04164, -37.06525, -37.08756, -37.10849, -37.12824, 
        -37.14695, -37.16551, -37.18436, -37.20356, -37.22327, -37.24286, 
        -37.26234, -37.28077, -37.30027, -37.31977, -37.33904, -37.35767, 
        -37.37538, -37.39202, -37.40769, -37.4227, -37.43758, -37.45285, 
        -37.46897, -37.48615, -37.50545, -37.52711, -37.55058, -37.57585, 
        -37.60236, -37.6296, -37.6577, -37.68709, -37.71783, -37.75024, 
        -37.78443, -37.82019, -37.85737, -37.8957, -37.93388, -37.97347, 
        -38.01311, -38.05204, -38.08967, -38.1256, -38.15953, -38.19181, 
        -38.22266, -38.25294, -38.28307, -38.3134, -38.34415, -38.37542, 
        -38.40721, -38.43944, -38.47175, -38.50385, -38.53585, -38.56693, 
        -38.59704, -38.62596, -38.6538, -38.68063, -38.70657, -38.73159, 
        -38.75557, -38.77835, -38.79953, -38.81903, -38.83735, -38.85433, 
        -38.87193, -38.88921, -38.90598, -38.92198, -38.93716, -38.95141, 
        -38.96524, -38.9781, -38.99018, -39.00135, -39.0118, -39.02178, 
        -39.03121, -39.03988, -39.04752, -39.0539, -39.05915, -39.06323, 
        -39.06645, -39.06879, -39.07039, -39.07145, -39.07225, -39.073, 
        -39.07352, -39.07371, -39.07289, -39.07036, -39.06568, -39.05838, 
        -39.04858, -39.03687, -39.0239, -39.01017, -38.99605, -38.98132, 
        -38.96592, -38.94866, -38.931, -38.91135, -38.88906, -38.86398, 
        -38.83604, -38.80564, -38.77349, -38.73985, -38.70467, -38.66767, 
        -38.62785, -38.58318, -38.53127, -38.46912, -38.39536, -38.30946, 
        -38.21355, -38.11242, -38.01288, -37.92302, -37.85092, -37.80285, 
        -37.78149,
  -30.04291, -30.08923, -30.13641, -30.1845, -30.23346, -30.28317, 
        -30.33348, -30.38398, -30.4344, -30.48455, -30.53353, -30.58362, 
        -30.63382, -30.6844, -30.7354, -30.7865, -30.83822, -30.89056, 
        -30.94337, -30.9963, -31.04884, -31.10047, -31.15089, -31.20007, 
        -31.24827, -31.29495, -31.34283, -31.3915, -31.44134, -31.49244, 
        -31.54459, -31.59738, -31.65042, -31.70349, -31.7565, -31.80942, 
        -31.86231, -31.91535, -31.96868, -32.02237, -32.07537, -32.12938, 
        -32.18304, -32.23609, -32.28848, -32.34041, -32.39217, -32.44397, 
        -32.49589, -32.54813, -32.6005, -32.65295, -32.70563, -32.75846, 
        -32.81139, -32.86419, -32.91557, -32.96726, -33.01807, -33.06786, 
        -33.1166, -33.16451, -33.2119, -33.25918, -33.30667, -33.35468, 
        -33.40337, -33.45275, -33.50267, -33.55292, -33.6035, -33.65414, 
        -33.70374, -33.75404, -33.80375, -33.85262, -33.90068, -33.94771, 
        -33.99441, -34.04118, -34.08774, -34.13457, -34.18137, -34.22771, 
        -34.27274, -34.3164, -34.35851, -34.39925, -34.43898, -34.47836, 
        -34.51691, -34.55713, -34.59832, -34.64044, -34.68296, -34.72524, 
        -34.76642, -34.80632, -34.84503, -34.88324, -34.92137, -34.95951, 
        -34.9974, -35.03485, -35.07155, -35.1075, -35.14273, -35.17731, 
        -35.21129, -35.2438, -35.27683, -35.30951, -35.3419, -35.37426, 
        -35.40668, -35.43921, -35.47178, -35.5043, -35.5369, -35.56961, 
        -35.60196, -35.63366, -35.66445, -35.69453, -35.72424, -35.75389, 
        -35.78361, -35.81342, -35.84247, -35.87289, -35.90378, -35.93499, 
        -35.96635, -35.99759, -36.0286, -36.05975, -36.09095, -36.12243, 
        -36.15442, -36.1868, -36.21944, -36.25211, -36.28456, -36.31657, 
        -36.34794, -36.37849, -36.4081, -36.4368, -36.46466, -36.49193, 
        -36.51798, -36.54516, -36.57277, -36.60088, -36.62925, -36.65753, 
        -36.68513, -36.71132, -36.73578, -36.7586, -36.78006, -36.80087, 
        -36.82174, -36.84328, -36.86591, -36.88969, -36.91438, -36.93948, 
        -36.96444, -36.98877, -37.01207, -37.03412, -37.05478, -37.07318, 
        -37.09174, -37.11004, -37.12859, -37.14764, -37.16684, -37.1862, 
        -37.20561, -37.22511, -37.24478, -37.26458, -37.28402, -37.30272, 
        -37.32049, -37.33707, -37.35252, -37.3672, -37.3817, -37.39668, 
        -37.41273, -37.43044, -37.45037, -37.47242, -37.49661, -37.52251, 
        -37.54931, -37.57608, -37.60486, -37.63504, -37.66697, -37.70086, 
        -37.73666, -37.77409, -37.81276, -37.8523, -37.89244, -37.93295, 
        -37.97321, -38.01288, -38.05113, -38.08756, -38.12217, -38.15516, 
        -38.18695, -38.21796, -38.24872, -38.27965, -38.31097, -38.34277, 
        -38.37495, -38.40734, -38.4397, -38.47178, -38.50354, -38.53438, 
        -38.56301, -38.59164, -38.61905, -38.64547, -38.67113, -38.6958, 
        -38.71965, -38.74256, -38.76336, -38.78305, -38.80193, -38.82007, 
        -38.83795, -38.85538, -38.87202, -38.88768, -38.9024, -38.91632, 
        -38.9296, -38.94219, -38.95386, -38.9647, -38.97482, -38.98441, 
        -38.99353, -39.00204, -39.0097, -39.01627, -39.0217, -39.02601, 
        -39.02937, -39.03187, -39.03362, -39.03474, -39.03543, -39.03582, 
        -39.03487, -39.03443, -39.0331, -39.03034, -39.02552, -39.0182, 
        -39.00836, -38.99651, -38.98332, -38.9694, -38.9551, -38.94054, 
        -38.92563, -38.91, -38.8931, -38.87418, -38.8527, -38.82846, 
        -38.80138, -38.77194, -38.74063, -38.70729, -38.6722, -38.63474, 
        -38.59383, -38.54767, -38.49378, -38.42943, -38.35339, -38.26521, 
        -38.16709, -38.06405, -37.96304, -37.87236, -37.80008, -37.75216, 
        -37.73102,
  -29.99861, -30.0447, -30.0916, -30.13927, -30.18779, -30.23613, 
        -30.28608, -30.33627, -30.38655, -30.43669, -30.48682, -30.53715, 
        -30.58797, -30.6393, -30.69104, -30.74309, -30.79553, -30.84825, 
        -30.90131, -30.95437, -31.0061, -31.05787, -31.10857, -31.15832, 
        -31.20718, -31.25564, -31.30423, -31.3535, -31.40374, -31.45506, 
        -31.50723, -31.55996, -31.6129, -31.66573, -31.71875, -31.77063, 
        -31.82355, -31.87694, -31.93066, -31.98478, -32.03914, -32.0934, 
        -32.1471, -32.19994, -32.25181, -32.30318, -32.35445, -32.40578, 
        -32.45739, -32.50909, -32.56095, -32.61183, -32.66375, -32.71598, 
        -32.76854, -32.821, -32.87322, -32.92465, -32.97506, -33.02428, 
        -33.07232, -33.11945, -33.16622, -33.21287, -33.25979, -33.3074, 
        -33.35587, -33.40423, -33.45429, -33.5048, -33.55545, -33.60624, 
        -33.65695, -33.70734, -33.75714, -33.80607, -33.85406, -33.90148, 
        -33.94845, -33.99533, -34.04216, -34.08922, -34.13617, -34.18228, 
        -34.22641, -34.27014, -34.31241, -34.35358, -34.39356, -34.43346, 
        -34.47345, -34.51403, -34.55553, -34.59779, -34.64022, -34.6823, 
        -34.72333, -34.76311, -34.80199, -34.84037, -34.87851, -34.91668, 
        -34.95364, -34.991, -35.02782, -35.06401, -35.0995, -35.13422, 
        -35.16835, -35.2019, -35.23497, -35.26774, -35.30031, -35.33289, 
        -35.36554, -35.39832, -35.43079, -35.46315, -35.49538, -35.52749, 
        -35.55919, -35.59026, -35.61959, -35.64926, -35.67858, -35.70789, 
        -35.73725, -35.76671, -35.79644, -35.82672, -35.85763, -35.88905, 
        -35.9206, -35.95213, -35.98331, -36.01448, -36.04549, -36.0768, 
        -36.1086, -36.14071, -36.1731, -36.20549, -36.23758, -36.26817, 
        -36.2992, -36.32948, -36.35899, -36.38786, -36.41578, -36.44297, 
        -36.46975, -36.49644, -36.52339, -36.55084, -36.57857, -36.60647, 
        -36.63391, -36.66037, -36.68534, -36.70875, -36.73086, -36.75214, 
        -36.77325, -36.79471, -36.81689, -36.8389, -36.86266, -36.8868, 
        -36.91094, -36.93457, -36.95738, -36.9791, -36.9995, -37.01865, 
        -37.03712, -37.05529, -37.07378, -37.09262, -37.1118, -37.13116, 
        -37.15061, -37.17012, -37.18972, -37.2093, -37.22856, -37.24722, 
        -37.26485, -37.28133, -37.2967, -37.31131, -37.32481, -37.33994, 
        -37.35627, -37.37442, -37.39472, -37.41722, -37.44186, -37.46806, 
        -37.49537, -37.52371, -37.55325, -37.58457, -37.61783, -37.65327, 
        -37.69078, -37.72991, -37.77016, -37.81107, -37.85244, -37.89372, 
        -37.93463, -37.9744, -38.01301, -38.04976, -38.08506, -38.11873, 
        -38.15165, -38.18328, -38.21381, -38.24546, -38.27734, -38.30947, 
        -38.34187, -38.3743, -38.4066, -38.4387, -38.47012, -38.50066, 
        -38.52999, -38.55827, -38.58546, -38.61164, -38.63695, -38.66163, 
        -38.68526, -38.70804, -38.72911, -38.74913, -38.76818, -38.78676, 
        -38.80481, -38.82222, -38.8387, -38.85402, -38.86825, -38.88168, 
        -38.89441, -38.90634, -38.91753, -38.92784, -38.93748, -38.94558, 
        -38.9544, -38.96286, -38.97064, -38.97745, -38.98334, -38.98807, 
        -38.99191, -38.99488, -38.99703, -38.99842, -38.99916, -38.99929, 
        -38.99887, -38.99786, -38.99592, -38.99273, -38.98772, -38.98033, 
        -38.97052, -38.95865, -38.94538, -38.93126, -38.91681, -38.90225, 
        -38.88742, -38.87212, -38.8558, -38.83747, -38.81673, -38.7933, 
        -38.76727, -38.73861, -38.70797, -38.67502, -38.63974, -38.60146, 
        -38.55925, -38.51138, -38.4556, -38.3895, -38.31147, -38.22152, 
        -38.12098, -38.01716, -37.91587, -37.82528, -37.75369, -37.7062, 
        -37.68512,
  -29.95711, -30.00209, -30.04859, -30.09589, -30.14397, -30.19285, 
        -30.24244, -30.2924, -30.34219, -30.39224, -30.44239, -30.49289, 
        -30.54399, -30.59578, -30.64817, -30.69985, -30.75297, -30.80639, 
        -30.85957, -30.91265, -30.96541, -31.01721, -31.06844, -31.11885, 
        -31.16844, -31.2176, -31.26683, -31.3165, -31.3669, -31.41816, 
        -31.46914, -31.52162, -31.5744, -31.62722, -31.68011, -31.73296, 
        -31.78625, -31.83993, -31.89405, -31.94847, -32.00298, -32.05724, 
        -32.11072, -32.16316, -32.21462, -32.26561, -32.31561, -32.36685, 
        -32.41839, -32.46989, -32.52138, -32.57262, -32.62374, -32.67517, 
        -32.72696, -32.779, -32.83081, -32.88187, -32.93178, -32.98023, 
        -33.02777, -33.07449, -33.12, -33.16636, -33.21305, -33.26041, 
        -33.30873, -33.35805, -33.4082, -33.45884, -33.50971, -33.56063, 
        -33.61152, -33.66207, -33.71198, -33.76101, -33.80904, -33.85643, 
        -33.90362, -33.94975, -33.99697, -34.04441, -34.09142, -34.13771, 
        -34.18295, -34.22679, -34.26936, -34.3107, -34.35114, -34.39141, 
        -34.43184, -34.47279, -34.51455, -34.55698, -34.59927, -34.64094, 
        -34.68179, -34.72068, -34.75998, -34.7985, -34.83691, -34.8751, 
        -34.91316, -34.95058, -34.98747, -35.0237, -35.05933, -35.09431, 
        -35.12863, -35.16219, -35.19525, -35.22801, -35.26067, -35.29344, 
        -35.32618, -35.35893, -35.39029, -35.4223, -35.45396, -35.48535, 
        -35.51649, -35.54713, -35.57698, -35.60627, -35.63536, -35.6643, 
        -35.69329, -35.72233, -35.75171, -35.78176, -35.81257, -35.844, 
        -35.87567, -35.90728, -35.93856, -35.96956, -35.9994, -36.0303, 
        -36.06168, -36.09351, -36.12545, -36.15753, -36.18929, -36.22062, 
        -36.25147, -36.28184, -36.31161, -36.34069, -36.3689, -36.39629, 
        -36.42308, -36.44946, -36.47586, -36.50251, -36.52953, -36.55654, 
        -36.58345, -36.60971, -36.63382, -36.65771, -36.68048, -36.70235, 
        -36.72372, -36.74509, -36.76673, -36.78885, -36.81156, -36.83465, 
        -36.85792, -36.88091, -36.90329, -36.92464, -36.94484, -36.96392, 
        -36.98228, -37.00053, -37.01904, -37.03776, -37.05703, -37.07639, 
        -37.09593, -37.11535, -37.13369, -37.15282, -37.17162, -37.18989, 
        -37.20729, -37.22363, -37.23901, -37.2538, -37.26866, -37.28426, 
        -37.30111, -37.31965, -37.34027, -37.36298, -37.38776, -37.41422, 
        -37.44195, -37.47108, -37.50183, -37.53452, -37.56934, -37.60648, 
        -37.64597, -37.68695, -37.72901, -37.77145, -37.81379, -37.85508, 
        -37.89642, -37.93631, -37.97486, -38.01194, -38.04764, -38.08224, 
        -38.11565, -38.14849, -38.18068, -38.21287, -38.2452, -38.2777, 
        -38.31023, -38.34257, -38.37465, -38.40636, -38.43744, -38.46757, 
        -38.49677, -38.52479, -38.55172, -38.57775, -38.60286, -38.62729, 
        -38.65085, -38.67375, -38.69519, -38.71565, -38.73524, -38.7541, 
        -38.77135, -38.78878, -38.80504, -38.81998, -38.83367, -38.84639, 
        -38.85836, -38.86959, -38.88008, -38.88983, -38.89895, -38.9077, 
        -38.91642, -38.92496, -38.93295, -38.94037, -38.94674, -38.95202, 
        -38.95642, -38.95995, -38.96263, -38.9644, -38.96529, -38.96532, 
        -38.96439, -38.9627, -38.96001, -38.95638, -38.95103, -38.94371, 
        -38.93397, -38.92226, -38.90887, -38.89455, -38.87986, -38.86507, 
        -38.85019, -38.83505, -38.81895, -38.80015, -38.78014, -38.75756, 
        -38.73241, -38.70462, -38.67452, -38.64178, -38.60625, -38.56723, 
        -38.5237, -38.47408, -38.41644, -38.34844, -38.26863, -38.17723, 
        -38.07692, -37.97239, -37.87124, -37.78217, -37.71178, -37.66525, 
        -37.64421,
  -29.91714, -29.96315, -30.00936, -30.05625, -30.10387, -30.15224, 
        -30.20137, -30.25076, -30.30037, -30.35018, -30.40028, -30.44996, 
        -30.50128, -30.55345, -30.60647, -30.65992, -30.71356, -30.76721, 
        -30.82063, -30.87372, -30.92621, -30.97825, -31.02981, -31.08071, 
        -31.1309, -31.17967, -31.22941, -31.27945, -31.33001, -31.38125, 
        -31.43311, -31.48553, -31.53823, -31.59093, -31.64369, -31.69666, 
        -31.75009, -31.80401, -31.85819, -31.91251, -31.96674, -32.01959, 
        -32.07265, -32.12472, -32.17598, -32.22684, -32.27783, -32.32925, 
        -32.38093, -32.4325, -32.48368, -32.53439, -32.58484, -32.63541, 
        -32.68645, -32.73781, -32.78905, -32.83847, -32.88758, -32.9356, 
        -32.98267, -33.02924, -33.07578, -33.12223, -33.16898, -33.21629, 
        -33.26444, -33.31361, -33.36366, -33.41425, -33.46517, -33.51624, 
        -33.56734, -33.61716, -33.66738, -33.71652, -33.76469, -33.81213, 
        -33.85945, -33.90682, -33.95446, -34.00211, -34.04937, -34.09582, 
        -34.14114, -34.18521, -34.22791, -34.26944, -34.31041, -34.3509, 
        -34.3916, -34.43192, -34.47409, -34.51639, -34.55878, -34.60072, 
        -34.64162, -34.68145, -34.72091, -34.75969, -34.79826, -34.83659, 
        -34.87466, -34.91208, -34.94882, -34.98511, -35.02091, -35.05607, 
        -35.09049, -35.12313, -35.15624, -35.18904, -35.22173, -35.25444, 
        -35.2871, -35.3195, -35.3514, -35.38282, -35.41385, -35.44469, 
        -35.47538, -35.50564, -35.53511, -35.56405, -35.59277, -35.62141, 
        -35.65007, -35.67881, -35.70798, -35.73671, -35.76724, -35.7984, 
        -35.82985, -35.86129, -35.89245, -35.92327, -35.95384, -35.98436, 
        -36.0153, -36.04662, -36.07826, -36.10997, -36.14157, -36.1729, 
        -36.20388, -36.23453, -36.26473, -36.29426, -36.3229, -36.35067, 
        -36.37753, -36.4028, -36.42868, -36.45456, -36.48049, -36.50679, 
        -36.53273, -36.55851, -36.58351, -36.6076, -36.63079, -36.65309, 
        -36.67468, -36.69579, -36.71678, -36.73795, -36.75964, -36.78178, 
        -36.80428, -36.82673, -36.84865, -36.86972, -36.88971, -36.90876, 
        -36.92625, -36.94471, -36.96323, -36.98217, -37.00158, -37.02102, 
        -37.0404, -37.05994, -37.07869, -37.09716, -37.11534, -37.13295, 
        -37.14999, -37.16626, -37.18173, -37.19685, -37.21231, -37.22854, 
        -37.24596, -37.26508, -37.28601, -37.30886, -37.33372, -37.36038, 
        -37.38867, -37.41868, -37.44964, -37.48397, -37.52034, -37.55955, 
        -37.60094, -37.64373, -37.6873, -37.73127, -37.77498, -37.81796, 
        -37.85985, -37.89993, -37.93839, -37.97572, -38.01174, -38.04683, 
        -38.08109, -38.11464, -38.14758, -38.18052, -38.21323, -38.24598, 
        -38.27839, -38.31031, -38.34198, -38.37314, -38.40373, -38.43358, 
        -38.46256, -38.49062, -38.5167, -38.54277, -38.5679, -38.59224, 
        -38.61596, -38.6389, -38.66087, -38.68189, -38.70198, -38.72128, 
        -38.73978, -38.75718, -38.77311, -38.78758, -38.80061, -38.81253, 
        -38.82365, -38.83404, -38.84377, -38.85284, -38.86155, -38.87017, 
        -38.87874, -38.8872, -38.89573, -38.90367, -38.91077, -38.91685, 
        -38.92193, -38.92607, -38.92927, -38.93136, -38.93229, -38.93201, 
        -38.93073, -38.92749, -38.92419, -38.91985, -38.91424, -38.9069, 
        -38.89737, -38.88588, -38.87239, -38.85786, -38.84282, -38.82764, 
        -38.8126, -38.79741, -38.78154, -38.76434, -38.74516, -38.72354, 
        -38.69926, -38.67225, -38.64251, -38.60974, -38.57373, -38.5337, 
        -38.48872, -38.43745, -38.37793, -38.30815, -38.2267, -38.13371, 
        -38.03259, -37.92831, -37.8283, -37.74041, -37.67134, -37.62582, 
        -37.6048,
  -29.8809, -29.92661, -29.97261, -30.01895, -30.06601, -30.1138, 
        -30.16125, -30.21018, -30.25944, -30.30908, -30.35933, -30.41026, 
        -30.46201, -30.51478, -30.56832, -30.62236, -30.67653, -30.73043, 
        -30.78377, -30.83666, -30.88912, -30.94022, -30.99193, -31.04309, 
        -31.09371, -31.14396, -31.19415, -31.24453, -31.29535, -31.34655, 
        -31.3984, -31.45071, -31.50329, -31.55591, -31.60859, -31.66158, 
        -31.71405, -31.7679, -31.82197, -31.8758, -31.92944, -31.98276, 
        -32.03532, -32.08696, -32.13809, -32.18899, -32.24015, -32.29185, 
        -32.34371, -32.3954, -32.44649, -32.49587, -32.54592, -32.59586, 
        -32.64608, -32.69659, -32.74696, -32.79655, -32.84508, -32.89258, 
        -32.93943, -32.98621, -33.03296, -33.07977, -33.1268, -33.1741, 
        -33.22219, -33.27111, -33.31985, -33.37025, -33.42101, -33.47221, 
        -33.52351, -33.57463, -33.62508, -33.67453, -33.72287, -33.77054, 
        -33.81805, -33.86571, -33.91367, -33.96154, -34.00899, -34.05544, 
        -34.10084, -34.14368, -34.18644, -34.22829, -34.26957, -34.31047, 
        -34.35158, -34.39325, -34.43569, -34.47837, -34.52108, -34.56316, 
        -34.60438, -34.64443, -34.68387, -34.72276, -34.7613, -34.79961, 
        -34.83757, -34.87401, -34.91085, -34.94719, -34.98301, -35.0182, 
        -35.05264, -35.08633, -35.11941, -35.15229, -35.18505, -35.21762, 
        -35.24992, -35.28181, -35.31306, -35.34366, -35.37416, -35.40448, 
        -35.43471, -35.4645, -35.49368, -35.52126, -35.54963, -35.57796, 
        -35.60634, -35.63484, -35.66368, -35.69309, -35.7232, -35.75379, 
        -35.78471, -35.81583, -35.84679, -35.8773, -35.9075, -35.9376, 
        -35.9681, -35.99902, -36.03035, -36.06187, -36.09351, -36.12492, 
        -36.15511, -36.18623, -36.21695, -36.24691, -36.27612, -36.30423, 
        -36.33126, -36.35741, -36.38295, -36.40821, -36.43333, -36.45854, 
        -36.48375, -36.50885, -36.5335, -36.55751, -36.58086, -36.6033, 
        -36.62485, -36.64562, -36.66594, -36.68623, -36.70577, -36.72718, 
        -36.74901, -36.77088, -36.79263, -36.81347, -36.83339, -36.85249, 
        -36.87112, -36.88973, -36.90848, -36.92765, -36.9472, -36.967, 
        -36.98639, -37.00558, -37.02393, -37.04152, -37.05892, -37.07606, 
        -37.09266, -37.10878, -37.12435, -37.13985, -37.15586, -37.17182, 
        -37.19003, -37.20972, -37.23105, -37.25415, -37.2792, -37.30605, 
        -37.33489, -37.36578, -37.3991, -37.43471, -37.47319, -37.51395, 
        -37.557, -37.60158, -37.64703, -37.69249, -37.73748, -37.78128, 
        -37.82341, -37.86377, -37.90244, -37.93961, -37.97584, -38.01146, 
        -38.04637, -38.08067, -38.11448, -38.14799, -38.18014, -38.21297, 
        -38.24516, -38.27675, -38.30779, -38.33827, -38.36821, -38.39759, 
        -38.42636, -38.45459, -38.48195, -38.50838, -38.53378, -38.55829, 
        -38.58202, -38.60516, -38.62754, -38.64925, -38.67002, -38.68983, 
        -38.70873, -38.72586, -38.74147, -38.75549, -38.76777, -38.77882, 
        -38.78915, -38.79867, -38.80767, -38.81632, -38.82474, -38.83307, 
        -38.84146, -38.84931, -38.85828, -38.86671, -38.87444, -38.88123, 
        -38.88705, -38.89181, -38.89539, -38.89759, -38.8984, -38.8978, 
        -38.89607, -38.89305, -38.88904, -38.88424, -38.87846, -38.87134, 
        -38.86218, -38.85089, -38.83768, -38.82286, -38.80742, -38.79185, 
        -38.77658, -38.76137, -38.74578, -38.72919, -38.71093, -38.69029, 
        -38.66685, -38.64043, -38.61084, -38.57775, -38.54107, -38.50012, 
        -38.45373, -38.40087, -38.33941, -38.26761, -38.18449, -38.0903, 
        -37.98828, -37.884, -37.78339, -37.69674, -37.62928, -37.58431, 
        -37.56296,
  -29.84662, -29.89199, -29.93657, -29.98253, -30.02904, -30.07618, 
        -30.12401, -30.17243, -30.22138, -30.27095, -30.32134, -30.37275, 
        -30.42517, -30.47849, -30.5327, -30.58728, -30.64083, -30.69487, 
        -30.74809, -30.80074, -30.85304, -30.9051, -30.95688, -31.00824, 
        -31.05919, -31.10986, -31.1605, -31.21121, -31.26212, -31.31342, 
        -31.36518, -31.41651, -31.46898, -31.52146, -31.57392, -31.62674, 
        -31.68018, -31.73367, -31.78723, -31.84048, -31.8934, -31.94581, 
        -31.99778, -32.04901, -32.10009, -32.15116, -32.20173, -32.25368, 
        -32.30566, -32.35741, -32.40847, -32.45874, -32.50848, -32.55801, 
        -32.6075, -32.65722, -32.70657, -32.75521, -32.80304, -32.85029, 
        -32.89728, -32.94444, -32.99075, -33.03809, -33.08556, -33.13298, 
        -33.18087, -33.22942, -33.27874, -33.32878, -33.37935, -33.43055, 
        -33.48203, -33.53348, -33.58434, -33.63415, -33.68291, -33.73087, 
        -33.77858, -33.82565, -33.87384, -33.92177, -33.96917, -34.01569, 
        -34.06101, -34.10478, -34.14751, -34.18941, -34.23088, -34.27221, 
        -34.31367, -34.35555, -34.39819, -34.44148, -34.4846, -34.52718, 
        -34.56875, -34.60818, -34.64765, -34.68647, -34.72491, -34.76306, 
        -34.80089, -34.83833, -34.87531, -34.91163, -34.9474, -34.98238, 
        -35.01675, -35.05032, -35.08354, -35.11657, -35.14928, -35.18167, 
        -35.2135, -35.24473, -35.27424, -35.30425, -35.33415, -35.36395, 
        -35.39365, -35.42291, -35.45158, -35.47977, -35.50776, -35.53565, 
        -35.56358, -35.59183, -35.62019, -35.64917, -35.67881, -35.70895, 
        -35.73942, -35.76998, -35.80029, -35.8304, -35.86033, -35.88911, 
        -35.91916, -35.9498, -35.98089, -36.01229, -36.04387, -36.07558, 
        -36.10703, -36.13849, -36.16948, -36.19996, -36.22952, -36.25795, 
        -36.28515, -36.31125, -36.33655, -36.36139, -36.386, -36.4105, 
        -36.43502, -36.45938, -36.4835, -36.50632, -36.52958, -36.55191, 
        -36.57316, -36.59327, -36.61277, -36.63206, -36.65197, -36.67249, 
        -36.69403, -36.71579, -36.73723, -36.7581, -36.7781, -36.79733, 
        -36.8161, -36.83487, -36.85391, -36.87341, -36.89331, -36.91328, 
        -36.93292, -36.95172, -36.96949, -36.98555, -37.00219, -37.01874, 
        -37.035, -37.05094, -37.06662, -37.0826, -37.09925, -37.11695, 
        -37.13577, -37.15608, -37.17785, -37.20126, -37.2265, -37.25389, 
        -37.28341, -37.31492, -37.3494, -37.38657, -37.42654, -37.46912, 
        -37.51385, -37.55999, -37.60692, -37.65384, -37.69989, -37.74446, 
        -37.78615, -37.82669, -37.86535, -37.90263, -37.93902, -37.97497, 
        -38.01053, -38.04569, -38.08021, -38.1143, -38.14782, -38.18061, 
        -38.21255, -38.2437, -38.27394, -38.30365, -38.33294, -38.36176, 
        -38.39036, -38.41872, -38.44658, -38.47355, -38.4994, -38.52409, 
        -38.54786, -38.57113, -38.59394, -38.6162, -38.63768, -38.65813, 
        -38.67722, -38.69443, -38.70863, -38.72206, -38.73383, -38.74422, 
        -38.75372, -38.76265, -38.77109, -38.77939, -38.78753, -38.79572, 
        -38.80438, -38.81353, -38.82269, -38.83148, -38.83961, -38.84693, 
        -38.85325, -38.85847, -38.86233, -38.86449, -38.86502, -38.86397, 
        -38.86155, -38.85796, -38.85347, -38.84836, -38.84254, -38.83582, 
        -38.8273, -38.81639, -38.80321, -38.78841, -38.77258, -38.75679, 
        -38.74134, -38.72626, -38.71109, -38.69509, -38.67759, -38.65682, 
        -38.63406, -38.60797, -38.57832, -38.54472, -38.50728, -38.46536, 
        -38.41794, -38.36357, -38.30042, -38.22643, -38.1411, -38.04507, 
        -37.94132, -37.83628, -37.73722, -37.65099, -37.58392, -37.53905, 
        -37.51754,
  -29.81296, -29.85794, -29.90313, -29.94854, -29.9944, -30.04085, 
        -30.08815, -30.13622, -30.18501, -30.23465, -30.28535, -30.33622, 
        -30.38927, -30.44324, -30.49801, -30.55313, -30.60806, -30.66212, 
        -30.71539, -30.76795, -30.82005, -30.87206, -30.9239, -30.97542, 
        -31.02657, -31.07756, -31.12757, -31.17847, -31.22951, -31.28081, 
        -31.33245, -31.38446, -31.43668, -31.48888, -31.54124, -31.59388, 
        -31.64689, -31.70004, -31.75303, -31.80561, -31.85775, -31.90853, 
        -31.95987, -32.01084, -32.06186, -32.11307, -32.16476, -32.21674, 
        -32.26874, -32.32017, -32.37109, -32.42125, -32.47076, -32.52, 
        -32.56897, -32.61778, -32.66635, -32.71338, -32.76085, -32.80805, 
        -32.85537, -32.90301, -32.9509, -32.99882, -33.04658, -33.09428, 
        -33.14198, -33.19018, -33.23912, -33.2888, -33.33932, -33.39047, 
        -33.44205, -33.49382, -33.54405, -33.59433, -33.64352, -33.69202, 
        -33.73997, -33.78812, -33.83652, -33.88479, -33.93197, -33.9784, 
        -34.02326, -34.06677, -34.10938, -34.15146, -34.19329, -34.2351, 
        -34.27701, -34.31935, -34.36132, -34.40488, -34.44864, -34.49168, 
        -34.53366, -34.57428, -34.61387, -34.65256, -34.69075, -34.72882, 
        -34.76656, -34.8042, -34.84127, -34.87764, -34.91319, -34.94792, 
        -34.9819, -35.01537, -35.04756, -35.08055, -35.11331, -35.14548, 
        -35.17688, -35.20747, -35.23726, -35.2667, -35.2959, -35.32503, 
        -35.354, -35.38259, -35.41065, -35.43832, -35.46588, -35.49338, 
        -35.52086, -35.5486, -35.57649, -35.60497, -35.63321, -35.66293, 
        -35.69287, -35.7229, -35.75281, -35.78238, -35.81194, -35.84141, 
        -35.87117, -35.90144, -35.93224, -35.96343, -35.9949, -36.02658, 
        -36.05812, -36.08961, -36.12083, -36.15151, -36.1813, -36.20988, 
        -36.23722, -36.26326, -36.2874, -36.312, -36.33622, -36.36031, 
        -36.38429, -36.40821, -36.43204, -36.45563, -36.47867, -36.50078, 
        -36.52164, -36.54126, -36.56002, -36.57873, -36.59785, -36.61795, 
        -36.63896, -36.66064, -36.6821, -36.70313, -36.72323, -36.74257, 
        -36.76146, -36.77931, -36.7985, -36.81816, -36.8383, -36.85859, 
        -36.87841, -36.89718, -36.91462, -36.93113, -36.94739, -36.96345, 
        -36.97937, -36.99519, -37.01097, -37.02719, -37.0443, -37.06261, 
        -37.08228, -37.1032, -37.12552, -37.14939, -37.17507, -37.20282, 
        -37.23284, -37.26536, -37.30071, -37.33817, -37.37954, -37.42363, 
        -37.46992, -37.51766, -37.56605, -37.61416, -37.6613, -37.70657, 
        -37.74962, -37.79036, -37.82903, -37.86631, -37.90299, -37.93919, 
        -37.97537, -38.01136, -38.04663, -38.08127, -38.11515, -38.14792, 
        -38.17941, -38.21008, -38.23965, -38.26862, -38.29719, -38.32564, 
        -38.35394, -38.38239, -38.41066, -38.43714, -38.46349, -38.48842, 
        -38.51235, -38.53576, -38.55879, -38.58143, -38.60337, -38.62414, 
        -38.64329, -38.66047, -38.67553, -38.68863, -38.69997, -38.70996, 
        -38.71901, -38.72747, -38.73565, -38.74371, -38.75187, -38.76027, 
        -38.76905, -38.77821, -38.78746, -38.79641, -38.80476, -38.81237, 
        -38.81905, -38.8245, -38.82831, -38.83039, -38.83051, -38.82895, 
        -38.82586, -38.82169, -38.81676, -38.81053, -38.80496, -38.79868, 
        -38.79073, -38.78041, -38.76763, -38.75291, -38.73714, -38.72147, 
        -38.70612, -38.69143, -38.67665, -38.66118, -38.64423, -38.62496, 
        -38.60267, -38.57678, -38.54698, -38.51316, -38.4753, -38.43262, 
        -38.38416, -38.3284, -38.26339, -38.18735, -38.0994, -38.00121, 
        -37.89559, -37.789, -37.68834, -37.60102, -37.53275, -37.4876, 
        -37.46587,
  -29.78176, -29.82617, -29.87077, -29.91558, -29.96083, -30.00688, 
        -30.05393, -30.10079, -30.14964, -30.19948, -30.25055, -30.30288, 
        -30.35638, -30.41098, -30.46626, -30.52178, -30.57688, -30.63105, 
        -30.68437, -30.73686, -30.78911, -30.84018, -30.8919, -30.94347, 
        -30.99486, -31.04602, -31.09718, -31.14832, -31.19943, -31.25041, 
        -31.30187, -31.35361, -31.4055, -31.45758, -31.50967, -31.56191, 
        -31.6135, -31.66613, -31.7184, -31.77022, -31.82163, -31.8727, 
        -31.92345, -31.97432, -32.02534, -32.07671, -32.12836, -32.18014, 
        -32.23167, -32.28275, -32.33318, -32.38296, -32.43123, -32.48018, 
        -32.52887, -32.57719, -32.62522, -32.67291, -32.72036, -32.76781, 
        -32.81571, -32.86389, -32.91235, -32.96072, -33.00871, -33.05641, 
        -33.10398, -33.15186, -33.20044, -33.24899, -33.29939, -33.35056, 
        -33.40245, -33.45459, -33.50627, -33.55709, -33.60695, -33.65587, 
        -33.7044, -33.75261, -33.80083, -33.84876, -33.89586, -33.94187, 
        -33.98645, -34.0297, -34.07125, -34.11361, -34.15591, -34.19825, 
        -34.24061, -34.28334, -34.32669, -34.37057, -34.41458, -34.45799, 
        -34.50026, -34.5412, -34.58078, -34.61944, -34.65753, -34.69555, 
        -34.73343, -34.77131, -34.80762, -34.84402, -34.87932, -34.91362, 
        -34.94711, -34.98022, -35.01315, -35.04602, -35.07869, -35.11056, 
        -35.14151, -35.17154, -35.20078, -35.22956, -35.25809, -35.28645, 
        -35.31454, -35.34221, -35.36957, -35.39668, -35.42271, -35.44984, 
        -35.47688, -35.5042, -35.53176, -35.55994, -35.58862, -35.61769, 
        -35.64698, -35.67656, -35.70597, -35.73514, -35.76438, -35.79362, 
        -35.82322, -35.85328, -35.88385, -35.91473, -35.9459, -35.97728, 
        -36.00859, -36.03885, -36.06994, -36.10044, -36.13011, -36.15867, 
        -36.18587, -36.21202, -36.23708, -36.26152, -36.28564, -36.3095, 
        -36.33318, -36.35691, -36.38058, -36.40405, -36.42694, -36.44882, 
        -36.46936, -36.48857, -36.50696, -36.52521, -36.54397, -36.56265, 
        -36.58342, -36.6049, -36.62643, -36.64759, -36.66791, -36.6874, 
        -36.70631, -36.72514, -36.74417, -36.76387, -36.78419, -36.80474, 
        -36.82474, -36.84369, -36.86127, -36.8778, -36.89373, -36.9096, 
        -36.92533, -36.94096, -36.95677, -36.97313, -36.99055, -37.00931, 
        -37.02848, -37.04999, -37.07291, -37.09742, -37.12378, -37.15219, 
        -37.18293, -37.21628, -37.25241, -37.29186, -37.3345, -37.38003, 
        -37.42777, -37.477, -37.52671, -37.57593, -37.62384, -37.6696, 
        -37.71287, -37.75361, -37.79249, -37.82969, -37.86639, -37.90337, 
        -37.94015, -37.97665, -38.01275, -38.04799, -38.08209, -38.11379, 
        -38.14495, -38.17492, -38.20396, -38.23217, -38.26008, -38.28804, 
        -38.3162, -38.34467, -38.3733, -38.40128, -38.42805, -38.45326, 
        -38.47741, -38.50083, -38.52381, -38.54646, -38.56852, -38.58934, 
        -38.60838, -38.62555, -38.6407, -38.6537, -38.66496, -38.67473, 
        -38.68356, -38.69182, -38.70004, -38.70837, -38.71696, -38.72559, 
        -38.73443, -38.74341, -38.75235, -38.75997, -38.76813, -38.77567, 
        -38.78246, -38.78796, -38.79174, -38.79368, -38.79331, -38.79115, 
        -38.78749, -38.78291, -38.7779, -38.77289, -38.76773, -38.76199, 
        -38.75464, -38.74484, -38.73244, -38.71812, -38.70287, -38.68763, 
        -38.6729, -38.65869, -38.64434, -38.62917, -38.6124, -38.59345, 
        -38.57154, -38.54584, -38.51599, -38.48183, -38.44342, -38.40028, 
        -38.35106, -38.29413, -38.22741, -38.14913, -38.05868, -37.95744, 
        -37.84912, -37.73952, -37.63606, -37.54631, -37.47644, -37.42915, 
        -37.40693,
  -29.75188, -29.79572, -29.83873, -29.88302, -29.9279, -29.97362, 
        -30.02048, -30.06855, -30.11763, -30.16779, -30.21916, -30.27177, 
        -30.32567, -30.38052, -30.43604, -30.49187, -30.54702, -30.60027, 
        -30.6537, -30.70624, -30.75852, -30.8105, -30.86233, -30.91391, 
        -30.96536, -31.01664, -31.06785, -31.11894, -31.16988, -31.22082, 
        -31.27202, -31.32354, -31.3743, -31.42605, -31.47787, -31.52979, 
        -31.58183, -31.63377, -31.6853, -31.73633, -31.78695, -31.83736, 
        -31.88785, -31.93857, -31.98966, -32.04115, -32.09264, -32.14292, 
        -32.19374, -32.24404, -32.29378, -32.34288, -32.39178, -32.4404, 
        -32.4888, -32.53699, -32.58493, -32.63271, -32.68053, -32.72859, 
        -32.77709, -32.82581, -32.87452, -32.92211, -32.97026, -33.01795, 
        -33.06544, -33.11319, -33.16166, -33.2111, -33.26155, -33.31302, 
        -33.36526, -33.41775, -33.46991, -33.52126, -33.57154, -33.62099, 
        -33.66967, -33.71814, -33.76528, -33.81288, -33.85955, -33.90505, 
        -33.94931, -33.99261, -34.03535, -34.07804, -34.12075, -34.16362, 
        -34.2065, -34.24954, -34.29301, -34.33696, -34.38102, -34.42461, 
        -34.467, -34.50803, -34.54681, -34.58562, -34.62389, -34.66216, 
        -34.7004, -34.73846, -34.77597, -34.8124, -34.84735, -34.88118, 
        -34.91423, -34.94693, -34.97957, -35.01207, -35.04438, -35.07595, 
        -35.10649, -35.13593, -35.16452, -35.19149, -35.2191, -35.24657, 
        -35.27376, -35.30063, -35.32718, -35.35381, -35.38061, -35.4074, 
        -35.43422, -35.46119, -35.48849, -35.51619, -35.54436, -35.57272, 
        -35.60139, -35.63032, -35.65936, -35.68834, -35.71733, -35.74645, 
        -35.77491, -35.80481, -35.83493, -35.8653, -35.89581, -35.92649, 
        -35.95729, -35.98807, -36.01871, -36.04889, -36.07825, -36.10652, 
        -36.13366, -36.1596, -36.18473, -36.20916, -36.23326, -36.25706, 
        -36.28069, -36.30439, -36.32806, -36.35152, -36.37335, -36.39516, 
        -36.41558, -36.43468, -36.45301, -36.47094, -36.48959, -36.50908, 
        -36.52963, -36.5508, -36.57246, -36.59367, -36.61419, -36.63383, 
        -36.65279, -36.67146, -36.69033, -36.70971, -36.72994, -36.75052, 
        -36.77068, -36.78984, -36.80775, -36.82462, -36.83986, -36.8558, 
        -36.87147, -36.88706, -36.90286, -36.91922, -36.93677, -36.95583, 
        -36.9763, -36.99826, -37.02167, -37.04689, -37.07408, -37.10334, 
        -37.13496, -37.16916, -37.20633, -37.2469, -37.29074, -37.33751, 
        -37.38674, -37.43747, -37.48848, -37.53872, -37.58718, -37.63327, 
        -37.67665, -37.71636, -37.75526, -37.79267, -37.82944, -37.86649, 
        -37.90393, -37.94114, -37.97795, -38.0137, -38.04794, -38.08054, 
        -38.11141, -38.14074, -38.16901, -38.19673, -38.22409, -38.25141, 
        -38.27952, -38.30804, -38.3368, -38.36499, -38.39195, -38.41743, 
        -38.44167, -38.46499, -38.48779, -38.51028, -38.53212, -38.5528, 
        -38.57188, -38.5891, -38.60423, -38.61652, -38.62784, -38.6376, 
        -38.64644, -38.65476, -38.66318, -38.67186, -38.68082, -38.68972, 
        -38.69849, -38.70714, -38.71558, -38.72392, -38.73172, -38.73888, 
        -38.74535, -38.75072, -38.75455, -38.75622, -38.75552, -38.7533, 
        -38.74934, -38.74478, -38.73978, -38.73504, -38.73027, -38.72489, 
        -38.71798, -38.70864, -38.69682, -38.68317, -38.66873, -38.65431, 
        -38.64037, -38.6267, -38.61271, -38.59772, -38.58109, -38.56227, 
        -38.54044, -38.51384, -38.48403, -38.44986, -38.41119, -38.36763, 
        -38.31785, -38.25988, -38.19158, -38.11108, -38.01775, -37.91324, 
        -37.80143, -37.6877, -37.58061, -37.48708, -37.41463, -37.3663, 
        -37.34324,
  -29.72253, -29.76605, -29.80949, -29.85322, -29.89769, -29.94327, 
        -29.99017, -30.03851, -30.08809, -30.1387, -30.19039, -30.24305, 
        -30.29595, -30.35087, -30.40654, -30.46221, -30.51731, -30.57149, 
        -30.6249, -30.67754, -30.72972, -30.78172, -30.83352, -30.88521, 
        -30.93667, -30.98799, -31.03909, -31.08901, -31.13977, -31.19053, 
        -31.24155, -31.29292, -31.3446, -31.39631, -31.44804, -31.49943, 
        -31.55092, -31.60206, -31.65266, -31.70278, -31.75263, -31.80252, 
        -31.85173, -31.90245, -31.95365, -32.00525, -32.05649, -32.10714, 
        -32.15704, -32.20621, -32.25489, -32.30335, -32.35159, -32.39997, 
        -32.44823, -32.49654, -32.54478, -32.59316, -32.64068, -32.68945, 
        -32.7385, -32.78755, -32.83638, -32.88497, -32.93308, -32.98068, 
        -33.02814, -33.07581, -33.12421, -33.17371, -33.22446, -33.27629, 
        -33.32897, -33.3819, -33.43453, -33.48537, -33.53612, -33.58595, 
        -33.63503, -33.68343, -33.7313, -33.77856, -33.82476, -33.86982, 
        -33.91396, -33.95713, -34.0001, -34.04338, -34.08667, -34.12992, 
        -34.17309, -34.21639, -34.25896, -34.30286, -34.34678, -34.39013, 
        -34.43249, -34.47359, -34.51355, -34.55269, -34.59128, -34.62993, 
        -34.66857, -34.707, -34.74465, -34.78082, -34.81563, -34.84901, 
        -34.88178, -34.914, -34.94621, -34.97726, -35.00903, -35.04008, 
        -35.07013, -35.09904, -35.12687, -35.15401, -35.18073, -35.20717, 
        -35.23343, -35.25961, -35.2856, -35.3119, -35.33838, -35.36495, 
        -35.39171, -35.41854, -35.44577, -35.47309, -35.50067, -35.5274, 
        -35.55522, -35.58356, -35.61223, -35.64093, -35.6699, -35.69901, 
        -35.72841, -35.75796, -35.78754, -35.81716, -35.84674, -35.87652, 
        -35.90648, -35.93662, -35.96666, -35.99633, -36.02526, -36.05316, 
        -36.07998, -36.10579, -36.13086, -36.15433, -36.17847, -36.20237, 
        -36.22612, -36.24991, -36.27365, -36.2972, -36.32012, -36.34194, 
        -36.36247, -36.38175, -36.40015, -36.41834, -36.43671, -36.45627, 
        -36.47657, -36.4977, -36.519, -36.54024, -36.56084, -36.58057, 
        -36.5995, -36.61796, -36.63554, -36.65471, -36.67439, -36.69466, 
        -36.71487, -36.73435, -36.75292, -36.77047, -36.78732, -36.80363, 
        -36.81937, -36.83496, -36.85067, -36.86721, -36.88468, -36.90373, 
        -36.92436, -36.94663, -36.97064, -36.99659, -37.02487, -37.05525, 
        -37.08797, -37.12343, -37.16183, -37.20353, -37.24747, -37.29559, 
        -37.34618, -37.39821, -37.45042, -37.50151, -37.55044, -37.5966, 
        -37.63992, -37.68058, -37.71914, -37.75666, -37.79392, -37.83131, 
        -37.86922, -37.90718, -37.9445, -37.98055, -38.01488, -38.04721, 
        -38.07752, -38.10607, -38.13345, -38.16031, -38.18736, -38.21469, 
        -38.24277, -38.27131, -38.30011, -38.32835, -38.35439, -38.37998, 
        -38.40411, -38.42728, -38.4499, -38.47192, -38.49334, -38.51366, 
        -38.53262, -38.54997, -38.56557, -38.57908, -38.59063, -38.60062, 
        -38.60955, -38.61816, -38.62677, -38.63575, -38.64471, -38.65367, 
        -38.66241, -38.67054, -38.6784, -38.68603, -38.69352, -38.7003, 
        -38.70635, -38.71146, -38.71506, -38.71658, -38.71617, -38.71385, 
        -38.71009, -38.70588, -38.70139, -38.69698, -38.69262, -38.6866, 
        -38.67994, -38.67094, -38.65975, -38.64693, -38.63342, -38.61993, 
        -38.60681, -38.59378, -38.58019, -38.56535, -38.54872, -38.52982, 
        -38.50804, -38.48246, -38.45271, -38.41858, -38.37994, -38.33628, 
        -38.28617, -38.22733, -38.15763, -38.07503, -37.97918, -37.87107, 
        -37.75498, -37.63671, -37.52533, -37.42704, -37.35064, -37.29987, 
        -37.27612,
  -29.69519, -29.73881, -29.78218, -29.82559, -29.86971, -29.91514, 
        -29.96208, -30.00961, -30.05951, -30.11048, -30.1623, -30.21503, 
        -30.26882, -30.32357, -30.37898, -30.43445, -30.48937, -30.54344, 
        -30.59662, -30.64916, -30.70128, -30.75326, -30.80411, -30.85578, 
        -30.90734, -30.95859, -31.00963, -31.06031, -31.11085, -31.16135, 
        -31.21221, -31.26348, -31.31509, -31.36681, -31.41828, -31.46934, 
        -31.52017, -31.5695, -31.61917, -31.66842, -31.71756, -31.76701, 
        -31.81709, -31.86786, -31.91915, -31.97049, -32.02132, -32.07129, 
        -32.12031, -32.16859, -32.21642, -32.26404, -32.3119, -32.35894, 
        -32.40715, -32.45567, -32.50442, -32.55353, -32.60291, -32.65247, 
        -32.70193, -32.75108, -32.7999, -32.84821, -32.89628, -32.94392, 
        -32.99137, -33.0391, -33.08755, -33.1361, -33.18695, -33.23913, 
        -33.29218, -33.34553, -33.39855, -33.45076, -33.50192, -33.55209, 
        -33.60136, -33.64986, -33.69764, -33.74447, -33.79025, -33.83497, 
        -33.87922, -33.92274, -33.96629, -34.00895, -34.05264, -34.09604, 
        -34.13926, -34.18255, -34.22601, -34.26976, -34.3134, -34.35654, 
        -34.39871, -34.43985, -34.48011, -34.51964, -34.55878, -34.59779, 
        -34.63673, -34.67521, -34.71269, -34.74765, -34.78199, -34.81517, 
        -34.84768, -34.87952, -34.9115, -34.94306, -34.97439, -35.00507, 
        -35.03455, -35.06284, -35.08995, -35.11631, -35.14209, -35.16768, 
        -35.19305, -35.21854, -35.24425, -35.27035, -35.29665, -35.32215, 
        -35.34871, -35.37538, -35.40251, -35.42949, -35.45642, -35.48378, 
        -35.51086, -35.53835, -35.56665, -35.59519, -35.62417, -35.65336, 
        -35.68248, -35.71165, -35.74062, -35.76925, -35.79784, -35.82657, 
        -35.85558, -35.88494, -35.91335, -35.94241, -35.97084, -35.99832, 
        -36.02477, -36.05036, -36.07531, -36.09991, -36.12418, -36.14828, 
        -36.17225, -36.19623, -36.22009, -36.24368, -36.26656, -36.28845, 
        -36.30909, -36.32866, -36.34733, -36.36591, -36.3844, -36.40387, 
        -36.42279, -36.44363, -36.46466, -36.48575, -36.50629, -36.52608, 
        -36.5451, -36.56361, -36.58202, -36.60076, -36.62012, -36.63978, 
        -36.65996, -36.67987, -36.69873, -36.71719, -36.73494, -36.75176, 
        -36.76791, -36.7834, -36.79908, -36.81547, -36.8329, -36.85209, 
        -36.87281, -36.8955, -36.91891, -36.94605, -36.97546, -37.00725, 
        -37.04145, -37.07845, -37.11827, -37.16143, -37.2078, -37.25714, 
        -37.30881, -37.36174, -37.41463, -37.46619, -37.5153, -37.56144, 
        -37.60453, -37.64499, -37.6835, -37.72115, -37.75872, -37.79678, 
        -37.83533, -37.87378, -37.9114, -37.94752, -37.98166, -38.01355, 
        -38.04217, -38.06986, -38.09652, -38.1226, -38.14922, -38.17628, 
        -38.20456, -38.23329, -38.26209, -38.29016, -38.31703, -38.34245, 
        -38.36653, -38.38957, -38.41195, -38.43372, -38.45474, -38.47482, 
        -38.49372, -38.51124, -38.52706, -38.5409, -38.55282, -38.56299, 
        -38.5721, -38.58081, -38.58946, -38.59847, -38.60726, -38.61619, 
        -38.62443, -38.63248, -38.63968, -38.64687, -38.6524, -38.65856, 
        -38.66423, -38.66908, -38.67253, -38.67428, -38.67414, -38.67243, 
        -38.66945, -38.66578, -38.66194, -38.65802, -38.65389, -38.64891, 
        -38.64241, -38.63384, -38.62337, -38.61145, -38.59879, -38.58619, 
        -38.57389, -38.56152, -38.54845, -38.53384, -38.51731, -38.49831, 
        -38.47633, -38.4507, -38.42097, -38.38692, -38.34836, -38.30478, 
        -38.25444, -38.19513, -38.12415, -38.03973, -37.94088, -37.82954, 
        -37.70926, -37.58652, -37.46961, -37.36626, -37.28493, -37.23099, 
        -37.20592,
  -29.66929, -29.71322, -29.75653, -29.79897, -29.84301, -29.88825, 
        -29.93517, -29.98375, -30.03366, -30.08453, -30.13633, -30.18895, 
        -30.24256, -30.29712, -30.3523, -30.40751, -30.46218, -30.51503, 
        -30.56801, -30.62038, -30.67229, -30.72421, -30.77596, -30.82774, 
        -30.87921, -30.93044, -30.98134, -31.0318, -31.08202, -31.13229, 
        -31.1829, -31.23406, -31.28461, -31.33615, -31.38739, -31.43809, 
        -31.48819, -31.53769, -31.5866, -31.63513, -31.68372, -31.73281, 
        -31.78272, -31.83337, -31.88457, -31.93558, -31.98589, -32.03521, 
        -32.08255, -32.13018, -32.17749, -32.22476, -32.27232, -32.32024, 
        -32.36858, -32.41734, -32.4666, -32.51637, -32.56649, -32.61663, 
        -32.66641, -32.71562, -32.76431, -32.81252, -32.85938, -32.90702, 
        -32.95455, -33.00229, -33.05067, -33.10014, -33.1511, -33.20343, 
        -33.25673, -33.31031, -33.36354, -33.41592, -33.46734, -33.51775, 
        -33.56725, -33.61587, -33.66349, -33.70916, -33.7548, -33.79957, 
        -33.844, -33.88808, -33.93226, -33.97641, -34.02027, -34.06372, 
        -34.10683, -34.14982, -34.19301, -34.2365, -34.27978, -34.32268, 
        -34.36477, -34.40622, -34.44687, -34.48587, -34.52539, -34.56465, 
        -34.60356, -34.6417, -34.6787, -34.71422, -34.74826, -34.78123, 
        -34.8135, -34.84535, -34.87708, -34.90844, -34.93938, -34.96955, 
        -34.99858, -35.02637, -35.05281, -35.07834, -35.10243, -35.1273, 
        -35.15216, -35.1773, -35.20279, -35.22869, -35.25483, -35.28106, 
        -35.30738, -35.3338, -35.36066, -35.38747, -35.41393, -35.44036, 
        -35.46706, -35.49394, -35.52177, -35.55034, -35.57914, -35.6083, 
        -35.63706, -35.66484, -35.69299, -35.72072, -35.74819, -35.77582, 
        -35.80397, -35.83261, -35.86139, -35.88983, -35.91768, -35.94471, 
        -35.97081, -35.99627, -36.02108, -36.04568, -36.07006, -36.09441, 
        -36.11861, -36.14273, -36.16671, -36.1903, -36.21315, -36.23405, 
        -36.25478, -36.27441, -36.29342, -36.31202, -36.33063, -36.34988, 
        -36.36975, -36.39027, -36.41114, -36.43199, -36.45245, -36.47235, 
        -36.4916, -36.51029, -36.52867, -36.54719, -36.56614, -36.58554, 
        -36.60543, -36.62537, -36.64497, -36.66426, -36.68267, -36.69908, 
        -36.71543, -36.73138, -36.74711, -36.76338, -36.78101, -36.80006, 
        -36.82065, -36.8436, -36.86906, -36.89739, -36.92813, -36.96163, 
        -36.99781, -37.03658, -37.07822, -37.12287, -37.17052, -37.22095, 
        -37.2734, -37.32684, -37.38, -37.43157, -37.48053, -37.52645, 
        -37.56933, -37.60964, -37.64823, -37.68515, -37.72322, -37.76188, 
        -37.80093, -37.83969, -37.87739, -37.91331, -37.94701, -37.97826, 
        -38.00708, -38.03398, -38.05969, -38.08509, -38.11126, -38.13851, 
        -38.16685, -38.19565, -38.2243, -38.25211, -38.27865, -38.30381, 
        -38.32779, -38.35078, -38.37305, -38.3947, -38.41559, -38.4356, 
        -38.45457, -38.4723, -38.48833, -38.50236, -38.51443, -38.52376, 
        -38.53294, -38.54158, -38.55005, -38.55876, -38.56743, -38.57567, 
        -38.58374, -38.59145, -38.59823, -38.60441, -38.61039, -38.61592, 
        -38.62113, -38.62566, -38.62913, -38.63127, -38.63184, -38.63107, 
        -38.62914, -38.62644, -38.62327, -38.61975, -38.61568, -38.61063, 
        -38.60412, -38.59587, -38.58606, -38.57488, -38.56313, -38.5514, 
        -38.53979, -38.52814, -38.51568, -38.50164, -38.48534, -38.46629, 
        -38.44412, -38.4183, -38.3886, -38.35357, -38.31517, -38.2718, 
        -38.22142, -38.16151, -38.08944, -38.0033, -37.902, -37.78766, 
        -37.66303, -37.53612, -37.41343, -37.30426, -37.21794, -37.16054, 
        -37.13417,
  -29.64328, -29.68765, -29.73149, -29.77527, -29.81945, -29.86471, 
        -29.91145, -29.95976, -30.00928, -30.05997, -30.11145, -30.16379, 
        -30.21709, -30.2703, -30.32517, -30.38016, -30.43464, -30.48834, 
        -30.54116, -30.59333, -30.64518, -30.69686, -30.74844, -30.80011, 
        -30.85145, -30.9026, -30.9533, -31.00249, -31.0524, -31.10234, 
        -31.15267, -31.20355, -31.25483, -31.30609, -31.35694, -31.4072, 
        -31.45681, -31.50575, -31.5541, -31.60211, -31.6503, -31.6991, 
        -31.74876, -31.79823, -31.84905, -31.89961, -31.94935, -31.99813, 
        -32.04607, -32.09345, -32.14066, -32.188, -32.23565, -32.28372, 
        -32.33223, -32.38122, -32.43082, -32.48104, -32.53157, -32.58106, 
        -32.63102, -32.68033, -32.72894, -32.77691, -32.8247, -32.8723, 
        -32.91987, -32.96762, -33.01598, -33.06526, -33.11612, -33.16837, 
        -33.2216, -33.27509, -33.32825, -33.3806, -33.43105, -33.48168, 
        -33.53121, -33.57994, -33.62766, -33.67447, -33.72014, -33.76536, 
        -33.81022, -33.85501, -33.89978, -33.94436, -33.98841, -34.03178, 
        -34.07458, -34.11723, -34.15998, -34.20207, -34.24519, -34.28798, 
        -34.33037, -34.37203, -34.41309, -34.4535, -34.49328, -34.53244, 
        -34.57093, -34.60843, -34.64465, -34.6796, -34.71326, -34.74611, 
        -34.77842, -34.81042, -34.84202, -34.87323, -34.90285, -34.93266, 
        -34.96128, -34.98854, -35.01447, -35.03944, -35.06396, -35.08835, 
        -35.11292, -35.13786, -35.16324, -35.18906, -35.21497, -35.24089, 
        -35.26679, -35.29283, -35.31911, -35.34546, -35.37159, -35.39736, 
        -35.42236, -35.44881, -35.4764, -35.50475, -35.53363, -35.56274, 
        -35.59135, -35.61956, -35.64695, -35.67377, -35.70031, -35.72708, 
        -35.75437, -35.78217, -35.81032, -35.83817, -35.86549, -35.89209, 
        -35.9179, -35.94307, -35.96779, -35.99238, -36.01586, -36.04031, 
        -36.06467, -36.08895, -36.11301, -36.13658, -36.15941, -36.18125, 
        -36.20198, -36.22155, -36.24044, -36.25896, -36.27766, -36.29683, 
        -36.31664, -36.33701, -36.35765, -36.37833, -36.39876, -36.41875, 
        -36.43821, -36.45712, -36.47562, -36.49309, -36.51184, -36.53098, 
        -36.55069, -36.57079, -36.59093, -36.61074, -36.62973, -36.64775, 
        -36.6646, -36.6806, -36.69645, -36.71295, -36.73047, -36.7496, 
        -36.77068, -36.79409, -36.82043, -36.8498, -36.88231, -36.9177, 
        -36.95584, -36.99674, -37.04034, -37.08667, -37.13558, -37.18689, 
        -37.23888, -37.29257, -37.34562, -37.39681, -37.4453, -37.49077, 
        -37.53341, -37.57369, -37.61246, -37.65089, -37.68948, -37.72859, 
        -37.76788, -37.80674, -37.84429, -37.87971, -37.9128, -37.94327, 
        -37.97128, -37.99731, -38.02232, -38.04724, -38.07306, -38.10019, 
        -38.12841, -38.15717, -38.18559, -38.21304, -38.23919, -38.26415, 
        -38.28696, -38.30997, -38.33227, -38.35392, -38.37488, -38.39508, 
        -38.41431, -38.43227, -38.44814, -38.46244, -38.47464, -38.48489, 
        -38.49392, -38.50229, -38.51042, -38.51872, -38.52699, -38.53514, 
        -38.54268, -38.54975, -38.55598, -38.56156, -38.56665, -38.57153, 
        -38.57618, -38.58038, -38.58406, -38.58672, -38.58827, -38.58865, 
        -38.58787, -38.58627, -38.58379, -38.58057, -38.57644, -38.57119, 
        -38.56455, -38.55546, -38.54608, -38.53566, -38.52464, -38.51345, 
        -38.50269, -38.49189, -38.48028, -38.46688, -38.45114, -38.43235, 
        -38.41017, -38.38416, -38.35427, -38.32032, -38.28216, -38.23868, 
        -38.18821, -38.12787, -38.05499, -37.96738, -37.86424, -37.74696, 
        -37.61925, -37.4877, -37.36005, -37.24578, -37.15478, -37.0934, 
        -37.06506,
  -29.61885, -29.66398, -29.7086, -29.75306, -29.79777, -29.84329, 
        -29.88998, -29.93789, -29.98591, -30.03606, -30.08703, -30.13887, 
        -30.1918, -30.24562, -30.30006, -30.35452, -30.40887, -30.46249, 
        -30.51525, -30.56731, -30.61898, -30.67047, -30.72187, -30.77218, 
        -30.82329, -30.87409, -30.9245, -30.97445, -31.02405, -31.07363, 
        -31.12359, -31.17414, -31.22495, -31.27576, -31.32617, -31.37608, 
        -31.42535, -31.47398, -31.52104, -31.56882, -31.61671, -31.66518, 
        -31.71458, -31.76461, -31.81496, -31.86495, -31.91423, -31.9627, 
        -32.01059, -32.05804, -32.10544, -32.15306, -32.20103, -32.24939, 
        -32.29715, -32.3464, -32.39622, -32.4466, -32.49723, -32.5479, 
        -32.598, -32.64731, -32.69582, -32.74373, -32.79135, -32.83894, 
        -32.88652, -32.93434, -32.98252, -33.03171, -33.08131, -33.13314, 
        -33.18599, -33.23906, -33.29186, -33.34393, -33.39516, -33.44547, 
        -33.49517, -33.54406, -33.59206, -33.63915, -33.68541, -33.73113, 
        -33.77658, -33.82198, -33.86729, -33.9123, -33.95552, -33.99889, 
        -34.04153, -34.08372, -34.12609, -34.16878, -34.21168, -34.25457, 
        -34.29716, -34.33928, -34.3809, -34.42166, -34.46141, -34.50029, 
        -34.53812, -34.57476, -34.61007, -34.64431, -34.67662, -34.70936, 
        -34.74168, -34.77374, -34.80547, -34.83662, -34.8671, -34.89662, 
        -34.92489, -34.95179, -34.97736, -35.00196, -35.02608, -35.05017, 
        -35.0746, -35.09938, -35.12466, -35.1503, -35.17589, -35.20135, 
        -35.22568, -35.25107, -35.27668, -35.30248, -35.32811, -35.35355, 
        -35.37907, -35.40526, -35.43248, -35.46068, -35.4896, -35.51848, 
        -35.54679, -35.57453, -35.60139, -35.62752, -35.65335, -35.67936, 
        -35.70593, -35.73306, -35.7605, -35.7868, -35.81363, -35.83981, 
        -35.86533, -35.89029, -35.91491, -35.93937, -35.96378, -35.98823, 
        -36.01273, -36.03713, -36.06131, -36.08497, -36.1078, -36.12948, 
        -36.15007, -36.16935, -36.18798, -36.20638, -36.22495, -36.24416, 
        -36.26403, -36.28335, -36.30399, -36.32459, -36.34492, -36.36489, 
        -36.38441, -36.40348, -36.42213, -36.44062, -36.45915, -36.47818, 
        -36.49787, -36.51799, -36.53836, -36.55869, -36.5783, -36.59679, 
        -36.6141, -36.63049, -36.64659, -36.66322, -36.68091, -36.70024, 
        -36.72166, -36.74576, -36.77301, -36.80266, -36.83674, -36.87404, 
        -36.91429, -36.95736, -37.00304, -37.0511, -37.10141, -37.15362, 
        -37.2071, -37.26078, -37.31361, -37.36425, -37.41199, -37.4569, 
        -37.49925, -37.53951, -37.57853, -37.61736, -37.65633, -37.69559, 
        -37.735, -37.7737, -37.81084, -37.84568, -37.87801, -37.90771, 
        -37.93494, -37.96035, -37.98372, -38.00821, -38.03369, -38.06047, 
        -38.08844, -38.11689, -38.14493, -38.17204, -38.19793, -38.22262, 
        -38.24641, -38.26943, -38.29183, -38.31364, -38.33485, -38.35537, 
        -38.37485, -38.39289, -38.40888, -38.42297, -38.4349, -38.44479, 
        -38.45367, -38.46194, -38.46983, -38.4778, -38.48575, -38.49347, 
        -38.50089, -38.50737, -38.51281, -38.51746, -38.52163, -38.52574, 
        -38.52868, -38.53265, -38.53648, -38.53959, -38.54209, -38.54369, 
        -38.54425, -38.54361, -38.54181, -38.53885, -38.53466, -38.52915, 
        -38.52221, -38.51399, -38.50477, -38.49474, -38.48436, -38.47406, 
        -38.46416, -38.45433, -38.44364, -38.43114, -38.41598, -38.39769, 
        -38.37569, -38.3498, -38.31977, -38.2858, -38.24757, -38.20411, 
        -38.15342, -38.09284, -38.01934, -37.93092, -37.82642, -37.70721, 
        -37.57694, -37.44176, -37.31008, -37.19168, -37.09615, -37.03109, 
        -36.99986,
  -29.59515, -29.64098, -29.68669, -29.73203, -29.77671, -29.82274, 
        -29.86952, -29.91699, -29.96543, -30.01484, -30.06521, -30.11666, 
        -30.16908, -30.22235, -30.27618, -30.33021, -30.38416, -30.43762, 
        -30.48941, -30.5415, -30.593, -30.64418, -30.6951, -30.74589, 
        -30.79649, -30.8469, -30.89705, -30.94681, -30.99623, -31.04546, 
        -31.09497, -31.14491, -31.19514, -31.24433, -31.29418, -31.34388, 
        -31.39299, -31.44163, -31.48974, -31.53744, -31.58517, -31.63342, 
        -31.68231, -31.73178, -31.78148, -31.83099, -31.87977, -31.92802, 
        -31.97612, -32.02299, -32.07098, -32.11922, -32.16773, -32.2164, 
        -32.26539, -32.31475, -32.36459, -32.41489, -32.46549, -32.51596, 
        -32.56609, -32.61546, -32.66391, -32.71172, -32.75922, -32.80574, 
        -32.85341, -32.90128, -32.94956, -32.99869, -33.04875, -33.10007, 
        -33.15216, -33.20452, -33.2565, -33.30809, -33.35893, -33.40906, 
        -33.45895, -33.50808, -33.55643, -33.60396, -33.64973, -33.69602, 
        -33.74206, -33.78794, -33.83368, -33.87896, -33.92342, -33.9669, 
        -34.00945, -34.05144, -34.09358, -34.13599, -34.17871, -34.22165, 
        -34.26457, -34.30723, -34.34921, -34.39022, -34.42903, -34.4674, 
        -34.50435, -34.53996, -34.57446, -34.60814, -34.64109, -34.67362, 
        -34.70592, -34.73806, -34.7699, -34.80107, -34.83145, -34.86075, 
        -34.88879, -34.91551, -34.94104, -34.96557, -34.98943, -35.01223, 
        -35.03648, -35.06104, -35.08612, -35.11129, -35.13641, -35.16124, 
        -35.18597, -35.2107, -35.23557, -35.26075, -35.2859, -35.31101, 
        -35.33628, -35.36218, -35.38909, -35.4171, -35.44576, -35.47445, 
        -35.50259, -35.52988, -35.55524, -35.58087, -35.60618, -35.63159, 
        -35.65756, -35.68409, -35.71092, -35.73768, -35.76406, -35.78986, 
        -35.81507, -35.83982, -35.86427, -35.88858, -35.9128, -35.93722, 
        -35.96178, -35.98642, -36.01077, -36.03451, -36.05735, -36.07898, 
        -36.09809, -36.1171, -36.13541, -36.15371, -36.17231, -36.19158, 
        -36.2115, -36.23196, -36.25262, -36.27313, -36.29327, -36.31313, 
        -36.33257, -36.35161, -36.37034, -36.38885, -36.40754, -36.42639, 
        -36.44576, -36.46589, -36.48648, -36.50717, -36.52726, -36.54626, 
        -36.56299, -36.57992, -36.59628, -36.61331, -36.63131, -36.65108, 
        -36.67302, -36.69781, -36.72601, -36.75789, -36.79347, -36.8325, 
        -36.87476, -36.91998, -36.96769, -37.01756, -37.06928, -37.12244, 
        -37.17641, -37.23027, -37.28277, -37.33311, -37.38003, -37.42431, 
        -37.46623, -37.50628, -37.5455, -37.58456, -37.62268, -37.66212, 
        -37.70146, -37.7397, -37.77624, -37.81042, -37.84199, -37.87091, 
        -37.89744, -37.92222, -37.94614, -37.97028, -37.9952, -38.02152, 
        -38.04899, -38.0769, -38.10451, -38.13121, -38.15681, -38.18144, 
        -38.20524, -38.22838, -38.25105, -38.2732, -38.29485, -38.31568, 
        -38.33528, -38.35338, -38.36918, -38.38281, -38.39415, -38.40394, 
        -38.41163, -38.41977, -38.42757, -38.43529, -38.44282, -38.4502, 
        -38.45708, -38.463, -38.46782, -38.47159, -38.47502, -38.4782, 
        -38.48164, -38.48545, -38.48905, -38.49264, -38.49592, -38.4985, 
        -38.50003, -38.50024, -38.49898, -38.49625, -38.49198, -38.48615, 
        -38.47884, -38.47042, -38.46119, -38.4515, -38.44174, -38.43214, 
        -38.42313, -38.41421, -38.40462, -38.39319, -38.37892, -38.36118, 
        -38.33958, -38.31398, -38.2841, -38.24999, -38.21163, -38.1669, 
        -38.11591, -38.05512, -37.9814, -37.89278, -37.78794, -37.66801, 
        -37.53621, -37.39898, -37.26446, -37.14258, -37.0431, -36.97441, 
        -36.94032,
  -29.57162, -29.61805, -29.6646, -29.71114, -29.75778, -29.80452, 
        -29.85126, -29.89858, -29.9464, -29.99525, -30.04526, -30.09628, 
        -30.14837, -30.19996, -30.25303, -30.30637, -30.35979, -30.41296, 
        -30.46574, -30.5178, -30.5693, -30.62021, -30.6706, -30.72073, 
        -30.77071, -30.82069, -30.87046, -30.91998, -30.96809, -31.01705, 
        -31.06601, -31.11518, -31.16454, -31.21399, -31.26346, -31.31275, 
        -31.36201, -31.41093, -31.4593, -31.50711, -31.55474, -31.60264, 
        -31.65103, -31.69987, -31.74776, -31.79679, -31.84528, -31.89356, 
        -31.94206, -31.99051, -32.03925, -32.08807, -32.13696, -32.18609, 
        -32.23525, -32.28462, -32.33438, -32.38452, -32.43489, -32.48527, 
        -32.53426, -32.58348, -32.63186, -32.67956, -32.72694, -32.77444, 
        -32.82222, -32.8703, -32.91878, -32.96775, -33.0176, -33.06815, 
        -33.11939, -33.17088, -33.22213, -33.27306, -33.32244, -33.37251, 
        -33.42234, -33.47164, -33.5204, -33.56846, -33.6158, -33.66258, 
        -33.70892, -33.75517, -33.80107, -33.84639, -33.89092, -33.93446, 
        -33.97709, -34.01927, -34.06134, -34.10365, -34.14537, -34.18842, 
        -34.23167, -34.27475, -34.31717, -34.35838, -34.39808, -34.43597, 
        -34.4721, -34.50681, -34.54058, -34.57363, -34.60623, -34.63858, 
        -34.67082, -34.70293, -34.73476, -34.76594, -34.79629, -34.82442, 
        -34.85239, -34.87918, -34.90488, -34.92945, -34.95319, -34.97696, 
        -35.00063, -35.02475, -35.04927, -35.07379, -35.09819, -35.1224, 
        -35.14642, -35.17054, -35.19474, -35.21922, -35.24391, -35.26881, 
        -35.29387, -35.31858, -35.34519, -35.37301, -35.40139, -35.42989, 
        -35.45768, -35.48452, -35.5104, -35.5357, -35.56057, -35.58554, 
        -35.61099, -35.63692, -35.66315, -35.68935, -35.71529, -35.74072, 
        -35.76558, -35.79009, -35.81435, -35.83849, -35.86274, -35.88614, 
        -35.91073, -35.93542, -35.95996, -35.9839, -36.00679, -36.02815, 
        -36.04796, -36.0666, -36.08475, -36.10301, -36.12169, -36.1412, 
        -36.16139, -36.1821, -36.2028, -36.22319, -36.24324, -36.26285, 
        -36.28206, -36.30107, -36.3198, -36.33817, -36.3557, -36.37434, 
        -36.39361, -36.41363, -36.43427, -36.45529, -36.47564, -36.49507, 
        -36.51336, -36.5306, -36.54756, -36.56513, -36.58373, -36.60398, 
        -36.62671, -36.65228, -36.68158, -36.71471, -36.75165, -36.79221, 
        -36.83609, -36.88317, -36.93277, -36.98436, -37.03747, -37.09167, 
        -37.14626, -37.19935, -37.25195, -37.30178, -37.34826, -37.39222, 
        -37.43333, -37.47307, -37.51223, -37.55124, -37.59043, -37.62981, 
        -37.6688, -37.70666, -37.74262, -37.77615, -37.807, -37.83519, 
        -37.86118, -37.88543, -37.90881, -37.93249, -37.95683, -37.98259, 
        -38.00935, -38.03656, -38.06352, -38.08979, -38.11518, -38.13977, 
        -38.16372, -38.18619, -38.20932, -38.23198, -38.25411, -38.27511, 
        -38.2947, -38.31255, -38.32788, -38.34082, -38.35174, -38.36127, 
        -38.37003, -38.37829, -38.38607, -38.39358, -38.40078, -38.40764, 
        -38.41386, -38.4191, -38.4232, -38.42625, -38.429, -38.43153, 
        -38.4345, -38.43798, -38.44159, -38.44526, -38.44905, -38.45222, 
        -38.45435, -38.45511, -38.45423, -38.45178, -38.44737, -38.44128, 
        -38.43364, -38.42498, -38.4157, -38.40524, -38.39598, -38.38712, 
        -38.37887, -38.37086, -38.36226, -38.35188, -38.33858, -38.32173, 
        -38.30072, -38.27546, -38.24566, -38.21158, -38.17305, -38.12906, 
        -38.07776, -38.0167, -37.9435, -37.85538, -37.75131, -37.63148, 
        -37.49987, -37.36179, -37.22591, -37.10191, -36.99947, -36.92705, 
        -36.8903,
  -29.55062, -29.59746, -29.64476, -29.69206, -29.73943, -29.78658, 
        -29.83355, -29.88062, -29.92822, -29.97582, -30.02565, -30.07648, 
        -30.12811, -30.18024, -30.23249, -30.28502, -30.33782, -30.39061, 
        -30.44312, -30.49513, -30.54654, -30.59718, -30.64719, -30.69576, 
        -30.74518, -30.79452, -30.84377, -30.89278, -30.94141, -30.98971, 
        -31.03805, -31.0865, -31.13522, -31.18401, -31.23304, -31.28249, 
        -31.33199, -31.38104, -31.42962, -31.47649, -31.52403, -31.5716, 
        -31.61946, -31.66759, -31.71602, -31.76441, -31.81288, -31.8615, 
        -31.91038, -31.95944, -32.00863, -32.05796, -32.10722, -32.15658, 
        -32.20492, -32.25441, -32.30408, -32.35407, -32.40419, -32.45422, 
        -32.50383, -32.55277, -32.60094, -32.64856, -32.69597, -32.74359, 
        -32.79158, -32.83989, -32.88862, -32.93773, -32.98726, -33.03634, 
        -33.08691, -33.13772, -33.18848, -33.23891, -33.28917, -33.33906, 
        -33.38879, -33.43822, -33.48712, -33.53544, -33.58316, -33.63017, 
        -33.67674, -33.72294, -33.76876, -33.81385, -33.8572, -33.9007, 
        -33.9435, -33.98589, -34.02819, -34.07074, -34.1137, -34.15705, 
        -34.20063, -34.24406, -34.28675, -34.32809, -34.3677, -34.40525, 
        -34.44083, -34.47492, -34.50797, -34.54043, -34.57259, -34.6036, 
        -34.6356, -34.66759, -34.6993, -34.73039, -34.76059, -34.78971, 
        -34.81771, -34.84457, -34.87028, -34.89494, -34.91893, -34.9423, 
        -34.96545, -34.98895, -35.01271, -35.03652, -35.06023, -35.08368, 
        -35.10722, -35.12967, -35.15343, -35.17742, -35.2016, -35.22625, 
        -35.25117, -35.27674, -35.30318, -35.3307, -35.35895, -35.38701, 
        -35.41435, -35.4407, -35.46606, -35.49083, -35.51527, -35.53972, 
        -35.56451, -35.58978, -35.61531, -35.64099, -35.66547, -35.69064, 
        -35.7153, -35.73979, -35.76401, -35.78802, -35.81245, -35.8369, 
        -35.86151, -35.88607, -35.91061, -35.93455, -35.9573, -35.97847, 
        -35.99809, -36.01657, -36.03475, -36.05313, -36.07211, -36.09195, 
        -36.11253, -36.13341, -36.15419, -36.17355, -36.19336, -36.2128, 
        -36.23194, -36.25059, -36.26927, -36.28768, -36.30577, -36.32409, 
        -36.34307, -36.36299, -36.38374, -36.40485, -36.42549, -36.44527, 
        -36.46387, -36.48166, -36.49924, -36.51736, -36.53674, -36.55784, 
        -36.5815, -36.60825, -36.63869, -36.67308, -36.71036, -36.75235, 
        -36.79782, -36.84629, -36.89742, -36.95057, -37.00488, -37.0599, 
        -37.11504, -37.16946, -37.22215, -37.2717, -37.31802, -37.36134, 
        -37.40191, -37.44122, -37.47998, -37.51884, -37.55801, -37.5973, 
        -37.63606, -37.67355, -37.70903, -37.74201, -37.77227, -37.79988, 
        -37.8252, -37.84892, -37.87197, -37.89392, -37.91771, -37.94274, 
        -37.96852, -37.99491, -38.02131, -38.04712, -38.0723, -38.09692, 
        -38.12118, -38.14516, -38.16885, -38.19203, -38.21437, -38.23545, 
        -38.25488, -38.27206, -38.28688, -38.29927, -38.30974, -38.31911, 
        -38.32794, -38.33636, -38.34413, -38.35127, -38.35807, -38.36446, 
        -38.36984, -38.37431, -38.37769, -38.38018, -38.38224, -38.38439, 
        -38.38698, -38.39016, -38.39264, -38.39651, -38.40053, -38.40406, 
        -38.40662, -38.40767, -38.40705, -38.40464, -38.40016, -38.39399, 
        -38.38617, -38.37733, -38.368, -38.35865, -38.34971, -38.34138, 
        -38.33372, -38.32642, -38.3185, -38.30899, -38.29668, -38.28069, 
        -38.26048, -38.23566, -38.20631, -38.17247, -38.13393, -38.08983, 
        -38.03857, -37.97782, -37.90529, -37.81832, -37.71561, -37.59747, 
        -37.46738, -37.3304, -37.19458, -37.0698, -36.96571, -36.89093, 
        -36.85139,
  -29.53134, -29.57833, -29.62582, -29.67357, -29.72023, -29.76758, 
        -29.81461, -29.8617, -29.90937, -29.95806, -30.00795, -30.05876, 
        -30.11008, -30.16166, -30.21326, -30.26499, -30.31703, -30.3693, 
        -30.42148, -30.47234, -30.52367, -30.57425, -30.62411, -30.6732, 
        -30.72203, -30.77078, -30.81912, -30.86734, -30.91518, -30.96268, 
        -31.01014, -31.0579, -31.10614, -31.15462, -31.20265, -31.25219, 
        -31.30171, -31.35097, -31.39967, -31.44748, -31.49478, -31.54187, 
        -31.58922, -31.63682, -31.68463, -31.73289, -31.78144, -31.8304, 
        -31.87976, -31.92834, -31.97788, -32.02739, -32.07694, -32.12645, 
        -32.17605, -32.22563, -32.27533, -32.3251, -32.37483, -32.42429, 
        -32.47325, -32.52167, -32.56953, -32.61727, -32.66489, -32.7128, 
        -32.76011, -32.80864, -32.85766, -32.90693, -32.9565, -33.0063, 
        -33.05645, -33.10691, -33.15739, -33.20769, -33.25795, -33.30788, 
        -33.35762, -33.40679, -33.45572, -33.50406, -33.55191, -33.59828, 
        -33.64485, -33.6908, -33.7361, -33.78071, -33.82468, -33.86804, 
        -33.91095, -33.95369, -33.99636, -34.0394, -34.08285, -34.12662, 
        -34.17054, -34.21419, -34.25705, -34.2985, -34.33804, -34.37443, 
        -34.40977, -34.44343, -34.47589, -34.50778, -34.53934, -34.57084, 
        -34.60245, -34.63409, -34.66552, -34.69638, -34.72641, -34.75542, 
        -34.78344, -34.81042, -34.83635, -34.8612, -34.88498, -34.90801, 
        -34.92963, -34.95237, -34.97519, -34.99816, -35.02122, -35.04421, 
        -35.0672, -35.09026, -35.11351, -35.13698, -35.16079, -35.18515, 
        -35.20989, -35.23557, -35.26198, -35.28919, -35.31697, -35.34466, 
        -35.37136, -35.39722, -35.42201, -35.44516, -35.46889, -35.49267, 
        -35.51667, -35.54104, -35.5658, -35.59089, -35.616, -35.64096, 
        -35.6656, -35.69016, -35.71448, -35.73877, -35.7632, -35.78781, 
        -35.81263, -35.83719, -35.86148, -35.88533, -35.90774, -35.92864, 
        -35.94812, -35.96565, -35.98401, -36.00274, -36.02214, -36.0424, 
        -36.06327, -36.08436, -36.10525, -36.12563, -36.14541, -36.16466, 
        -36.18364, -36.20222, -36.22064, -36.23877, -36.25656, -36.27465, 
        -36.29344, -36.31318, -36.33391, -36.35508, -36.37601, -36.3961, 
        -36.41513, -36.43348, -36.4507, -36.46958, -36.48966, -36.51177, 
        -36.53654, -36.56456, -36.59631, -36.632, -36.67152, -36.71473, 
        -36.76164, -36.81141, -36.86378, -36.9179, -36.97321, -37.029, 
        -37.08455, -37.13922, -37.1918, -37.2413, -37.28746, -37.33013, 
        -37.37041, -37.40923, -37.44768, -37.48637, -37.52551, -37.56458, 
        -37.60215, -37.63933, -37.67442, -37.70704, -37.73689, -37.76402, 
        -37.78884, -37.81205, -37.83461, -37.85712, -37.88013, -37.9042, 
        -37.92923, -37.95458, -37.98017, -38.00546, -38.03046, -38.05521, 
        -38.0799, -38.10443, -38.12873, -38.15243, -38.17483, -38.19554, 
        -38.21439, -38.23108, -38.24528, -38.25721, -38.26743, -38.2768, 
        -38.28571, -38.29411, -38.30101, -38.30782, -38.31425, -38.31993, 
        -38.32442, -38.32801, -38.33076, -38.33276, -38.33442, -38.33635, 
        -38.33881, -38.3418, -38.34526, -38.34904, -38.35302, -38.3566, 
        -38.35925, -38.36048, -38.35982, -38.35746, -38.35299, -38.34681, 
        -38.33909, -38.33021, -38.32091, -38.31166, -38.30288, -38.29475, 
        -38.28732, -38.28019, -38.27259, -38.26367, -38.25213, -38.23699, 
        -38.2177, -38.19366, -38.16502, -38.13169, -38.09344, -38.04962, 
        -37.99866, -37.93856, -37.86594, -37.78053, -37.68011, -37.56483, 
        -37.43723, -37.30293, -37.16905, -37.04496, -36.94046, -36.86407, 
        -36.82131,
  -29.51248, -29.55956, -29.607, -29.65463, -29.70217, -29.7494, 
        -29.79642, -29.84361, -29.89151, -29.94047, -29.9905, -30.0413, 
        -30.09245, -30.14364, -30.19374, -30.24493, -30.29636, -30.34804, 
        -30.39976, -30.45129, -30.50242, -30.55291, -30.60264, -30.65158, 
        -30.69991, -30.74782, -30.79532, -30.84243, -30.88915, -30.93468, 
        -30.98139, -31.02861, -31.07652, -31.12514, -31.17439, -31.22407, 
        -31.27378, -31.32309, -31.3716, -31.41919, -31.46608, -31.51272, 
        -31.55951, -31.60662, -31.65316, -31.70121, -31.74985, -31.79904, 
        -31.84864, -31.89843, -31.94819, -31.9979, -32.04764, -32.09744, 
        -32.14726, -32.19703, -32.2467, -32.2962, -32.34539, -32.3941, 
        -32.4413, -32.48913, -32.53679, -32.58455, -32.63255, -32.68089, 
        -32.72962, -32.77868, -32.82797, -32.8773, -32.92685, -32.97649, 
        -33.02646, -33.07679, -33.12732, -33.1778, -33.22804, -33.27697, 
        -33.32655, -33.37576, -33.4246, -33.47301, -33.52095, -33.5683, 
        -33.61491, -33.66066, -33.70553, -33.74961, -33.79309, -33.83617, 
        -33.87907, -33.92201, -33.96519, -34.00878, -34.05276, -34.096, 
        -34.14025, -34.18409, -34.22707, -34.26859, -34.30817, -34.34553, 
        -34.3807, -34.41404, -34.44608, -34.47737, -34.50831, -34.53924, 
        -34.57031, -34.60145, -34.63246, -34.66291, -34.69255, -34.72129, 
        -34.74813, -34.77506, -34.80103, -34.82587, -34.84954, -34.87229, 
        -34.89447, -34.91652, -34.93863, -34.9609, -34.98333, -35.00586, 
        -35.02847, -35.05117, -35.07404, -35.09717, -35.12074, -35.14487, 
        -35.16967, -35.19526, -35.22066, -35.24776, -35.27516, -35.30221, 
        -35.32833, -35.35332, -35.37726, -35.40043, -35.42318, -35.44584, 
        -35.46873, -35.49209, -35.51606, -35.54062, -35.56556, -35.59059, 
        -35.61553, -35.64035, -35.66507, -35.68977, -35.71454, -35.73939, 
        -35.76319, -35.78772, -35.81175, -35.83496, -35.85697, -35.87761, 
        -35.89703, -35.91575, -35.93442, -35.95356, -35.97343, -35.99402, 
        -36.01512, -36.03635, -36.05732, -36.07775, -36.09754, -36.11677, 
        -36.13564, -36.15422, -36.17249, -36.19041, -36.20811, -36.22603, 
        -36.24365, -36.26336, -36.28407, -36.30526, -36.32629, -36.34661, 
        -36.36606, -36.38494, -36.4038, -36.42338, -36.44439, -36.46755, 
        -36.49356, -36.52296, -36.5561, -36.59325, -36.63418, -36.67873, 
        -36.72667, -36.77759, -36.83091, -36.88588, -36.94173, -36.99779, 
        -37.05341, -37.10781, -37.15903, -37.20821, -37.25405, -37.29662, 
        -37.33677, -37.3756, -37.41412, -37.45293, -37.49202, -37.53111, 
        -37.56943, -37.60631, -37.64112, -37.67338, -37.70282, -37.72948, 
        -37.75381, -37.77651, -37.79845, -37.82034, -37.84273, -37.86592, 
        -37.8899, -37.91444, -37.93925, -37.9641, -37.98895, -38.01387, 
        -38.03889, -38.0639, -38.08854, -38.11127, -38.13353, -38.15393, 
        -38.17228, -38.18847, -38.20237, -38.21415, -38.22434, -38.2336, 
        -38.24235, -38.2506, -38.25815, -38.26479, -38.27051, -38.27532, 
        -38.27915, -38.28211, -38.28432, -38.28604, -38.28764, -38.28954, 
        -38.29197, -38.29495, -38.29836, -38.30206, -38.30583, -38.30925, 
        -38.31177, -38.3129, -38.31234, -38.30997, -38.30574, -38.29969, 
        -38.29206, -38.28328, -38.27393, -38.26462, -38.25576, -38.24659, 
        -38.23907, -38.23186, -38.22437, -38.21558, -38.20467, -38.19036, 
        -38.1719, -38.14888, -38.12113, -38.0886, -38.05109, -38.00787, 
        -37.95763, -37.89849, -37.82831, -37.74503, -37.64745, -37.53576, 
        -37.41231, -37.28188, -37.15152, -37.02993, -36.9263, -36.84901, 
        -36.80358,
  -29.4961, -29.54301, -29.59016, -29.63736, -29.68443, -29.73128, 
        -29.77818, -29.82558, -29.87386, -29.92319, -29.97242, -30.02318, 
        -30.07408, -30.12496, -30.17571, -30.2266, -30.27757, -30.3287, 
        -30.37987, -30.43094, -30.48178, -30.53224, -30.582, -30.63095, 
        -30.67771, -30.7248, -30.77105, -30.81683, -30.86225, -30.90766, 
        -30.95369, -31.00059, -31.04858, -31.09772, -31.14749, -31.19757, 
        -31.24738, -31.29653, -31.34464, -31.39066, -31.43692, -31.48292, 
        -31.52914, -31.57586, -31.6232, -31.67131, -31.72014, -31.76946, 
        -31.81902, -31.8688, -31.91855, -31.96827, -32.01812, -32.0681, 
        -32.11818, -32.16708, -32.21679, -32.26603, -32.31462, -32.36254, 
        -32.40995, -32.45722, -32.50467, -32.5527, -32.60116, -32.64998, 
        -32.6991, -32.74841, -32.79787, -32.84741, -32.89682, -32.94632, 
        -32.99522, -33.04565, -33.09647, -33.14738, -33.19785, -33.24794, 
        -33.29754, -33.34671, -33.39548, -33.44389, -33.4919, -33.53936, 
        -33.58602, -33.63171, -33.6763, -33.71987, -33.76284, -33.8045, 
        -33.84725, -33.89033, -33.93389, -33.97796, -34.02243, -34.06705, 
        -34.11154, -34.1555, -34.19851, -34.24007, -34.27976, -34.31725, 
        -34.35248, -34.38559, -34.41726, -34.44795, -34.47823, -34.50854, 
        -34.53801, -34.56861, -34.59903, -34.62898, -34.65806, -34.68639, 
        -34.71378, -34.74038, -34.76623, -34.79091, -34.81441, -34.83699, 
        -34.85884, -34.88043, -34.90197, -34.92364, -34.94557, -34.96767, 
        -34.98993, -35.01232, -35.03386, -35.05671, -35.07995, -35.10394, 
        -35.12873, -35.15434, -35.18067, -35.20755, -35.23443, -35.26091, 
        -35.28631, -35.31041, -35.33342, -35.35546, -35.37693, -35.3982, 
        -35.41976, -35.44199, -35.46508, -35.48921, -35.51411, -35.53838, 
        -35.56378, -35.58923, -35.61439, -35.63958, -35.66485, -35.69005, 
        -35.71498, -35.73928, -35.7628, -35.78534, -35.80672, -35.827, 
        -35.8465, -35.86542, -35.88447, -35.90404, -35.92427, -35.94511, 
        -35.96634, -35.98763, -36.00858, -36.02921, -36.04827, -36.0677, 
        -36.0867, -36.10538, -36.12357, -36.14148, -36.15908, -36.17708, 
        -36.19565, -36.21558, -36.23635, -36.25756, -36.27861, -36.29909, 
        -36.31889, -36.33826, -36.35774, -36.37799, -36.39979, -36.42389, 
        -36.45112, -36.48194, -36.51661, -36.55515, -36.59758, -36.6434, 
        -36.69149, -36.74327, -36.79729, -36.85271, -36.90881, -36.96484, 
        -37.0201, -37.07389, -37.12542, -37.17395, -37.21949, -37.26227, 
        -37.30272, -37.34202, -37.38107, -37.42028, -37.45969, -37.49873, 
        -37.53682, -37.57339, -37.60787, -37.63971, -37.66891, -37.6952, 
        -37.71911, -37.74137, -37.76281, -37.78416, -37.80588, -37.82721, 
        -37.85022, -37.87381, -37.89791, -37.92223, -37.94689, -37.97191, 
        -37.99714, -38.02231, -38.04696, -38.07042, -38.09223, -38.11206, 
        -38.1298, -38.14586, -38.15976, -38.17168, -38.182, -38.19124, 
        -38.19979, -38.20774, -38.21497, -38.22114, -38.22628, -38.23048, 
        -38.23355, -38.23602, -38.23786, -38.23952, -38.2412, -38.24323, 
        -38.24573, -38.2488, -38.25216, -38.25565, -38.25806, -38.26113, 
        -38.26335, -38.26431, -38.26377, -38.26163, -38.25767, -38.25194, 
        -38.24456, -38.2359, -38.22653, -38.21708, -38.20797, -38.1996, 
        -38.19178, -38.18427, -38.17655, -38.16779, -38.15705, -38.14331, 
        -38.12561, -38.10366, -38.07713, -38.04571, -38.00928, -37.96711, 
        -37.91796, -37.86021, -37.79183, -37.71104, -37.61687, -37.50946, 
        -37.39098, -37.26573, -37.14024, -37.02261, -36.92107, -36.84371, 
        -36.79635,
  -29.48055, -29.52744, -29.57437, -29.621, -29.66735, -29.71268, 
        -29.75942, -29.80697, -29.85562, -29.90533, -29.95571, -30.0065, 
        -30.0573, -30.10797, -30.15855, -30.20906, -30.2597, -30.3103, 
        -30.36086, -30.41137, -30.4608, -30.51108, -30.56076, -30.60939, 
        -30.65686, -30.70272, -30.74783, -30.7922, -30.83637, -30.88082, 
        -30.92631, -30.97323, -31.02173, -31.07158, -31.12215, -31.17195, 
        -31.22158, -31.27035, -31.31787, -31.36411, -31.4095, -31.45474, 
        -31.50035, -31.5467, -31.59392, -31.64204, -31.69102, -31.7402, 
        -31.78975, -31.83937, -31.888, -31.93767, -31.98751, -32.0376, 
        -32.08774, -32.13773, -32.18742, -32.23641, -32.28457, -32.33192, 
        -32.3787, -32.42561, -32.47305, -32.52129, -32.57019, -32.61943, 
        -32.6689, -32.7174, -32.76686, -32.81617, -32.86533, -32.9146, 
        -32.96432, -33.01495, -33.06612, -33.11745, -33.16846, -33.2189, 
        -33.26872, -33.31804, -33.36687, -33.41542, -33.4636, -33.51121, 
        -33.55716, -33.60292, -33.64742, -33.69072, -33.73333, -33.77554, 
        -33.81802, -33.86107, -33.90482, -33.94917, -33.99389, -34.03869, 
        -34.08324, -34.1272, -34.17015, -34.21166, -34.25138, -34.28896, 
        -34.32326, -34.3564, -34.38781, -34.41808, -34.44776, -34.47749, 
        -34.50758, -34.53763, -34.56753, -34.5969, -34.62545, -34.65314, 
        -34.67998, -34.70594, -34.73123, -34.75521, -34.77863, -34.8012, 
        -34.82291, -34.84322, -34.86443, -34.88574, -34.90722, -34.9289, 
        -34.95076, -34.97276, -34.99483, -35.01733, -35.04032, -35.06413, 
        -35.08893, -35.1145, -35.14073, -35.16728, -35.19363, -35.21936, 
        -35.24399, -35.26722, -35.2892, -35.31011, -35.32915, -35.34895, 
        -35.36908, -35.39004, -35.4123, -35.43598, -35.46088, -35.48652, 
        -35.51248, -35.53857, -35.56443, -35.5901, -35.61591, -35.64149, 
        -35.66647, -35.6905, -35.71348, -35.73529, -35.75612, -35.77609, 
        -35.79539, -35.81451, -35.8329, -35.85282, -35.87336, -35.89441, 
        -35.9157, -35.93705, -35.95815, -35.9788, -35.9992, -36.01914, 
        -36.0385, -36.05734, -36.0756, -36.09365, -36.11155, -36.12981, 
        -36.14888, -36.16896, -36.18994, -36.21123, -36.2323, -36.25281, 
        -36.27279, -36.29251, -36.31251, -36.33229, -36.35471, -36.37971, 
        -36.40796, -36.44016, -36.47631, -36.51637, -36.56021, -36.60744, 
        -36.65759, -36.71015, -36.76456, -36.8201, -36.87608, -36.93169, 
        -36.98624, -37.03901, -37.08977, -37.13784, -37.18324, -37.2262, 
        -37.26723, -37.30765, -37.34768, -37.38771, -37.42754, -37.4667, 
        -37.50464, -37.53984, -37.57393, -37.60545, -37.63424, -37.66002, 
        -37.68364, -37.7055, -37.72642, -37.74723, -37.76826, -37.78972, 
        -37.81176, -37.83445, -37.85775, -37.88165, -37.90609, -37.93108, 
        -37.95633, -37.98134, -38.00563, -38.02852, -38.04953, -38.06883, 
        -38.08657, -38.10236, -38.11655, -38.12895, -38.13952, -38.14877, 
        -38.15709, -38.16464, -38.17134, -38.17705, -38.18058, -38.18398, 
        -38.18665, -38.18871, -38.19044, -38.19221, -38.19418, -38.19644, 
        -38.19914, -38.20219, -38.20546, -38.20873, -38.21175, -38.21433, 
        -38.21614, -38.2169, -38.21638, -38.21444, -38.21099, -38.20565, 
        -38.19864, -38.19016, -38.18076, -38.17126, -38.16203, -38.15332, 
        -38.14525, -38.13741, -38.12933, -38.12032, -38.10957, -38.09618, 
        -38.0793, -38.05832, -38.03297, -38.00291, -37.96781, -37.92704, 
        -37.87928, -37.8233, -37.75705, -37.67937, -37.58814, -37.48561, 
        -37.37289, -37.25385, -37.13434, -37.02164, -36.92341, -36.84689, 
        -36.79795,
  -29.46536, -29.51132, -29.55783, -29.60394, -29.64982, -29.69582, 
        -29.74244, -29.79012, -29.83903, -29.889, -29.93964, -29.99052, 
        -30.04134, -30.09196, -30.14237, -30.19165, -30.24182, -30.29186, 
        -30.34176, -30.39164, -30.4416, -30.49149, -30.54078, -30.58886, 
        -30.63536, -30.68032, -30.72414, -30.76731, -30.81044, -30.85425, 
        -30.8985, -30.94572, -30.99497, -31.04575, -31.09714, -31.14818, 
        -31.19804, -31.24635, -31.29305, -31.33836, -31.38286, -31.42728, 
        -31.47227, -31.51825, -31.56536, -31.6125, -31.66138, -31.71062, 
        -31.76, -31.80939, -31.85881, -31.90837, -31.95815, -32.00814, 
        -32.05818, -32.1081, -32.15768, -32.20659, -32.25455, -32.3016, 
        -32.34816, -32.39388, -32.44134, -32.48973, -32.53888, -32.58841, 
        -32.63803, -32.68757, -32.73687, -32.78582, -32.83456, -32.88348, 
        -32.93307, -32.98378, -33.03527, -33.08703, -33.13852, -33.18939, 
        -33.2386, -33.28825, -33.33747, -33.38633, -33.43485, -33.48288, 
        -33.5301, -33.57612, -33.62074, -33.66402, -33.70637, -33.74834, 
        -33.79053, -33.83342, -33.87716, -33.92155, -33.96629, -34.01102, 
        -34.05444, -34.0982, -34.14093, -34.18224, -34.22183, -34.2594, 
        -34.2948, -34.32803, -34.35938, -34.38942, -34.41886, -34.4483, 
        -34.47796, -34.50769, -34.53714, -34.56596, -34.59395, -34.62099, 
        -34.64713, -34.67135, -34.69569, -34.71918, -34.74195, -34.76411, 
        -34.78575, -34.80708, -34.82822, -34.8493, -34.87041, -34.89162, 
        -34.91296, -34.93439, -34.95596, -34.97791, -35.00058, -35.02423, 
        -35.0489, -35.07439, -35.10035, -35.1254, -35.15105, -35.17598, 
        -35.19984, -35.22235, -35.24345, -35.26325, -35.2821, -35.30056, 
        -35.31932, -35.33907, -35.36041, -35.3836, -35.40847, -35.43429, 
        -35.46064, -35.48712, -35.51357, -35.53996, -35.56625, -35.59212, 
        -35.61709, -35.63983, -35.66227, -35.68353, -35.70385, -35.72346, 
        -35.74271, -35.76197, -35.7816, -35.8018, -35.82257, -35.84378, 
        -35.86523, -35.88673, -35.90804, -35.92906, -35.94975, -35.97004, 
        -35.98982, -36.00899, -36.02755, -36.04581, -36.06418, -36.08309, 
        -36.10286, -36.12251, -36.14374, -36.1651, -36.18613, -36.20663, 
        -36.22669, -36.24663, -36.26692, -36.28816, -36.3112, -36.33696, 
        -36.36623, -36.39955, -36.43703, -36.47857, -36.5238, -36.57227, 
        -36.62345, -36.6767, -36.73138, -36.78685, -36.84241, -36.89734, 
        -36.95095, -37.00279, -37.05257, -37.10016, -37.14459, -37.18815, 
        -37.23037, -37.27188, -37.31309, -37.35407, -37.39451, -37.43394, 
        -37.47189, -37.50792, -37.54163, -37.57268, -37.60088, -37.6263, 
        -37.6494, -37.67088, -37.69139, -37.71155, -37.73169, -37.7523, 
        -37.77342, -37.79526, -37.8179, -37.84137, -37.8656, -37.89043, 
        -37.91542, -37.93999, -37.96354, -37.98562, -38.00604, -38.02394, 
        -38.04148, -38.05763, -38.07221, -38.08493, -38.09579, -38.10506, 
        -38.11314, -38.12027, -38.12645, -38.13154, -38.13546, -38.13829, 
        -38.14043, -38.14224, -38.14405, -38.14604, -38.14829, -38.15084, 
        -38.15373, -38.15685, -38.15999, -38.16297, -38.1656, -38.1677, 
        -38.1691, -38.16959, -38.16905, -38.16734, -38.16427, -38.15953, 
        -38.15303, -38.14492, -38.13577, -38.12626, -38.117, -38.10829, 
        -38.10003, -38.09096, -38.08253, -38.07318, -38.06223, -38.04895, 
        -38.03256, -38.01247, -37.98829, -37.95965, -37.9261, -37.88691, 
        -37.84101, -37.78707, -37.72358, -37.64929, -37.56352, -37.46663, 
        -37.3604, -37.24839, -37.13575, -37.0289, -36.93472, -36.8596, 
        -36.80874,
  -29.44917, -29.4961, -29.54244, -29.58824, -29.63382, -29.67965, 
        -29.7263, -29.77415, -29.82327, -29.87341, -29.9232, -29.97425, 
        -30.02522, -30.07589, -30.12619, -30.17617, -30.22586, -30.27526, 
        -30.32449, -30.37375, -30.42316, -30.47244, -30.52098, -30.56815, 
        -30.61356, -30.65635, -30.69901, -30.74112, -30.78351, -30.82703, 
        -30.87244, -30.92023, -30.97031, -31.02207, -31.07425, -31.12566, 
        -31.17543, -31.22321, -31.26908, -31.3135, -31.35605, -31.39976, 
        -31.44412, -31.4897, -31.53661, -31.58484, -31.63373, -31.68288, 
        -31.73209, -31.78131, -31.8306, -31.88, -31.92953, -31.97913, 
        -32.02879, -32.07845, -32.12692, -32.17587, -32.22392, -32.27106, 
        -32.31767, -32.36442, -32.4119, -32.46031, -32.5095, -32.55911, 
        -32.60873, -32.65827, -32.70724, -32.75566, -32.80385, -32.85235, 
        -32.90179, -32.95147, -33.00314, -33.05519, -33.10703, -33.15831, 
        -33.209, -33.25918, -33.30894, -33.35838, -33.40739, -33.45586, 
        -33.5035, -33.54992, -33.59488, -33.63837, -33.68086, -33.72274, 
        -33.76365, -33.80637, -33.84992, -33.89418, -33.93878, -33.9833, 
        -34.0274, -34.07075, -34.11301, -34.15393, -34.19324, -34.23068, 
        -34.26617, -34.29956, -34.33102, -34.36108, -34.39047, -34.41978, 
        -34.44925, -34.47778, -34.50691, -34.53538, -34.5629, -34.58936, 
        -34.6147, -34.63893, -34.66204, -34.68445, -34.70647, -34.72844, 
        -34.74993, -34.77152, -34.79271, -34.81377, -34.83458, -34.85532, 
        -34.87609, -34.89673, -34.9175, -34.93773, -34.95987, -34.98317, 
        -35.00758, -35.03276, -35.0582, -35.08342, -35.10826, -35.13232, 
        -35.15541, -35.17718, -35.19764, -35.2168, -35.23476, -35.25225, 
        -35.26996, -35.2887, -35.30919, -35.33176, -35.35624, -35.38204, 
        -35.40738, -35.43409, -35.46108, -35.48792, -35.51441, -35.54038, 
        -35.56529, -35.58875, -35.61084, -35.63177, -35.6518, -35.67124, 
        -35.69048, -35.70994, -35.72984, -35.75028, -35.77121, -35.79252, 
        -35.81414, -35.83583, -35.85742, -35.87877, -35.89985, -35.9196, 
        -35.93982, -35.95933, -35.9782, -35.99683, -36.01585, -36.03569, 
        -36.05642, -36.07778, -36.09931, -36.12075, -36.14169, -36.16213, 
        -36.18225, -36.20235, -36.2229, -36.24456, -36.26817, -36.29468, 
        -36.32483, -36.35914, -36.39773, -36.44061, -36.4871, -36.5367, 
        -36.58888, -36.6418, -36.69676, -36.75205, -36.80711, -36.8612, 
        -36.91382, -36.9647, -37.01377, -37.06115, -37.10668, -37.15096, 
        -37.19427, -37.23693, -37.27923, -37.32107, -37.36213, -37.40198, 
        -37.44015, -37.47612, -37.50952, -37.54002, -37.56768, -37.59261, 
        -37.61523, -37.63637, -37.65644, -37.67593, -37.6953, -37.71495, 
        -37.73423, -37.75537, -37.7775, -37.80062, -37.82461, -37.84911, 
        -37.87356, -37.89732, -37.9199, -37.94116, -37.96084, -37.97944, 
        -37.997, -38.01341, -38.02836, -38.04143, -38.05252, -38.06182, 
        -38.06972, -38.07652, -38.08229, -38.08684, -38.09021, -38.09249, 
        -38.0942, -38.09585, -38.09764, -38.09976, -38.10221, -38.1049, 
        -38.10786, -38.1109, -38.11395, -38.11674, -38.11915, -38.12094, 
        -38.12104, -38.12133, -38.12073, -38.11916, -38.11647, -38.11232, 
        -38.10644, -38.09891, -38.09025, -38.08095, -38.07191, -38.06348, 
        -38.05527, -38.04716, -38.03853, -38.02888, -38.01753, -38.00426, 
        -37.98807, -37.96851, -37.94532, -37.91809, -37.88622, -37.84896, 
        -37.8052, -37.75379, -37.69348, -37.62318, -37.54238, -37.45152, 
        -37.35234, -37.24799, -37.14292, -37.04242, -36.95313, -36.87997, 
        -36.82768,
  -29.43397, -29.4805, -29.52666, -29.57231, -29.61785, -29.66381, 
        -29.70971, -29.75787, -29.80723, -29.8576, -29.90858, -29.95979, 
        -30.01087, -30.06155, -30.11169, -30.16132, -30.21051, -30.25941, 
        -30.3081, -30.35676, -30.40448, -30.45283, -30.50026, -30.54613, 
        -30.59029, -30.63298, -30.67464, -30.71608, -30.75809, -30.80162, 
        -30.84732, -30.89564, -30.94641, -30.9987, -31.0514, -31.10196, 
        -31.15159, -31.19894, -31.24419, -31.28799, -31.33086, -31.37386, 
        -31.41781, -31.4629, -31.50962, -31.55771, -31.60651, -31.6557, 
        -31.70497, -31.75424, -31.80352, -31.85169, -31.90091, -31.95009, 
        -31.99933, -32.04859, -32.09785, -32.1468, -32.19495, -32.24229, 
        -32.28906, -32.33591, -32.38338, -32.4317, -32.48071, -32.53019, 
        -32.57986, -32.62803, -32.67677, -32.72458, -32.77255, -32.82064, 
        -32.86989, -32.92047, -32.9721, -33.0243, -33.07639, -33.12809, 
        -33.17939, -33.23026, -33.2806, -33.33061, -33.38023, -33.42924, 
        -33.47722, -33.52299, -33.56831, -33.61217, -33.65495, -33.69705, 
        -33.73904, -33.78162, -33.82502, -33.86913, -33.91355, -33.95782, 
        -34.00153, -34.04439, -34.08611, -34.12649, -34.16543, -34.20273, 
        -34.23826, -34.2708, -34.30246, -34.33274, -34.36232, -34.39162, 
        -34.42101, -34.45032, -34.47921, -34.50732, -34.53441, -34.5603, 
        -34.58491, -34.6083, -34.63044, -34.65196, -34.67337, -34.69469, 
        -34.71608, -34.73727, -34.75739, -34.7782, -34.79866, -34.81877, 
        -34.83876, -34.85853, -34.87844, -34.8989, -34.92038, -34.94299, 
        -34.96681, -34.99131, -35.01594, -35.04036, -35.06427, -35.08751, 
        -35.10983, -35.1311, -35.15115, -35.16984, -35.18742, -35.20339, 
        -35.22037, -35.23826, -35.25794, -35.27962, -35.30326, -35.3285, 
        -35.35458, -35.38108, -35.40794, -35.435, -35.46185, -35.48779, 
        -35.51255, -35.53595, -35.55801, -35.57896, -35.59903, -35.61861, 
        -35.63807, -35.65774, -35.67791, -35.6985, -35.71866, -35.74013, 
        -35.76201, -35.78406, -35.80606, -35.82782, -35.84932, -35.8705, 
        -35.89119, -35.91108, -35.93038, -35.9495, -35.96917, -35.98979, 
        -36.01123, -36.03307, -36.05497, -36.07634, -36.09719, -36.11757, 
        -36.13779, -36.15813, -36.17906, -36.20123, -36.22437, -36.25164, 
        -36.28273, -36.31796, -36.3575, -36.40134, -36.44893, -36.49954, 
        -36.5526, -36.60726, -36.66259, -36.71796, -36.77262, -36.82611, 
        -36.87807, -36.92837, -36.97708, -37.02425, -37.07011, -37.11488, 
        -37.15878, -37.20214, -37.24506, -37.28745, -37.32893, -37.36916, 
        -37.40763, -37.44379, -37.47712, -37.50636, -37.53363, -37.55828, 
        -37.58066, -37.6016, -37.62119, -37.63995, -37.65864, -37.67747, 
        -37.69699, -37.71755, -37.73926, -37.76206, -37.78566, -37.80965, 
        -37.83344, -37.85633, -37.87803, -37.89836, -37.9175, -37.93568, 
        -37.95293, -37.96914, -37.98415, -37.99727, -38.0085, -38.0179, 
        -38.02571, -38.03233, -38.03762, -38.04169, -38.04456, -38.04637, 
        -38.04668, -38.04796, -38.04956, -38.05171, -38.05426, -38.05712, 
        -38.06012, -38.06322, -38.06647, -38.06907, -38.07139, -38.07293, 
        -38.0738, -38.07388, -38.07315, -38.07171, -38.06946, -38.06592, 
        -38.06091, -38.05438, -38.04654, -38.03808, -38.02941, -38.0211, 
        -38.01291, -38.00462, -37.99561, -37.98564, -37.97393, -37.96036, 
        -37.94438, -37.92517, -37.90292, -37.87704, -37.8468, -37.81144, 
        -37.76991, -37.72125, -37.66444, -37.59844, -37.52295, -37.43853, 
        -37.34666, -37.24915, -37.15184, -37.05834, -36.97402, -36.90318, 
        -36.85081,
  -29.41928, -29.46443, -29.51023, -29.55581, -29.6015, -29.64775, 
        -29.69501, -29.74345, -29.79301, -29.84348, -29.89451, -29.94575, 
        -29.99681, -30.04737, -30.09731, -30.14663, -30.19449, -30.24298, 
        -30.29123, -30.33932, -30.38717, -30.43441, -30.4805, -30.52504, 
        -30.56796, -30.60956, -30.65048, -30.69147, -30.73337, -30.77702, 
        -30.8231, -30.87094, -30.92222, -30.975, -31.0279, -31.07955, 
        -31.12899, -31.176, -31.22083, -31.26413, -31.30665, -31.34924, 
        -31.39272, -31.43746, -31.48395, -31.53189, -31.57976, -31.62905, 
        -31.67846, -31.72786, -31.77716, -31.82624, -31.87504, -31.92362, 
        -31.97219, -32.02093, -32.06984, -32.11866, -32.16694, -32.2145, 
        -32.26153, -32.30852, -32.35492, -32.403, -32.45175, -32.50096, 
        -32.55028, -32.59927, -32.64764, -32.69542, -32.743, -32.79096, 
        -32.84007, -32.89033, -32.94188, -32.9941, -33.04644, -33.09855, 
        -33.1503, -33.20071, -33.25174, -33.30237, -33.35249, -33.40188, 
        -33.45024, -33.49731, -33.54297, -33.58731, -33.63059, -33.67318, 
        -33.71559, -33.75835, -33.80177, -33.84577, -33.88998, -33.93393, 
        -33.97719, -34.01847, -34.0596, -34.09948, -34.13804, -34.17517, 
        -34.21068, -34.24437, -34.27631, -34.30688, -34.33667, -34.36609, 
        -34.3954, -34.42449, -34.45304, -34.48074, -34.50736, -34.53273, 
        -34.55674, -34.57941, -34.59995, -34.62077, -34.64137, -34.66206, 
        -34.6829, -34.70374, -34.72438, -34.74469, -34.7646, -34.7841, 
        -34.80324, -34.82216, -34.84118, -34.86076, -34.88132, -34.90308, 
        -34.92591, -34.94936, -34.97295, -34.99633, -35.01828, -35.04068, 
        -35.0624, -35.08323, -35.10298, -35.12155, -35.13903, -35.15578, 
        -35.17244, -35.18981, -35.20868, -35.22938, -35.25202, -35.27623, 
        -35.30151, -35.3275, -35.35406, -35.38097, -35.40775, -35.43381, 
        -35.45858, -35.48204, -35.50327, -35.52447, -35.54487, -35.5648, 
        -35.58462, -35.60466, -35.62508, -35.6459, -35.66713, -35.6888, 
        -35.71095, -35.73339, -35.75585, -35.77813, -35.8001, -35.8217, 
        -35.84276, -35.86309, -35.88282, -35.90245, -35.92269, -35.94389, 
        -35.96591, -35.98818, -36.00916, -36.03055, -36.05137, -36.07185, 
        -36.0923, -36.11303, -36.13447, -36.15723, -36.18213, -36.21013, 
        -36.24174, -36.27774, -36.31837, -36.3631, -36.41174, -36.46347, 
        -36.51742, -36.57269, -36.62844, -36.68393, -36.7385, -36.79174, 
        -36.84338, -36.89333, -36.94174, -36.98881, -37.03474, -37.07868, 
        -37.12285, -37.16645, -37.20958, -37.25212, -37.29383, -37.3343, 
        -37.37304, -37.40942, -37.44293, -37.47325, -37.50052, -37.52511, 
        -37.54751, -37.56816, -37.58742, -37.60574, -37.62367, -37.64181, 
        -37.66066, -37.68084, -37.70223, -37.7247, -37.74788, -37.77126, 
        -37.79423, -37.81625, -37.83704, -37.85657, -37.87498, -37.89247, 
        -37.90916, -37.92393, -37.93849, -37.95148, -37.9627, -37.97216, 
        -37.98004, -37.98648, -37.99152, -37.99519, -37.99756, -37.99891, 
        -37.99975, -38.00064, -38.002, -38.004, -38.00657, -38.00952, 
        -38.01268, -38.01591, -38.01904, -38.02182, -38.02407, -38.02565, 
        -38.02639, -38.02629, -38.02548, -38.02412, -38.02223, -38.01949, 
        -38.01549, -38.01004, -38.00327, -37.99569, -37.98776, -37.97977, 
        -37.97161, -37.96308, -37.95367, -37.9431, -37.93009, -37.91627, 
        -37.90024, -37.88167, -37.86027, -37.83559, -37.80693, -37.77344, 
        -37.73425, -37.68847, -37.63523, -37.57376, -37.50378, -37.42577, 
        -37.3412, -37.25248, -37.16288, -37.07626, -36.99691, -36.92904, 
        -36.87666,
  -29.4042, -29.44991, -29.49547, -29.54111, -29.58708, -29.63367, 
        -29.68132, -29.72992, -29.77938, -29.82973, -29.88058, -29.93067, 
        -29.98161, -30.03199, -30.08169, -30.13084, -30.17949, -30.22765, 
        -30.27558, -30.32318, -30.36998, -30.41592, -30.46046, -30.50359, 
        -30.54553, -30.58635, -30.6259, -30.66678, -30.70877, -30.75273, 
        -30.79912, -30.84833, -30.89986, -30.95283, -31.00579, -31.0575, 
        -31.10662, -31.15347, -31.19806, -31.2412, -31.28354, -31.32496, 
        -31.36819, -31.41281, -31.45914, -31.50697, -31.55589, -31.60532, 
        -31.65504, -31.70468, -31.75408, -31.80296, -31.8513, -31.89915, 
        -31.94687, -31.99482, -32.04321, -32.0907, -32.13899, -32.18677, 
        -32.23412, -32.28133, -32.32866, -32.37645, -32.4248, -32.47363, 
        -32.52272, -32.57162, -32.6199, -32.66761, -32.71552, -32.76319, 
        -32.81177, -32.86172, -32.91191, -32.96387, -33.0164, -33.06888, 
        -33.12114, -33.17316, -33.22476, -33.27592, -33.32645, -33.37615, 
        -33.42473, -33.472, -33.51803, -33.5629, -33.60699, -33.65048, 
        -33.69363, -33.73584, -33.77936, -33.82329, -33.86728, -33.91085, 
        -33.95362, -33.9953, -34.03585, -34.07528, -34.11349, -34.15046, 
        -34.18592, -34.21972, -34.2519, -34.28278, -34.3128, -34.3423, 
        -34.37151, -34.40027, -34.42735, -34.45457, -34.4807, -34.50555, 
        -34.52903, -34.55119, -34.57222, -34.59248, -34.61239, -34.63235, 
        -34.65245, -34.67263, -34.69268, -34.71239, -34.73175, -34.75055, 
        -34.7688, -34.7867, -34.8047, -34.82334, -34.84187, -34.86243, 
        -34.88411, -34.90619, -34.9285, -34.95085, -34.97292, -34.99455, 
        -35.01563, -35.03598, -35.05537, -35.07385, -35.09136, -35.10816, 
        -35.12477, -35.14191, -35.16024, -35.18016, -35.20167, -35.22467, 
        -35.24882, -35.2729, -35.29893, -35.32553, -35.35221, -35.37815, 
        -35.40302, -35.42667, -35.44926, -35.47089, -35.49182, -35.51229, 
        -35.53261, -35.55292, -35.57357, -35.59451, -35.61586, -35.63772, 
        -35.66014, -35.68298, -35.70593, -35.72871, -35.75115, -35.77318, 
        -35.79367, -35.81445, -35.83464, -35.85468, -35.87545, -35.89714, 
        -35.9196, -35.94208, -35.96401, -35.98539, -36.00618, -36.02684, 
        -36.04771, -36.069, -36.09132, -36.11494, -36.14071, -36.16934, 
        -36.20183, -36.23843, -36.27996, -36.32566, -36.37545, -36.42818, 
        -36.48296, -36.53881, -36.59405, -36.64978, -36.7045, -36.75783, 
        -36.80945, -36.85922, -36.90723, -36.95404, -36.99977, -37.04457, 
        -37.08862, -37.1321, -37.17488, -37.21719, -37.25879, -37.29933, 
        -37.33828, -37.37498, -37.40879, -37.43945, -37.46703, -37.49182, 
        -37.51434, -37.53496, -37.55394, -37.57185, -37.58931, -37.60696, 
        -37.62533, -37.64512, -37.66528, -37.68745, -37.71022, -37.73295, 
        -37.7551, -37.77621, -37.79612, -37.81491, -37.83258, -37.84917, 
        -37.86511, -37.87999, -37.89374, -37.90619, -37.91719, -37.92661, 
        -37.93446, -37.94079, -37.94548, -37.94892, -37.95095, -37.95189, 
        -37.95249, -37.95305, -37.95401, -37.9557, -37.95816, -37.96109, 
        -37.96439, -37.96772, -37.97099, -37.97402, -37.97647, -37.97822, 
        -37.97897, -37.97878, -37.97679, -37.97539, -37.97372, -37.97167, 
        -37.96871, -37.9645, -37.95903, -37.95257, -37.9455, -37.93796, 
        -37.93002, -37.92126, -37.91149, -37.90048, -37.88805, -37.87395, 
        -37.85793, -37.83985, -37.81929, -37.79581, -37.76857, -37.73686, 
        -37.6999, -37.657, -37.60737, -37.55033, -37.48579, -37.414, 
        -37.3364, -37.25513, -37.17291, -37.09283, -37.0188, -36.95414, 
        -36.90242,
  -29.39207, -29.43718, -29.48257, -29.52827, -29.57448, -29.62138, 
        -29.66904, -29.71649, -29.76567, -29.81545, -29.86567, -29.91633, 
        -29.96681, -30.01687, -30.06637, -30.11533, -30.16372, -30.21168, 
        -30.25921, -30.30618, -30.35211, -30.39578, -30.43908, -30.4812, 
        -30.52228, -30.56281, -30.60334, -30.64442, -30.68676, -30.73105, 
        -30.77781, -30.82721, -30.87884, -30.93175, -30.9846, -31.03609, 
        -31.08426, -31.13088, -31.17531, -31.21822, -31.26059, -31.30308, 
        -31.34634, -31.39099, -31.43736, -31.48531, -31.53434, -31.58412, 
        -31.634, -31.68388, -31.73326, -31.78186, -31.82859, -31.87555, 
        -31.92226, -31.96938, -32.01694, -32.06492, -32.11307, -32.161, 
        -32.20864, -32.25609, -32.30346, -32.35098, -32.39885, -32.44723, 
        -32.49591, -32.54465, -32.59209, -32.64018, -32.68821, -32.73611, 
        -32.78448, -32.83396, -32.88469, -32.93655, -32.98894, -33.04182, 
        -33.09452, -33.14695, -33.19898, -33.25045, -33.30133, -33.35121, 
        -33.39999, -33.44759, -33.49307, -33.53868, -33.58361, -33.62806, 
        -33.67211, -33.71597, -33.75986, -33.80379, -33.84756, -33.89074, 
        -33.93305, -33.97422, -34.01425, -34.0532, -34.09109, -34.12782, 
        -34.16322, -34.1971, -34.22842, -34.25957, -34.2898, -34.31939, 
        -34.34834, -34.37665, -34.40418, -34.43078, -34.45633, -34.48071, 
        -34.50377, -34.52559, -34.54626, -34.56606, -34.58536, -34.60439, 
        -34.6235, -34.64268, -34.66185, -34.67984, -34.69843, -34.71655, 
        -34.73404, -34.75116, -34.76852, -34.78618, -34.80458, -34.82381, 
        -34.84375, -34.86427, -34.88506, -34.90602, -34.92699, -34.94761, 
        -34.96805, -34.98801, -35.00729, -35.02571, -35.04328, -35.06021, 
        -35.07592, -35.09293, -35.11097, -35.13028, -35.15089, -35.17265, 
        -35.19568, -35.2198, -35.24505, -35.27119, -35.29747, -35.32333, 
        -35.34836, -35.37216, -35.39515, -35.41726, -35.43873, -35.45972, 
        -35.48043, -35.50109, -35.52182, -35.54292, -35.5644, -35.58545, 
        -35.6083, -35.63171, -35.65518, -35.67854, -35.70161, -35.72408, 
        -35.74602, -35.76713, -35.7878, -35.80817, -35.82918, -35.85123, 
        -35.8739, -35.89653, -35.91868, -35.94022, -35.96134, -35.98244, 
        -36.00386, -36.02606, -36.04911, -36.07367, -36.10023, -36.1297, 
        -36.16183, -36.19928, -36.24139, -36.28812, -36.33865, -36.39224, 
        -36.44784, -36.50449, -36.56131, -36.6176, -36.67271, -36.72617, 
        -36.77769, -36.82731, -36.87487, -36.92104, -36.96627, -37.01068, 
        -37.05437, -37.09744, -37.13993, -37.18185, -37.22315, -37.2636, 
        -37.30262, -37.33953, -37.37381, -37.40499, -37.43223, -37.45748, 
        -37.48039, -37.50121, -37.52024, -37.53796, -37.55503, -37.57212, 
        -37.59005, -37.60932, -37.63, -37.65177, -37.6741, -37.69621, 
        -37.71764, -37.73794, -37.75695, -37.77471, -37.79141, -37.80694, 
        -37.82166, -37.83552, -37.84846, -37.86039, -37.87111, -37.88051, 
        -37.88844, -37.89476, -37.89932, -37.90258, -37.90417, -37.905, 
        -37.90512, -37.90547, -37.90522, -37.90671, -37.90893, -37.91188, 
        -37.9153, -37.9189, -37.92244, -37.92575, -37.92841, -37.93018, 
        -37.93077, -37.93034, -37.92918, -37.92775, -37.92633, -37.92484, 
        -37.92291, -37.91999, -37.91586, -37.91065, -37.90445, -37.89749, 
        -37.88971, -37.88079, -37.87062, -37.85916, -37.84626, -37.83191, 
        -37.81601, -37.79842, -37.7788, -37.75653, -37.73081, -37.70082, 
        -37.66611, -37.62597, -37.57981, -37.52694, -37.46745, -37.40159, 
        -37.33039, -37.25578, -37.18021, -37.10519, -37.03628, -36.97479, 
        -36.92423,
  -29.3815, -29.4262, -29.47039, -29.51616, -29.56259, -29.60963, 
        -29.65719, -29.70516, -29.75348, -29.80234, -29.85165, -29.90133, 
        -29.95098, -30.00059, -30.04985, -30.09863, -30.14688, -30.19355, 
        -30.24058, -30.28684, -30.33187, -30.37566, -30.41798, -30.45947, 
        -30.50031, -30.54099, -30.58201, -30.62375, -30.66684, -30.71174, 
        -30.75867, -30.80709, -30.8585, -30.91103, -30.96333, -31.01449, 
        -31.06351, -31.11003, -31.15443, -31.19757, -31.24002, -31.28265, 
        -31.32612, -31.37096, -31.41752, -31.46568, -31.515, -31.56394, 
        -31.61421, -31.66413, -31.71344, -31.76171, -31.8087, -31.85472, 
        -31.90036, -31.94632, -31.99285, -32.04017, -32.08797, -32.13603, 
        -32.184, -32.23176, -32.27925, -32.3256, -32.37305, -32.42091, 
        -32.46919, -32.51779, -32.56648, -32.61498, -32.6633, -32.71158, 
        -32.75993, -32.80907, -32.85916, -32.91064, -32.96317, -33.01614, 
        -33.06914, -33.12204, -33.17347, -33.22525, -33.27632, -33.32646, 
        -33.37556, -33.42354, -33.47053, -33.51687, -33.56274, -33.60818, 
        -33.65318, -33.69773, -33.742, -33.786, -33.82956, -33.87243, 
        -33.91433, -33.9551, -33.99377, -34.03239, -34.07, -34.10652, 
        -34.14181, -34.1757, -34.2082, -34.23949, -34.26986, -34.29939, 
        -34.32798, -34.35572, -34.3825, -34.4084, -34.43336, -34.45714, 
        -34.4798, -34.50146, -34.52182, -34.54013, -34.55899, -34.57708, 
        -34.59489, -34.61272, -34.63065, -34.64863, -34.6664, -34.68378, 
        -34.70063, -34.71734, -34.73396, -34.75079, -34.76811, -34.78588, 
        -34.80409, -34.8227, -34.84172, -34.86116, -34.88081, -34.89965, 
        -34.91945, -34.93892, -34.95795, -34.97618, -34.99356, -35.01053, 
        -35.02736, -35.04443, -35.06232, -35.08112, -35.10099, -35.12188, 
        -35.1438, -35.16703, -35.19153, -35.21709, -35.24302, -35.26868, 
        -35.29358, -35.31783, -35.34107, -35.36261, -35.38473, -35.40608, 
        -35.42711, -35.44788, -35.46873, -35.48986, -35.51154, -35.53403, 
        -35.55743, -35.58135, -35.6055, -35.62947, -35.65319, -35.67622, 
        -35.69846, -35.71995, -35.74085, -35.76169, -35.78283, -35.80505, 
        -35.82791, -35.85072, -35.87331, -35.89537, -35.91602, -35.93779, 
        -35.96003, -35.98302, -36.00717, -36.03264, -36.06012, -36.0904, 
        -36.12433, -36.16258, -36.20549, -36.25301, -36.30437, -36.35865, 
        -36.41482, -36.47198, -36.52932, -36.58613, -36.64165, -36.69532, 
        -36.74675, -36.79586, -36.84293, -36.88837, -36.93288, -36.97674, 
        -37.02001, -37.06167, -37.10388, -37.14523, -37.186, -37.22616, 
        -37.26513, -37.3023, -37.33686, -37.36871, -37.39781, -37.42407, 
        -37.44761, -37.46891, -37.48818, -37.50586, -37.52273, -37.53928, 
        -37.55659, -37.57518, -37.59518, -37.61634, -37.63812, -37.65976, 
        -37.68052, -37.70008, -37.71824, -37.73499, -37.75051, -37.76493, 
        -37.77842, -37.79111, -37.80208, -37.81335, -37.82376, -37.83307, 
        -37.841, -37.8473, -37.85182, -37.85484, -37.85633, -37.85669, 
        -37.85682, -37.8569, -37.85766, -37.85916, -37.86147, -37.86458, 
        -37.8682, -37.87207, -37.87589, -37.87936, -37.88203, -37.88358, 
        -37.88387, -37.88307, -37.88159, -37.88005, -37.87885, -37.87791, 
        -37.87696, -37.87516, -37.87234, -37.86836, -37.86303, -37.85675, 
        -37.84934, -37.84043, -37.82998, -37.81814, -37.80489, -37.79033, 
        -37.7735, -37.75646, -37.73774, -37.71667, -37.69233, -37.66404, 
        -37.63134, -37.59381, -37.5509, -37.50208, -37.44719, -37.38658, 
        -37.32103, -37.25196, -37.1823, -37.11413, -37.04962, -36.99142, 
        -36.9419,
  -29.37125, -29.41564, -29.46073, -29.50661, -29.55321, -29.60033, 
        -29.64765, -29.69492, -29.74217, -29.7896, -29.83744, -29.88576, 
        -29.93332, -29.98221, -30.03109, -30.0796, -30.12757, -30.1749, 
        -30.22139, -30.26691, -30.31132, -30.35438, -30.39631, -30.43756, 
        -30.47857, -30.51999, -30.56197, -30.60376, -30.64779, -30.69345, 
        -30.74107, -30.7904, -30.84141, -30.89331, -30.9452, -30.99573, 
        -31.04444, -31.09073, -31.13504, -31.17811, -31.22074, -31.26365, 
        -31.30647, -31.35163, -31.3984, -31.44677, -31.49632, -31.54668, 
        -31.59705, -31.64722, -31.69637, -31.74413, -31.79037, -31.83538, 
        -31.87985, -31.9244, -31.96979, -32.01627, -32.0627, -32.11074, 
        -32.15904, -32.20717, -32.25492, -32.3023, -32.3495, -32.39688, 
        -32.44461, -32.49302, -32.54193, -32.59074, -32.63948, -32.68803, 
        -32.73667, -32.78568, -32.83559, -32.88567, -32.93777, -32.99083, 
        -33.04412, -33.09731, -33.1501, -33.20228, -33.2538, -33.30415, 
        -33.35365, -33.40211, -33.4498, -33.49683, -33.54348, -33.58976, 
        -33.63562, -33.68083, -33.72445, -33.76847, -33.81174, -33.85441, 
        -33.89618, -33.93681, -33.97635, -34.01482, -34.05222, -34.08859, 
        -34.12381, -34.15774, -34.19038, -34.22181, -34.2522, -34.28156, 
        -34.30953, -34.33644, -34.3623, -34.38636, -34.41056, -34.4339, 
        -34.45608, -34.47729, -34.49757, -34.51672, -34.53452, -34.55146, 
        -34.56818, -34.58456, -34.60106, -34.61767, -34.63432, -34.65085, 
        -34.66715, -34.68345, -34.69968, -34.71596, -34.73224, -34.7475, 
        -34.76386, -34.78048, -34.79749, -34.81516, -34.83344, -34.85227, 
        -34.87142, -34.89025, -34.90876, -34.92668, -34.94403, -34.96097, 
        -34.97786, -34.99512, -35.01286, -35.03113, -35.05032, -35.0704, 
        -35.09166, -35.11414, -35.13698, -35.16193, -35.18739, -35.21281, 
        -35.23766, -35.26195, -35.28566, -35.30869, -35.33109, -35.35286, 
        -35.3741, -35.39504, -35.41594, -35.43719, -35.45918, -35.48213, 
        -35.50607, -35.53056, -35.55538, -35.58007, -35.60433, -35.62791, 
        -35.6506, -35.67224, -35.69236, -35.71332, -35.7348, -35.75711, 
        -35.78023, -35.80363, -35.82685, -35.84974, -35.87229, -35.89501, 
        -35.91821, -35.94218, -35.96719, -35.99374, -36.02223, -36.05342, 
        -36.08828, -36.12734, -36.17107, -36.21932, -36.2713, -36.32605, 
        -36.38266, -36.44019, -36.49792, -36.55502, -36.60992, -36.66371, 
        -36.71489, -36.7634, -36.80956, -36.85412, -36.89783, -36.94101, 
        -36.98393, -37.02625, -37.06784, -37.10884, -37.14934, -37.18932, 
        -37.22807, -37.2653, -37.30017, -37.33277, -37.36264, -37.3901, 
        -37.41466, -37.43691, -37.4566, -37.4744, -37.49084, -37.50711, 
        -37.52372, -37.54132, -37.56046, -37.58086, -37.60098, -37.62204, 
        -37.64225, -37.66112, -37.67844, -37.69419, -37.70856, -37.72178, 
        -37.73402, -37.74555, -37.75655, -37.76715, -37.77724, -37.7864, 
        -37.7943, -37.80061, -37.80508, -37.80787, -37.80918, -37.80952, 
        -37.80944, -37.80981, -37.81073, -37.81259, -37.81528, -37.81861, 
        -37.82249, -37.82669, -37.83058, -37.83411, -37.83642, -37.83742, 
        -37.83703, -37.83562, -37.83374, -37.83207, -37.83, -37.8296, 
        -37.82926, -37.8287, -37.82707, -37.82414, -37.81975, -37.81424, 
        -37.80732, -37.79874, -37.78837, -37.77631, -37.76292, -37.74831, 
        -37.73266, -37.71608, -37.69807, -37.67794, -37.65485, -37.62806, 
        -37.59731, -37.56226, -37.52246, -37.47745, -37.42686, -37.37086, 
        -37.31028, -37.24646, -37.18156, -37.11781, -37.0574, -37.00212, 
        -36.95412,
  -29.36304, -29.40717, -29.45216, -29.49814, -29.54494, -29.59212, 
        -29.63922, -29.68576, -29.73075, -29.77651, -29.82249, -29.86912, 
        -29.91633, -29.96425, -30.01243, -30.06053, -30.10819, -30.15508, 
        -30.20112, -30.24589, -30.28973, -30.33238, -30.3734, -30.41495, 
        -30.45663, -30.49897, -30.54208, -30.58632, -30.63184, -30.67858, 
        -30.72673, -30.77625, -30.82674, -30.87794, -30.92893, -30.97878, 
        -31.02678, -31.07167, -31.11586, -31.15892, -31.20177, -31.24502, 
        -31.28924, -31.33471, -31.38172, -31.43023, -31.47999, -31.53053, 
        -31.58124, -31.63134, -31.68031, -31.72757, -31.77311, -31.81618, 
        -31.85942, -31.90273, -31.94687, -31.9924, -32.03934, -32.08731, 
        -32.13583, -32.18432, -32.23244, -32.27997, -32.32711, -32.37416, 
        -32.42158, -32.46975, -32.51834, -32.56644, -32.61536, -32.66429, 
        -32.71325, -32.76243, -32.81235, -32.86325, -32.91516, -32.96793, 
        -33.02116, -33.07456, -33.12775, -33.18037, -33.23226, -33.28323, 
        -33.33327, -33.38247, -33.43075, -33.47753, -33.5248, -33.57172, 
        -33.61818, -33.66386, -33.70873, -33.75269, -33.79597, -33.83851, 
        -33.8803, -33.92107, -33.96077, -33.99926, -34.03658, -34.07293, 
        -34.10816, -34.14224, -34.17509, -34.20575, -34.23614, -34.26492, 
        -34.29214, -34.31799, -34.34263, -34.36656, -34.39, -34.41261, 
        -34.43448, -34.45515, -34.47502, -34.49367, -34.51075, -34.52681, 
        -34.54216, -34.55715, -34.57197, -34.58692, -34.60112, -34.61661, 
        -34.63241, -34.64847, -34.66441, -34.68005, -34.69528, -34.71011, 
        -34.72461, -34.73915, -34.75411, -34.76982, -34.78651, -34.80405, 
        -34.82227, -34.84063, -34.85881, -34.87642, -34.8936, -34.91055, 
        -34.92751, -34.94371, -34.96123, -34.97905, -34.99741, -35.01683, 
        -35.03751, -35.05947, -35.08279, -35.10734, -35.13239, -35.15746, 
        -35.18228, -35.20673, -35.23073, -35.25411, -35.27681, -35.29876, 
        -35.32006, -35.3411, -35.36209, -35.38353, -35.40596, -35.42944, 
        -35.4529, -35.47807, -35.50358, -35.52885, -35.5536, -35.57753, 
        -35.60037, -35.62228, -35.64357, -35.66485, -35.68671, -35.70951, 
        -35.73313, -35.75723, -35.78138, -35.80534, -35.82909, -35.85294, 
        -35.87703, -35.90193, -35.92798, -35.95548, -35.98515, -36.01745, 
        -36.05329, -36.09232, -36.13697, -36.18583, -36.23835, -36.29339, 
        -36.35018, -36.40782, -36.46584, -36.52331, -36.57907, -36.63277, 
        -36.6837, -36.73145, -36.77666, -36.82023, -36.86295, -36.90545, 
        -36.94778, -36.98977, -37.03117, -37.07203, -37.11219, -37.15192, 
        -37.19065, -37.22754, -37.26287, -37.29589, -37.3269, -37.35544, 
        -37.38011, -37.40311, -37.42343, -37.44146, -37.45786, -37.47374, 
        -37.48967, -37.50642, -37.52459, -37.54409, -37.56441, -37.58476, 
        -37.60431, -37.6225, -37.639, -37.65379, -37.66709, -37.67917, 
        -37.69032, -37.70077, -37.71089, -37.72084, -37.73054, -37.73949, 
        -37.74732, -37.75352, -37.75792, -37.76051, -37.76166, -37.76209, 
        -37.76229, -37.76295, -37.76459, -37.76708, -37.76942, -37.7732, 
        -37.77738, -37.78167, -37.78522, -37.78836, -37.79007, -37.79015, 
        -37.78875, -37.78655, -37.78428, -37.78251, -37.78141, -37.78127, 
        -37.7814, -37.78157, -37.7809, -37.77918, -37.77589, -37.77138, 
        -37.76523, -37.75727, -37.74739, -37.73564, -37.7223, -37.70787, 
        -37.69254, -37.67628, -37.6587, -37.63913, -37.61694, -37.59159, 
        -37.56264, -37.53005, -37.49334, -37.45184, -37.40514, -37.35331, 
        -37.29703, -37.23769, -37.17702, -37.11718, -37.05989, -37.00704, 
        -36.95908,
  -29.35515, -29.39915, -29.44414, -29.48906, -29.53594, -29.58314, 
        -29.62997, -29.67575, -29.72067, -29.76505, -29.80934, -29.85428, 
        -29.90009, -29.94673, -29.99394, -30.04145, -30.08865, -30.13423, 
        -30.17976, -30.22407, -30.26753, -30.31029, -30.35247, -30.39455, 
        -30.43703, -30.4803, -30.52477, -30.57051, -30.6174, -30.66537, 
        -30.71415, -30.7638, -30.81297, -30.8635, -30.91363, -30.96255, 
        -31.00978, -31.05521, -31.09913, -31.14226, -31.18526, -31.22875, 
        -31.27321, -31.31899, -31.36622, -31.41481, -31.46469, -31.51533, 
        -31.56501, -31.61493, -31.66367, -31.7106, -31.75559, -31.79885, 
        -31.84107, -31.88334, -31.92639, -31.97093, -32.01723, -32.06494, 
        -32.11346, -32.16221, -32.21062, -32.25841, -32.30469, -32.35174, 
        -32.39884, -32.44651, -32.49499, -32.54436, -32.59346, -32.64262, 
        -32.69181, -32.74141, -32.79155, -32.84234, -32.89402, -32.94635, 
        -32.99924, -33.05257, -33.10592, -33.15801, -33.21052, -33.26223, 
        -33.31314, -33.36309, -33.4122, -33.46055, -33.50838, -33.55577, 
        -33.60254, -33.64859, -33.69362, -33.73777, -33.7809, -33.82351, 
        -33.86545, -33.90649, -33.94643, -33.9841, -34.02168, -34.05815, 
        -34.09362, -34.12804, -34.16127, -34.19308, -34.22325, -34.2515, 
        -34.27771, -34.30226, -34.32556, -34.34816, -34.37037, -34.39222, 
        -34.41335, -34.43366, -34.45286, -34.47083, -34.48625, -34.50138, 
        -34.51558, -34.52914, -34.54234, -34.55575, -34.56956, -34.58388, 
        -34.59886, -34.61426, -34.62962, -34.6445, -34.65866, -34.67197, 
        -34.68473, -34.69733, -34.71024, -34.72394, -34.73895, -34.7549, 
        -34.77225, -34.789, -34.80689, -34.8244, -34.84151, -34.85839, 
        -34.87532, -34.89228, -34.90944, -34.92672, -34.94448, -34.96326, 
        -34.98304, -35.00473, -35.028, -35.05226, -35.07692, -35.1018, 
        -35.12661, -35.15112, -35.17532, -35.19894, -35.22182, -35.24295, 
        -35.26423, -35.28524, -35.30624, -35.32794, -35.35073, -35.37467, 
        -35.39972, -35.42554, -35.45158, -35.47742, -35.5026, -35.52677, 
        -35.54985, -35.57206, -35.59359, -35.61541, -35.63799, -35.66146, 
        -35.68585, -35.71082, -35.73603, -35.76114, -35.78619, -35.81003, 
        -35.8352, -35.86107, -35.88818, -35.91688, -35.94761, -35.98111, 
        -36.01806, -36.0591, -36.10456, -36.15416, -36.20715, -36.26258, 
        -36.31966, -36.37756, -36.43539, -36.4928, -36.54839, -36.60169, 
        -36.65205, -36.69921, -36.74339, -36.78596, -36.82776, -36.8693, 
        -36.91092, -36.95249, -36.99273, -37.03347, -37.07363, -37.11297, 
        -37.15138, -37.1882, -37.22344, -37.25706, -37.28877, -37.31823, 
        -37.34506, -37.36888, -37.38995, -37.40845, -37.42498, -37.44062, 
        -37.45602, -37.4721, -37.48928, -37.50777, -37.52709, -37.54658, 
        -37.56537, -37.58282, -37.59855, -37.61255, -37.6249, -37.63609, 
        -37.64633, -37.65586, -37.66511, -37.67436, -37.68254, -37.69107, 
        -37.6986, -37.70469, -37.70889, -37.71144, -37.7127, -37.71333, 
        -37.71401, -37.71543, -37.71783, -37.7212, -37.72514, -37.72961, 
        -37.73393, -37.73787, -37.74112, -37.74332, -37.74379, -37.74271, 
        -37.74031, -37.73738, -37.73462, -37.73268, -37.73161, -37.73135, 
        -37.73173, -37.73212, -37.73221, -37.73141, -37.72949, -37.7263, 
        -37.7214, -37.71457, -37.70567, -37.6947, -37.68199, -37.66795, 
        -37.65284, -37.6366, -37.61808, -37.59878, -37.57727, -37.55312, 
        -37.52602, -37.49576, -37.4618, -37.42356, -37.38054, -37.33248, 
        -37.28022, -37.22488, -37.16806, -37.11149, -37.05689, -37.00582, 
        -36.95945,
  -29.34666, -29.39031, -29.43505, -29.48086, -29.52757, -29.57461, 
        -29.62113, -29.66654, -29.71068, -29.754, -29.79691, -29.8404, 
        -29.88493, -29.92932, -29.97559, -30.02229, -30.06893, -30.11501, 
        -30.1602, -30.20438, -30.24778, -30.29058, -30.33316, -30.37595, 
        -30.41929, -30.46361, -30.5093, -30.55624, -30.60344, -30.65235, 
        -30.70175, -30.75141, -30.80129, -30.85096, -30.90026, -30.94831, 
        -30.99494, -31.03989, -31.08376, -31.12686, -31.17002, -31.21374, 
        -31.25836, -31.30333, -31.35065, -31.39925, -31.44898, -31.49939, 
        -31.54989, -31.59971, -31.64835, -31.69504, -31.73962, -31.78237, 
        -31.82397, -31.86542, -31.90753, -31.95119, -31.99671, -32.04293, 
        -32.09118, -32.13988, -32.18843, -32.23647, -32.28392, -32.33111, 
        -32.37824, -32.42599, -32.47435, -32.52322, -32.5726, -32.62198, 
        -32.6715, -32.72137, -32.77149, -32.8222, -32.87251, -32.92446, 
        -32.9771, -33.03015, -33.08368, -33.13728, -33.19053, -33.24315, 
        -33.29495, -33.34579, -33.39564, -33.44463, -33.49293, -33.54068, 
        -33.58777, -33.63403, -33.67918, -33.72239, -33.76571, -33.8084, 
        -33.85049, -33.8918, -33.932, -33.97103, -34.00893, -34.0458, 
        -34.08172, -34.11663, -34.15027, -34.18229, -34.21225, -34.23981, 
        -34.26496, -34.28817, -34.31005, -34.33126, -34.35118, -34.37189, 
        -34.39219, -34.41175, -34.4303, -34.44748, -34.46315, -34.47741, 
        -34.49044, -34.50265, -34.51447, -34.52637, -34.5387, -34.55176, 
        -34.56563, -34.57998, -34.59427, -34.60806, -34.62092, -34.63283, 
        -34.64301, -34.65389, -34.66497, -34.67691, -34.69011, -34.70473, 
        -34.72121, -34.73844, -34.75581, -34.77318, -34.79011, -34.80674, 
        -34.82332, -34.83995, -34.85654, -34.87327, -34.8904, -34.90874, 
        -34.9285, -34.95003, -34.97308, -34.9971, -35.02056, -35.04515, 
        -35.06982, -35.09444, -35.11872, -35.14254, -35.1656, -35.18763, 
        -35.20897, -35.23, -35.25108, -35.27288, -35.29585, -35.32013, 
        -35.34562, -35.37192, -35.3985, -35.42482, -35.45037, -35.47483, 
        -35.49822, -35.52081, -35.54308, -35.5647, -35.58812, -35.61251, 
        -35.63779, -35.66369, -35.68988, -35.71608, -35.74215, -35.76819, 
        -35.79433, -35.82129, -35.84948, -35.87942, -35.91152, -35.94638, 
        -35.98458, -36.02674, -36.07305, -36.12344, -36.17695, -36.23273, 
        -36.28994, -36.34779, -36.40562, -36.4626, -36.51787, -36.56956, 
        -36.61911, -36.66548, -36.70906, -36.75072, -36.79148, -36.83207, 
        -36.87301, -36.91399, -36.95482, -36.99533, -37.03526, -37.07441, 
        -37.11242, -37.14907, -37.1843, -37.21807, -37.25031, -37.28063, 
        -37.30833, -37.33304, -37.35471, -37.37366, -37.39059, -37.40634, 
        -37.42159, -37.43707, -37.45338, -37.47075, -37.48902, -37.50751, 
        -37.52444, -37.5411, -37.55606, -37.56934, -37.58105, -37.59153, 
        -37.60093, -37.60967, -37.61813, -37.62659, -37.63501, -37.64309, 
        -37.65007, -37.6557, -37.65983, -37.66246, -37.66398, -37.6651, 
        -37.6664, -37.66859, -37.67191, -37.67619, -37.68103, -37.686, 
        -37.69035, -37.69362, -37.69598, -37.6968, -37.69605, -37.69371, 
        -37.69036, -37.68669, -37.68345, -37.68106, -37.67968, -37.67931, 
        -37.67953, -37.67916, -37.67975, -37.67986, -37.67924, -37.6775, 
        -37.67428, -37.66906, -37.66166, -37.65194, -37.64021, -37.62671, 
        -37.61181, -37.59553, -37.57784, -37.55862, -37.53762, -37.51454, 
        -37.48913, -37.46105, -37.4298, -37.3945, -37.35476, -37.31026, 
        -37.26173, -37.21006, -37.15679, -37.10316, -37.0507, -37.0008, 
        -36.95445,
  -29.33933, -29.38264, -29.42683, -29.47219, -29.51845, -29.56502, 
        -29.61127, -29.65632, -29.69903, -29.74169, -29.78403, -29.82665, 
        -29.87002, -29.91448, -29.95983, -30.00574, -30.05173, -30.09739, 
        -30.14238, -30.18654, -30.23006, -30.27309, -30.31614, -30.35855, 
        -30.40264, -30.44792, -30.49465, -30.54267, -30.59156, -30.64105, 
        -30.69079, -30.74037, -30.78976, -30.83881, -30.88744, -30.9349, 
        -30.98082, -31.02561, -31.06841, -31.11171, -31.15506, -31.19901, 
        -31.24391, -31.28996, -31.33723, -31.38563, -31.435, -31.48492, 
        -31.53495, -31.58454, -31.63291, -31.6795, -31.72405, -31.7667, 
        -31.80708, -31.84803, -31.88952, -31.9324, -31.97706, -32.02348, 
        -32.07116, -32.11948, -32.16787, -32.21595, -32.2635, -32.3109, 
        -32.35838, -32.40613, -32.45449, -32.50341, -32.55167, -32.60116, 
        -32.65095, -32.70106, -32.75126, -32.8019, -32.85291, -32.90459, 
        -32.95676, -33.00942, -33.06309, -33.11723, -33.17134, -33.22493, 
        -33.27765, -33.32922, -33.37966, -33.42921, -33.47709, -33.52523, 
        -33.57259, -33.61906, -33.66446, -33.70888, -33.75243, -33.79531, 
        -33.83757, -33.87912, -33.91957, -33.95891, -33.9972, -34.0345, 
        -34.07101, -34.10649, -34.14061, -34.17281, -34.20157, -34.22846, 
        -34.25266, -34.27467, -34.29524, -34.31516, -34.33475, -34.35422, 
        -34.37342, -34.39204, -34.4097, -34.42598, -34.44067, -34.45406, 
        -34.46602, -34.47701, -34.48748, -34.49791, -34.50884, -34.52041, 
        -34.53185, -34.54485, -34.55774, -34.57004, -34.58139, -34.59187, 
        -34.60163, -34.61103, -34.62057, -34.63089, -34.64253, -34.6561, 
        -34.67168, -34.68834, -34.70537, -34.72229, -34.73882, -34.75505, 
        -34.77098, -34.78693, -34.80286, -34.81805, -34.83493, -34.85306, 
        -34.87284, -34.89444, -34.91743, -34.94125, -34.96544, -34.98968, 
        -35.01427, -35.03889, -35.06335, -35.08728, -35.11029, -35.13241, 
        -35.15366, -35.17451, -35.19557, -35.21745, -35.2406, -35.2652, 
        -35.29105, -35.31776, -35.34377, -35.37049, -35.39634, -35.42105, 
        -35.44475, -35.46786, -35.49093, -35.51471, -35.5393, -35.56483, 
        -35.5911, -35.6179, -35.64495, -35.67207, -35.69904, -35.72598, 
        -35.75328, -35.78126, -35.81068, -35.84185, -35.87534, -35.91155, 
        -35.9511, -35.99442, -36.04179, -36.09188, -36.14596, -36.20215, 
        -36.25955, -36.31741, -36.375, -36.43158, -36.48619, -36.53814, 
        -36.58703, -36.63276, -36.67571, -36.71675, -36.75653, -36.79613, 
        -36.83606, -36.87628, -36.91655, -36.95691, -36.99667, -37.03552, 
        -37.07313, -37.10951, -37.14465, -37.17852, -37.21099, -37.2417, 
        -37.26996, -37.29523, -37.31656, -37.33619, -37.35373, -37.37002, 
        -37.3854, -37.40056, -37.41606, -37.4323, -37.44926, -37.4666, 
        -37.48353, -37.49938, -37.51369, -37.52634, -37.53745, -37.54723, 
        -37.55601, -37.56408, -37.57182, -37.57955, -37.58714, -37.59447, 
        -37.6008, -37.60617, -37.61016, -37.61289, -37.61473, -37.61628, 
        -37.61826, -37.62128, -37.62552, -37.63069, -37.63628, -37.64149, 
        -37.64459, -37.64725, -37.64837, -37.6477, -37.64546, -37.64187, 
        -37.63755, -37.63323, -37.62945, -37.62661, -37.62477, -37.62392, 
        -37.62392, -37.62455, -37.62553, -37.62654, -37.6272, -37.62711, 
        -37.62574, -37.62248, -37.61689, -37.60881, -37.5983, -37.58557, 
        -37.57093, -37.55459, -37.5367, -37.51746, -37.49693, -37.47496, 
        -37.45125, -37.42533, -37.39653, -37.36409, -37.32733, -37.28608, 
        -37.2409, -37.19273, -37.14249, -37.0915, -37.04099, -36.99179, 
        -36.94508,
  -29.33234, -29.37487, -29.41834, -29.46295, -29.50743, -29.55336, 
        -29.5991, -29.64388, -29.68749, -29.73013, -29.77225, -29.81455, 
        -29.85765, -29.90132, -29.94587, -29.99112, -30.03658, -30.08184, 
        -30.12566, -30.16984, -30.21357, -30.25697, -30.30052, -30.34461, 
        -30.38942, -30.43542, -30.48286, -30.53145, -30.58089, -30.63058, 
        -30.68006, -30.7295, -30.77834, -30.82576, -30.87361, -30.92052, 
        -30.9664, -31.01136, -31.0553, -31.09907, -31.14276, -31.18701, 
        -31.23217, -31.27831, -31.32541, -31.37336, -31.422, -31.4711, 
        -31.52039, -31.56845, -31.61654, -31.66316, -31.70802, -31.75093, 
        -31.79251, -31.83334, -31.87438, -31.91648, -31.96021, -32.00563, 
        -32.05245, -32.10006, -32.14803, -32.19605, -32.2436, -32.29028, 
        -32.33796, -32.38584, -32.43451, -32.48349, -32.53275, -32.5823, 
        -32.63221, -32.68236, -32.73259, -32.78342, -32.83406, -32.88529, 
        -32.93704, -32.98986, -33.04358, -33.09819, -33.15205, -33.20643, 
        -33.2599, -33.31218, -33.363, -33.41302, -33.46229, -33.51102, 
        -33.55898, -33.60583, -33.65166, -33.69654, -33.74053, -33.78352, 
        -33.82591, -33.86749, -33.90815, -33.94767, -33.98524, -34.02305, 
        -34.06, -34.09599, -34.13057, -34.16297, -34.19243, -34.21873, 
        -34.24228, -34.26353, -34.28323, -34.30205, -34.32039, -34.33863, 
        -34.35661, -34.37406, -34.39061, -34.40571, -34.41953, -34.43067, 
        -34.44156, -34.45126, -34.46048, -34.46953, -34.47896, -34.48919, 
        -34.49994, -34.51115, -34.52232, -34.53284, -34.54263, -34.55174, 
        -34.56015, -34.56821, -34.57647, -34.58549, -34.59614, -34.60889, 
        -34.62353, -34.63955, -34.65501, -34.67131, -34.68708, -34.7024, 
        -34.71745, -34.73257, -34.74786, -34.76373, -34.7806, -34.799, 
        -34.81902, -34.84083, -34.86372, -34.88725, -34.91114, -34.93515, 
        -34.95931, -34.9838, -35.00825, -35.0322, -35.05522, -35.07715, 
        -35.09719, -35.1179, -35.13889, -35.16095, -35.18443, -35.20941, 
        -35.23561, -35.26266, -35.28993, -35.31699, -35.34301, -35.36781, 
        -35.39174, -35.4154, -35.43959, -35.46462, -35.49059, -35.51741, 
        -35.54473, -35.57236, -35.60012, -35.62785, -35.65554, -35.68336, 
        -35.71164, -35.73987, -35.77044, -35.80296, -35.83786, -35.87552, 
        -35.91653, -35.9612, -36.00956, -36.06145, -36.11609, -36.17267, 
        -36.23022, -36.28797, -36.34533, -36.40123, -36.45518, -36.5066, 
        -36.55489, -36.60013, -36.64268, -36.68318, -36.72219, -36.76077, 
        -36.79955, -36.83897, -36.87883, -36.91843, -36.95693, -36.99544, 
        -37.03273, -37.06871, -37.10361, -37.13739, -37.16982, -37.20047, 
        -37.2289, -37.25458, -37.27749, -37.29801, -37.31655, -37.3337, 
        -37.34951, -37.3646, -37.37949, -37.39465, -37.41028, -37.42619, 
        -37.44199, -37.45686, -37.47044, -37.4825, -37.49302, -37.5023, 
        -37.51052, -37.51803, -37.52515, -37.53216, -37.53897, -37.54545, 
        -37.5503, -37.55513, -37.55904, -37.56171, -37.56401, -37.56624, 
        -37.56886, -37.57264, -37.57757, -37.58341, -37.58936, -37.59453, 
        -37.59822, -37.59995, -37.59961, -37.59742, -37.59381, -37.58904, 
        -37.58391, -37.57898, -37.57466, -37.57122, -37.5689, -37.56752, 
        -37.56721, -37.56771, -37.56903, -37.5709, -37.57278, -37.57437, 
        -37.57499, -37.5738, -37.57024, -37.56396, -37.55479, -37.543, 
        -37.52876, -37.51251, -37.49466, -37.47554, -37.45555, -37.43383, 
        -37.41188, -37.38823, -37.36181, -37.33195, -37.29787, -37.25954, 
        -37.21743, -37.17225, -37.12503, -37.07632, -37.0272, -36.97863, 
        -36.93149,
  -29.32437, -29.36605, -29.40868, -29.4523, -29.49694, -29.54217, 
        -29.58737, -29.63186, -29.67548, -29.71819, -29.76051, -29.80281, 
        -29.84563, -29.88918, -29.93224, -29.97703, -30.02225, -30.0674, 
        -30.11222, -30.1566, -30.20046, -30.24408, -30.28805, -30.33264, 
        -30.37818, -30.42492, -30.47297, -30.52206, -30.57158, -30.62035, 
        -30.66964, -30.7184, -30.76658, -30.8142, -30.86129, -30.90764, 
        -30.95342, -30.99867, -31.04346, -31.08797, -31.13251, -31.17736, 
        -31.22276, -31.26879, -31.31434, -31.36143, -31.4091, -31.45711, 
        -31.50556, -31.55412, -31.60214, -31.649, -31.69412, -31.73759, 
        -31.77948, -31.82043, -31.86124, -31.90271, -31.94546, -31.98975, 
        -32.03448, -32.08125, -32.12864, -32.17634, -32.22412, -32.27192, 
        -32.31988, -32.36803, -32.41661, -32.46555, -32.51471, -32.56404, 
        -32.61357, -32.66352, -32.71372, -32.76448, -32.8153, -32.86596, 
        -32.91755, -32.97046, -33.02458, -33.07955, -33.1349, -33.1899, 
        -33.24387, -33.29649, -33.34772, -33.39832, -33.44809, -33.49747, 
        -33.54601, -33.5935, -33.6399, -33.68534, -33.72869, -33.77212, 
        -33.8146, -33.85612, -33.89669, -33.93633, -33.97511, -34.01317, 
        -34.05064, -34.08702, -34.12189, -34.1542, -34.18352, -34.20967, 
        -34.23273, -34.25344, -34.2726, -34.29064, -34.30809, -34.32421, 
        -34.34101, -34.35721, -34.37241, -34.38633, -34.39871, -34.40969, 
        -34.4192, -34.42755, -34.43548, -34.44321, -34.45126, -34.45978, 
        -34.46885, -34.47808, -34.48724, -34.49596, -34.5041, -34.51168, 
        -34.51883, -34.52478, -34.5321, -34.54038, -34.55044, -34.56247, 
        -34.57635, -34.59143, -34.60698, -34.62222, -34.63691, -34.65112, 
        -34.66515, -34.67936, -34.69413, -34.70988, -34.72701, -34.74594, 
        -34.76634, -34.78827, -34.8111, -34.83437, -34.85786, -34.88055, 
        -34.90453, -34.92875, -34.953, -34.97672, -34.99948, -35.02106, 
        -35.04182, -35.06237, -35.08348, -35.10568, -35.12943, -35.15474, 
        -35.18131, -35.20866, -35.23623, -35.26339, -35.28959, -35.31452, 
        -35.33875, -35.36295, -35.38808, -35.41432, -35.44165, -35.46883, 
        -35.49733, -35.5258, -35.55418, -35.58245, -35.61072, -35.63926, 
        -35.66847, -35.69879, -35.73068, -35.76466, -35.80101, -35.84031, 
        -35.88292, -35.92889, -35.97834, -36.03094, -36.08595, -36.14267, 
        -36.20024, -36.25783, -36.31469, -36.37016, -36.42354, -36.47435, 
        -36.52227, -36.5663, -36.6087, -36.64868, -36.68723, -36.72509, 
        -36.76315, -36.8018, -36.84087, -36.88017, -36.91886, -36.95692, 
        -36.99371, -37.02926, -37.06361, -37.09701, -37.12905, -37.15946, 
        -37.18779, -37.21375, -37.23735, -37.25879, -37.27861, -37.29662, 
        -37.3131, -37.32826, -37.34268, -37.3569, -37.37116, -37.38557, 
        -37.39992, -37.41363, -37.4253, -37.4367, -37.44672, -37.45556, 
        -37.46339, -37.47046, -37.47706, -37.48344, -37.48957, -37.49533, 
        -37.5005, -37.50503, -37.5086, -37.51165, -37.51417, -37.51705, 
        -37.52038, -37.52483, -37.53028, -37.53627, -37.54216, -37.54694, 
        -37.54984, -37.55046, -37.54881, -37.54509, -37.54033, -37.53474, 
        -37.52886, -37.52327, -37.51843, -37.51451, -37.51167, -37.5099, 
        -37.50941, -37.51014, -37.5118, -37.5133, -37.51631, -37.51931, 
        -37.52155, -37.52225, -37.52053, -37.51588, -37.50809, -37.49737, 
        -37.48395, -37.46825, -37.45093, -37.43248, -37.41342, -37.39407, 
        -37.37395, -37.35233, -37.32816, -37.30063, -37.26899, -37.23322, 
        -37.19383, -37.15137, -37.10649, -37.05986, -37.01194, -36.96393, 
        -36.91649,
  -29.31758, -29.35833, -29.39996, -29.4426, -29.48631, -29.53074, 
        -29.57543, -29.61976, -29.66343, -29.70548, -29.74811, -29.79067, 
        -29.83351, -29.87679, -29.92074, -29.9654, -30.01054, -30.05574, 
        -30.10066, -30.14507, -30.18932, -30.23343, -30.27785, -30.32291, 
        -30.36811, -30.41541, -30.46382, -30.51319, -30.5627, -30.6122, 
        -30.66121, -30.70941, -30.75692, -30.80377, -30.84996, -30.89592, 
        -30.94161, -30.98737, -31.03316, -31.07787, -31.12353, -31.16916, 
        -31.21484, -31.26053, -31.30628, -31.35223, -31.3985, -31.4453, 
        -31.49278, -31.54076, -31.58868, -31.63588, -31.68167, -31.72568, 
        -31.76807, -31.80834, -31.84908, -31.89011, -31.93198, -31.97511, 
        -32.01961, -32.06539, -32.11204, -32.15947, -32.20721, -32.2552, 
        -32.30335, -32.35161, -32.40014, -32.44883, -32.49762, -32.54553, 
        -32.5947, -32.64434, -32.69447, -32.74535, -32.79671, -32.84846, 
        -32.90121, -32.95448, -33.00863, -33.06372, -33.11923, -33.17456, 
        -33.22869, -33.28154, -33.33317, -33.38403, -33.43457, -33.48363, 
        -33.53289, -33.58116, -33.6283, -33.67442, -33.7193, -33.76292, 
        -33.80541, -33.84676, -33.88718, -33.92673, -33.96559, -34.00384, 
        -34.04151, -34.07817, -34.11304, -34.14542, -34.17469, -34.19957, 
        -34.22245, -34.24305, -34.26194, -34.27959, -34.29634, -34.31252, 
        -34.32822, -34.34319, -34.35708, -34.36958, -34.38057, -34.38993, 
        -34.39796, -34.40488, -34.41142, -34.41792, -34.42462, -34.43163, 
        -34.43885, -34.44513, -34.45223, -34.45901, -34.46538, -34.47146, 
        -34.47725, -34.48315, -34.48965, -34.49742, -34.50705, -34.51855, 
        -34.53166, -34.54568, -34.55993, -34.57381, -34.58729, -34.60032, 
        -34.61332, -34.62674, -34.64114, -34.65701, -34.67356, -34.69294, 
        -34.71401, -34.73592, -34.75851, -34.7814, -34.80453, -34.82788, 
        -34.85167, -34.87573, -34.89965, -34.92296, -34.94522, -34.96629, 
        -34.9867, -35.00707, -35.02819, -35.05059, -35.07463, -35.10025, 
        -35.12714, -35.15479, -35.18266, -35.20904, -35.23529, -35.26031, 
        -35.28471, -35.30947, -35.33535, -35.36271, -35.39151, -35.42094, 
        -35.45061, -35.48003, -35.50906, -35.53788, -35.56678, -35.59608, 
        -35.62627, -35.65777, -35.69099, -35.72642, -35.76435, -35.8053, 
        -35.84947, -35.89676, -35.94725, -36.00035, -36.0545, -36.11101, 
        -36.16826, -36.22545, -36.28196, -36.33696, -36.38995, -36.44047, 
        -36.48829, -36.53326, -36.57555, -36.6154, -36.65357, -36.69095, 
        -36.72849, -36.76663, -36.80525, -36.84379, -36.88181, -36.91882, 
        -36.95495, -36.98984, -37.02357, -37.05642, -37.08791, -37.11783, 
        -37.14583, -37.17192, -37.19621, -37.21771, -37.23858, -37.2577, 
        -37.27483, -37.29028, -37.30441, -37.31779, -37.33075, -37.34362, 
        -37.35632, -37.36862, -37.3802, -37.39088, -37.40049, -37.40906, 
        -37.41667, -37.42346, -37.42973, -37.43562, -37.44121, -37.4464, 
        -37.45117, -37.4552, -37.45872, -37.46179, -37.46469, -37.46823, 
        -37.4724, -37.47745, -37.48294, -37.48869, -37.4938, -37.49775, 
        -37.49947, -37.49894, -37.49519, -37.49041, -37.48469, -37.47832, 
        -37.47187, -37.46576, -37.46028, -37.4558, -37.45266, -37.45084, 
        -37.45046, -37.45118, -37.45318, -37.45625, -37.46012, -37.46418, 
        -37.46774, -37.46988, -37.46969, -37.46651, -37.46007, -37.45049, 
        -37.43835, -37.4239, -37.40775, -37.39056, -37.37284, -37.35491, 
        -37.33648, -37.31679, -37.2947, -37.2692, -37.23978, -37.20642, 
        -37.16951, -37.12951, -37.08672, -37.04162, -36.99494, -36.94736, 
        -36.8998,
  -29.31086, -29.35059, -29.39131, -29.43314, -29.47608, -29.51883, 
        -29.56301, -29.60711, -29.65076, -29.69399, -29.73689, -29.7797, 
        -29.82269, -29.86606, -29.91009, -29.95482, -30.00004, -30.04531, 
        -30.09032, -30.13399, -30.17843, -30.22301, -30.26804, -30.3139, 
        -30.36079, -30.40876, -30.45766, -30.50711, -30.55683, -30.60604, 
        -30.6544, -30.70192, -30.74854, -30.79454, -30.83904, -30.88457, 
        -30.93047, -30.97688, -31.02381, -31.07092, -31.11781, -31.16424, 
        -31.21009, -31.25533, -31.30006, -31.34464, -31.38942, -31.43492, 
        -31.48145, -31.52896, -31.5759, -31.62349, -31.66991, -31.71459, 
        -31.75761, -31.79922, -31.83999, -31.88066, -31.92174, -31.9638, 
        -32.00719, -32.05195, -32.09796, -32.14496, -32.19262, -32.24049, 
        -32.28784, -32.33599, -32.38425, -32.43243, -32.48064, -32.52899, 
        -32.57769, -32.627, -32.67723, -32.72838, -32.78036, -32.83303, 
        -32.88646, -32.94045, -32.99507, -33.05032, -33.10602, -33.16045, 
        -33.21484, -33.26787, -33.31972, -33.37075, -33.42147, -33.47192, 
        -33.52188, -33.57091, -33.6187, -33.66525, -33.71045, -33.75422, 
        -33.79662, -33.83781, -33.87806, -33.91756, -33.95642, -33.99374, 
        -34.03157, -34.06834, -34.10324, -34.13573, -34.16479, -34.19064, 
        -34.21341, -34.23405, -34.2527, -34.27001, -34.28628, -34.30171, 
        -34.31642, -34.3303, -34.34304, -34.35418, -34.36367, -34.37152, 
        -34.37802, -34.3825, -34.38762, -34.39275, -34.39812, -34.40361, 
        -34.40916, -34.41455, -34.41971, -34.42459, -34.4291, -34.43344, 
        -34.43779, -34.44255, -34.4482, -34.45544, -34.46462, -34.47557, 
        -34.48789, -34.50084, -34.51369, -34.52519, -34.53733, -34.54927, 
        -34.56137, -34.57417, -34.58831, -34.60427, -34.62219, -34.64198, 
        -34.66326, -34.6852, -34.70758, -34.73011, -34.75293, -34.77612, 
        -34.79972, -34.82353, -34.8471, -34.86988, -34.89154, -34.91216, 
        -34.93223, -34.95148, -34.97255, -34.99503, -35.0192, -35.045, 
        -35.07211, -35.09998, -35.12814, -35.15578, -35.18223, -35.20748, 
        -35.23213, -35.25721, -35.28371, -35.31197, -35.34175, -35.37235, 
        -35.40318, -35.43362, -35.46354, -35.49322, -35.52294, -35.55314, 
        -35.58445, -35.6172, -35.65083, -35.68774, -35.72728, -35.76985, 
        -35.81541, -35.86401, -35.91527, -35.96869, -36.02375, -36.07987, 
        -36.13664, -36.19334, -36.24926, -36.30398, -36.35668, -36.40699, 
        -36.45475, -36.49976, -36.542, -36.58174, -36.61973, -36.65698, 
        -36.69437, -36.73236, -36.77062, -36.80864, -36.84585, -36.88205, 
        -36.91597, -36.94981, -36.98268, -37.01471, -37.04554, -37.07497, 
        -37.10282, -37.12907, -37.15382, -37.17715, -37.19894, -37.2188, 
        -37.23666, -37.25243, -37.26646, -37.2792, -37.29105, -37.30241, 
        -37.31346, -37.32417, -37.33444, -37.34419, -37.3532, -37.36154, 
        -37.36906, -37.37583, -37.38197, -37.38766, -37.39296, -37.39775, 
        -37.40203, -37.40568, -37.40787, -37.41099, -37.41447, -37.41858, 
        -37.42332, -37.42872, -37.43435, -37.43971, -37.44417, -37.44692, 
        -37.44762, -37.44609, -37.44208, -37.43644, -37.42975, -37.42271, 
        -37.41582, -37.40927, -37.40343, -37.39868, -37.39523, -37.39343, 
        -37.39306, -37.39402, -37.39633, -37.39976, -37.40404, -37.40866, 
        -37.41301, -37.41614, -37.41705, -37.41516, -37.41011, -37.40209, 
        -37.39153, -37.37887, -37.36464, -37.34914, -37.33309, -37.31672, 
        -37.29984, -37.28171, -37.2603, -37.23663, -37.20919, -37.17799, 
        -37.14329, -37.10534, -37.06443, -37.02084, -36.97516, -36.92816, 
        -36.88075,
  -29.30346, -29.34234, -29.38237, -29.42353, -29.46589, -29.50907, 
        -29.5527, -29.59644, -29.64, -29.68329, -29.72631, -29.76932, 
        -29.8125, -29.85612, -29.9004, -29.94441, -29.9898, -30.03519, 
        -30.08035, -30.12517, -30.17003, -30.21514, -30.26089, -30.30753, 
        -30.35517, -30.40374, -30.45306, -30.5028, -30.55238, -30.60034, 
        -30.64829, -30.69513, -30.74101, -30.78626, -30.83129, -30.87659, 
        -30.92264, -30.96971, -31.01762, -31.06604, -31.11407, -31.1612, 
        -31.20713, -31.25177, -31.29549, -31.33773, -31.38115, -31.42549, 
        -31.47116, -31.51816, -31.56617, -31.61401, -31.66095, -31.70627, 
        -31.74975, -31.79169, -31.83248, -31.87285, -31.91332, -31.95453, 
        -31.99702, -32.03991, -32.08525, -32.1317, -32.17906, -32.22677, 
        -32.27482, -32.32287, -32.37081, -32.41858, -32.46627, -32.5141, 
        -32.5624, -32.61152, -32.66179, -32.71334, -32.7661, -32.81967, 
        -32.87307, -32.9279, -32.98301, -33.03853, -33.0943, -33.14976, 
        -33.20431, -33.25739, -33.30933, -33.36046, -33.41118, -33.46186, 
        -33.51219, -33.56177, -33.61009, -33.65696, -33.70224, -33.7459, 
        -33.78708, -33.82802, -33.868, -33.9072, -33.94603, -33.98442, 
        -34.02234, -34.05921, -34.0942, -34.12654, -34.15561, -34.1813, 
        -34.20419, -34.22461, -34.24326, -34.26003, -34.27593, -34.29073, 
        -34.30364, -34.31676, -34.32845, -34.33843, -34.34658, -34.35299, 
        -34.35799, -34.36209, -34.36579, -34.36957, -34.37359, -34.37778, 
        -34.38191, -34.38572, -34.38916, -34.39224, -34.39484, -34.39732, 
        -34.39996, -34.40322, -34.40677, -34.41321, -34.42178, -34.43214, 
        -34.44361, -34.45543, -34.467, -34.47827, -34.48928, -34.50027, 
        -34.51164, -34.52399, -34.53793, -34.554, -34.57218, -34.59219, 
        -34.61344, -34.63531, -34.65733, -34.6795, -34.70198, -34.72501, 
        -34.74749, -34.77106, -34.79426, -34.81662, -34.83778, -34.85794, 
        -34.87772, -34.89775, -34.91872, -34.94117, -34.96531, -34.99114, 
        -35.01839, -35.04658, -35.07501, -35.10289, -35.12961, -35.15504, 
        -35.17993, -35.20531, -35.23218, -35.26095, -35.2914, -35.32302, 
        -35.35384, -35.38544, -35.41648, -35.44728, -35.47825, -35.50974, 
        -35.54241, -35.57663, -35.61283, -35.65132, -35.69238, -35.73637, 
        -35.7833, -35.83294, -35.88483, -35.9384, -35.99316, -36.04884, 
        -36.10489, -36.16111, -36.21667, -36.27099, -36.32343, -36.37363, 
        -36.42125, -36.46597, -36.50803, -36.5466, -36.58445, -36.6218, 
        -36.65947, -36.69749, -36.73556, -36.77308, -36.80952, -36.84461, 
        -36.87836, -36.91093, -36.94251, -36.97353, -37.00363, -37.03265, 
        -37.06044, -37.08681, -37.11184, -37.1357, -37.1581, -37.17862, 
        -37.19701, -37.21327, -37.22746, -37.23987, -37.25093, -37.26106, 
        -37.27044, -37.2795, -37.28831, -37.29691, -37.30417, -37.31223, 
        -37.31974, -37.32663, -37.33289, -37.33859, -37.34371, -37.34823, 
        -37.3521, -37.35532, -37.35822, -37.36129, -37.36508, -37.36969, 
        -37.37508, -37.38087, -37.38644, -37.39129, -37.39494, -37.39681, 
        -37.39651, -37.39376, -37.38903, -37.38256, -37.37519, -37.36763, 
        -37.36032, -37.35353, -37.34755, -37.34269, -37.33914, -37.33727, 
        -37.33704, -37.33822, -37.34066, -37.34422, -37.34851, -37.35234, 
        -37.35699, -37.3607, -37.36247, -37.3616, -37.35789, -37.35159, 
        -37.34298, -37.33258, -37.32056, -37.30738, -37.29327, -37.27838, 
        -37.26266, -37.24566, -37.22658, -37.20438, -37.17865, -37.14939, 
        -37.1167, -37.08064, -37.04144, -36.99932, -36.95483, -36.90861, 
        -36.86156,
  -29.29778, -29.33602, -29.37563, -29.4166, -29.45858, -29.50131, 
        -29.54438, -29.58759, -29.63079, -29.674, -29.71611, -29.75922, 
        -29.80248, -29.84641, -29.89107, -29.93638, -29.98201, -30.02757, 
        -30.07291, -30.11802, -30.16332, -30.20909, -30.25561, -30.30304, 
        -30.35135, -30.39945, -30.4492, -30.49914, -30.54874, -30.59745, 
        -30.6449, -30.6912, -30.73655, -30.78133, -30.82602, -30.87125, 
        -30.91758, -30.96511, -31.01379, -31.06296, -31.11083, -31.15834, 
        -31.20432, -31.2485, -31.29136, -31.33354, -31.37579, -31.41913, 
        -31.46428, -31.51085, -31.55861, -31.60669, -31.6538, -31.69951, 
        -31.74332, -31.78539, -31.82514, -31.86523, -31.90519, -31.94585, 
        -31.98765, -32.03087, -32.07547, -32.12149, -32.16838, -32.21591, 
        -32.26366, -32.31131, -32.35898, -32.4063, -32.45362, -32.50102, 
        -32.548, -32.59702, -32.64755, -32.69942, -32.75311, -32.80753, 
        -32.8629, -32.9186, -32.97423, -33.03009, -33.08586, -33.14128, 
        -33.19588, -33.2489, -33.30095, -33.35194, -33.40267, -33.45338, 
        -33.50283, -33.55262, -33.60128, -33.64824, -33.69342, -33.73664, 
        -33.77841, -33.81895, -33.85857, -33.89764, -33.93641, -33.97489, 
        -34.01285, -34.04981, -34.08476, -34.11705, -34.14602, -34.17163, 
        -34.19332, -34.21365, -34.23196, -34.24838, -34.26357, -34.27767, 
        -34.29126, -34.30362, -34.31455, -34.32368, -34.33081, -34.33613, 
        -34.33992, -34.34265, -34.34485, -34.34725, -34.34996, -34.35296, 
        -34.35587, -34.35847, -34.35955, -34.36098, -34.36176, -34.36221, 
        -34.36293, -34.36437, -34.36745, -34.37277, -34.38043, -34.39001, 
        -34.40049, -34.41123, -34.42175, -34.43195, -34.44206, -34.45232, 
        -34.46313, -34.47525, -34.48909, -34.50517, -34.52346, -34.54247, 
        -34.5635, -34.58503, -34.60666, -34.62851, -34.6508, -34.67371, 
        -34.69713, -34.72043, -34.74321, -34.76519, -34.78593, -34.80581, 
        -34.82536, -34.84517, -34.86599, -34.88826, -34.91232, -34.93812, 
        -34.96544, -34.99377, -35.02237, -35.05045, -35.07635, -35.10206, 
        -35.12724, -35.15279, -35.17987, -35.20885, -35.23965, -35.2718, 
        -35.30473, -35.3373, -35.37003, -35.40231, -35.43493, -35.46811, 
        -35.50239, -35.53826, -35.57608, -35.61615, -35.65872, -35.70401, 
        -35.7521, -35.80264, -35.85505, -35.90875, -35.96328, -36.01844, 
        -36.07304, -36.12868, -36.18389, -36.23796, -36.29018, -36.34007, 
        -36.38717, -36.43132, -36.47294, -36.51206, -36.55001, -36.5876, 
        -36.62552, -36.66365, -36.70158, -36.7386, -36.77422, -36.80816, 
        -36.84047, -36.87152, -36.90176, -36.93147, -36.96072, -36.98945, 
        -37.01715, -37.04364, -37.06895, -37.09303, -37.11559, -37.13547, 
        -37.15438, -37.17105, -37.18569, -37.19827, -37.209, -37.2182, 
        -37.22624, -37.23378, -37.24101, -37.24828, -37.25576, -37.26327, 
        -37.27087, -37.27792, -37.28442, -37.29021, -37.29523, -37.29943, 
        -37.30301, -37.30574, -37.30835, -37.31136, -37.31532, -37.32031, 
        -37.32619, -37.33228, -37.3379, -37.34241, -37.34529, -37.34642, 
        -37.34533, -37.34194, -37.33648, -37.32947, -37.32156, -37.31256, 
        -37.30504, -37.29824, -37.29245, -37.28764, -37.28405, -37.28215, 
        -37.28183, -37.28297, -37.28537, -37.28878, -37.293, -37.29765, 
        -37.30241, -37.3064, -37.30884, -37.30902, -37.30667, -37.30207, 
        -37.29558, -37.28745, -37.27766, -37.26655, -37.25435, -37.24096, 
        -37.22635, -37.21046, -37.19228, -37.17136, -37.14696, -37.11937, 
        -37.08852, -37.05432, -37.01687, -36.9764, -36.93321, -36.88803, 
        -36.84149,
  -29.29355, -29.33142, -29.371, -29.41208, -29.45396, -29.49649, 
        -29.53818, -29.58075, -29.62334, -29.66603, -29.70897, -29.75216, 
        -29.7956, -29.83969, -29.88455, -29.93011, -29.97598, -30.02187, 
        -30.06756, -30.11314, -30.15797, -30.20432, -30.25154, -30.29964, 
        -30.34854, -30.39809, -30.44822, -30.49832, -30.54793, -30.59628, 
        -30.64329, -30.68909, -30.73388, -30.77839, -30.82308, -30.86748, 
        -30.91408, -30.96207, -31.01126, -31.06086, -31.11011, -31.15777, 
        -31.20357, -31.24735, -31.28956, -31.33095, -31.37244, -31.41516, 
        -31.45942, -31.50584, -31.55314, -31.59993, -31.64706, -31.69296, 
        -31.73688, -31.77905, -31.81968, -31.85953, -31.89924, -31.93932, 
        -31.98067, -32.02334, -32.06744, -32.11276, -32.15929, -32.20634, 
        -32.25354, -32.29992, -32.34713, -32.39421, -32.44139, -32.48879, 
        -32.53685, -32.58602, -32.63663, -32.68912, -32.74334, -32.799, 
        -32.85493, -32.911, -32.96708, -33.02302, -33.07871, -33.13404, 
        -33.18747, -33.24067, -33.29274, -33.34363, -33.39433, -33.44488, 
        -33.49545, -33.54543, -33.59415, -33.64109, -33.68607, -33.72884, 
        -33.77023, -33.81029, -33.84939, -33.88824, -33.92686, -33.96527, 
        -34.00227, -34.03912, -34.07402, -34.1062, -34.1349, -34.16037, 
        -34.18278, -34.20277, -34.2205, -34.2367, -34.2515, -34.26517, 
        -34.27832, -34.29007, -34.30031, -34.3087, -34.31506, -34.3193, 
        -34.32215, -34.32384, -34.32357, -34.32458, -34.32591, -34.3277, 
        -34.32962, -34.33126, -34.33214, -34.33212, -34.33121, -34.32974, 
        -34.32832, -34.32779, -34.32919, -34.33317, -34.33969, -34.34818, 
        -34.35766, -34.36738, -34.37696, -34.38633, -34.39484, -34.40461, 
        -34.41513, -34.42698, -34.44079, -34.45687, -34.47502, -34.49475, 
        -34.51538, -34.53643, -34.55769, -34.5793, -34.60142, -34.62431, 
        -34.64758, -34.67061, -34.69303, -34.71474, -34.73513, -34.75479, 
        -34.77405, -34.79376, -34.81436, -34.83558, -34.85952, -34.88533, 
        -34.91271, -34.941, -34.9695, -34.99749, -35.0245, -35.05033, 
        -35.07573, -35.10163, -35.12883, -35.15786, -35.18891, -35.22164, 
        -35.25516, -35.28905, -35.32344, -35.35765, -35.39219, -35.42724, 
        -35.46331, -35.50092, -35.54037, -35.58203, -35.62499, -35.67155, 
        -35.72061, -35.7719, -35.82481, -35.87867, -35.93315, -35.98808, 
        -36.04333, -36.09863, -36.15349, -36.20727, -36.25906, -36.30844, 
        -36.35493, -36.39838, -36.43924, -36.47813, -36.51606, -36.55378, 
        -36.59176, -36.62979, -36.66732, -36.70372, -36.73844, -36.77122, 
        -36.80212, -36.83158, -36.85926, -36.88762, -36.91579, -36.94393, 
        -36.97153, -36.99812, -37.02338, -37.04736, -37.06989, -37.09107, 
        -37.11018, -37.12744, -37.14248, -37.15548, -37.16618, -37.17492, 
        -37.18219, -37.18863, -37.19458, -37.2007, -37.20733, -37.21439, 
        -37.22181, -37.22903, -37.23565, -37.24142, -37.2462, -37.25005, 
        -37.25331, -37.25564, -37.25803, -37.26105, -37.26512, -37.26945, 
        -37.27568, -37.28199, -37.28773, -37.29217, -37.29481, -37.29546, 
        -37.29388, -37.28991, -37.28389, -37.27632, -37.2679, -37.25952, 
        -37.25194, -37.24538, -37.2398, -37.23533, -37.23193, -37.23002, 
        -37.22948, -37.23036, -37.23244, -37.23553, -37.23944, -37.24396, 
        -37.2487, -37.25301, -37.25612, -37.25731, -37.25623, -37.2532, 
        -37.24847, -37.24226, -37.23452, -37.22527, -37.21456, -37.20248, 
        -37.18927, -37.17445, -37.15733, -37.13756, -37.11481, -37.08757, 
        -37.05851, -37.02598, -36.99025, -36.95152, -36.90978, -36.86572, 
        -36.81972 ;
    } // group puerto_rico_virgin_islands_geoid18
  } // group puerto_rico_virgin_islands_geoid18
}

netcdf GGXFspec-E6_no-data {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:content = "deviationsOfTheVertical" ;
		:title = "PRVI DOV 2018" ;
		:product_version = "2018" ;
		:summary = "PRVI hybrid deflection model. Deflections are at the Earth\'s surface" ;
		:source_file = "GGXFspec-E6_no-data.ggxf" ;
		:extent_description = "US Puerto Rico and Virgin Islands - onshore." ;
		:geospatial_lat_min = 17.67 ;
		:geospatial_lon_min = -65.09 ;
		:geospatial_lat_max = 18.42 ;
		:geospatial_lon_max = -64.6 ;
		:institution = "National Geodetic Survey, National Oceanic and Atmospheric Administration" ;
		:deliveryPoint = "1315 East West Hwy" ;
		:city = "Silver Spring" ;
		:postalCode = "20910" ;
		:country = "United States of America" ;
		:publisher_url = "https://geodesy.noaa.gov/PC_PROD/GEOID18/Format_ascii/g2018p0.asc.zip" ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:parameters.count = 2LL ;
		:parameters.0.parameterName = "deviationEast" ;
		:parameters.0.unitName = "arc-second" ;
		:parameters.0.unitSiRatio = 4.84813681109536e-06 ;
		:parameters.1.parameterName = "deviationNorth" ;
		:parameters.1.unitName = "arc-second" ;
		:parameters.1.unitSiRatio = 4.84813681109536e-06 ;
		:_NCProperties = "version=2,netcdf=4.9.0,hdf5=1.12.2" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: Puerto\ Rico\ Virgin\ Islands\ DEFLEC18 {

  // group attributes:
  		:interpolationMethod = "biquadratic" ;

  group: Puerto\ Rico\ Virgin\ Islands\ DEFLEC18 {
    dimensions:
    	iNodeCount = 361 ;
    	jNodeCount = 301 ;
    variables:
    	float deviationEast(iNodeCount, jNodeCount) ;
    		deviationEast:_Storage = "contiguous" ;
    		deviationEast:_Endianness = "little" ;
    	float deviationNorth(iNodeCount, jNodeCount) ;
    		deviationNorth:_Storage = "contiguous" ;
    		deviationNorth:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 15., 0.016666666666667, 0., -69., 0., 0.016666666666667 ;
    } // group Puerto\ Rico\ Virgin\ Islands\ DEFLEC18
  } // group Puerto\ Rico\ Virgin\ Islands\ DEFLEC18
}

netcdf GGXFspec-E3_grid-incomplete {
types:
  compound ggxfParameterType {
    char parameterName(32) ;
    char parameterSet(32) ;
    char unit(16) ;
    double unitSiRatio ;
    int sourceCrsAxis ;
    float parameterMinimumValue ;
    float parameterMaximumValue ;
    float noDataFlag ;
  }; // ggxfParameterType

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:title = "National Transformation v2_0" ;
		:summary = "Transformation of geodetic latitude and longitude referenced to NAD27 to latitude and longitude referenced to NAD83(Original)." ;
		:source_file = "27to83.gxt" ;
		:content = "geographic2dOffsets" ;
		:date_issued = "1995-02" ;
		:publisher_institution = "Geodetic Survey Division, Natural Resources Canada" ;
		:publisher_url = "https://webapp.geod.nrcan.gc.ca/geod/data-donnees/transformations.php" ;
		:license = "https://open.canada.ca/en/open-government-licence-canada" ;
		:geospatial_lat_min = 40. ;
		:geospatial_lon_min = -141. ;
		:geospatial_lat_max = 60. ;
		:geospatial_lon_max = -88. ;
		:extent_description = "Canada south of 60°N" ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:targetCrsWkt = "GEOGCRS[\"NAD83(Original)\",\n  DATUM[\"North American Datum 1983\",\n    ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:operationAccuracy = 1.5 ;
		ggxfParameterType :parameters = 
    {{"latitudeOffset"}, {"offset"}, {"arc-second"}, 4.84813681109536e-06, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"longitudeOffset"}, {"offset"}, {"arc-second"}, 4.84813681109536e-06, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"latitudeOffsetUncertainty"}, {"offsetUncertainty"}, {"metre"}, 1, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"longitudeOffsetUncertainty"}, {"offsetUncertainty"}, {"metre"}, 1, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38} ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: National\ Transformation\ v2_0 {
  dimensions:
  	offsetCount = 2 ;
  	offsetUncertaintyCount = 2 ;

  // group attributes:
  		:uncertaintyMeasure = "2CEE" ;
  		:interpolationMethod = "bilinear" ;

  group: CAwest {
    dimensions:
    	iNodeCount = 649 ;
    	jNodeCount = 157 ;
    variables:
    	float offset(jNodeCount, iNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.083333333333333, -142., 0.083333333333333, 0. ;
    		:gridPriority = 1LL ;
    } // group CAwest

  group: CAeast {
    dimensions:
    	iNodeCount = 529 ;
    	jNodeCount = 241 ;
    variables:
    	float offset(jNodeCount, iNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.083333333333333, -88., 0.083333333333333, 0. ;
    		:gridPriority = 2LL ;

    group: ONtronto {
      dimensions:
      	iNodeCount = 351 ;
      	jNodeCount = 511 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.666666667, 0., -0.00833333, -81.75, 0.1, 0.008333333 ;
      		:gridPriority = 1LL ;
      } // group ONtronto

    group: ONsarnia {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 121 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 43.41666667, 0., -0.00833333, -82.5833333, 0.1, 0.00083333 ;
      		:gridPriority = 2LL ;
      } // group ONsarnia

    group: ONwinsor {
      dimensions:
      	iNodeCount = 171 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 42.41666667, 0., -0.00833333, -83.1666667, 0.1, 0.00833333 ;
      		:gridPriority = 3LL ;
      } // group ONwinsor
    } // group CAeast
  } // group National\ Transformation\ v2_0
}

netcdf SAGeoid2010_Dataset {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:content = "geoidModel" ;
		:comment = "hybrid geoid" ;
		:title = "South_African_geoid_2010" ;
		:summary = "Model for converting ellipsoidal heights determined using NGI\'s TrigNet to orthometric heights on the South African Land Levelling Datum, to an accuracy of 10 cm (design requirements). Accuracy is 7cm absolute and relative <2cm + GNSS related error." ;
		:source_file = "SAGeoid2010_Dataset.ggxf" ;
		:geospatial_lat_min = -34.89 ;
		:geospatial_lon_min = 16.45 ;
		:geospatial_lat_max = -22.13 ;
		:geospatial_lon_max = 32.96 ;
		:extent_description = "South Africa - mainland onshore." ;
		:interpolationCrsWkt = "GEOGCRS[\"ITRF2005\",\n  DYNAMIC[FRAMEEPOCH[2000.0]],\n    DATUM[\"International Terrestrial Reference Frame 2005\",\n      ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"ITRF2005\",\n  DYNAMIC[FRAMEEPOCH[2000.0]],\n    TRF[\"International Terrestrial Reference Frame 2005\",\n      ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,3],\n  AXIS[\"Geodetic latitude (Lat)\",north,\n    ANGLEUNIT[\"degree\",0.0174532925199433]],\n  AXIS[\"Geodetic longitude (Lon)\",east,\n    ANGLEUNIT[\"degree\",0.0174532925199433]],\n  AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1]]]\n" ;
		:targetCrsWkt = "VERTCRS[\"VI LLD height\",\n  VDATUM[\"South Africa Land Levelling Datum\"],\n  CS[vertical,1],\n  AXIS[\"Gravity-related height (H)\",up],\n  LENGTHUNIT[\"metre\",1]]\n" ;
		:operationAccuracy = 0.07 ;
		:institution = "Chief Directorate: National Geospatial Information" ;
		:deliveryPoint = "Private Bag X10" ;
		:city = "Mowbray" ;
		:postalCode = "7705" ;
		:country = "South Africa" ;
		:publisher_url = "ftp://ftp.trignet.co.za/South_African_Geoid" ;
		:parameters.count = 1LL ;
		:parameters.0.parameterName = "geoidHeight" ;
		:parameters.0.sourceCrsAxis = 2LL ;
		:parameters.0.unitName = "metre" ;
		:parameters.0.unitSiRatio = 1. ;
		:_NCProperties = "version=2,netcdf=4.9.0,hdf5=1.12.2" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: SA\ geoid\ 2010 {

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: SA\ geoid\ 2010 {
    dimensions:
    	iNodeCount = 409 ;
    	jNodeCount = 313 ;
    variables:
    	float geoidHeight(jNodeCount, iNodeCount) ;
    		geoidHeight:_Storage = "contiguous" ;
    		geoidHeight:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -35., 0., 0.04166666666667, 16., 0.04166666666667, 0. ;
    } // group SA\ geoid\ 2010
  } // group SA\ geoid\ 2010
}

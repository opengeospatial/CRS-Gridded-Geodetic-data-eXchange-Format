netcdf ca_ntv2 {
types:
  compound ggxfParameterType {
    char parameterName(32) ;
    char parameterSet(32) ;
    char unit(16) ;
    double unitSiRatio ;
    int sourceCrsAxis ;
    float parameterMinimumValue ;
    float parameterMaximumValue ;
    float noDataFlag ;
  }; // ggxfParameterType

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "27to83.gxt" ;
		:title = "Canadian National NAD27-NAD83(Original) NTV2 transformation" ;
		:summary = "Canadian National NAD27-NAD83(Original) NTV2 transformation" ;
		:content = "geographic2dOffsets" ;
		:product_version = "National Transformation v2_0" ;
		:date_issued = "1995-02" ;
		:publisher_institution = "Geodetic Survey Division, Natural Resources Canada" ;
		:publisher_url = "https://webapp.geod.nrcan.gc.ca/geod/data-donnees/transformations.php" ;
		:license = "https://open.canada.ca/en/open-government-licence-canada" ;
		:geospatial_lat_min = 40. ;
		:geospatial_lon_min = -141. ;
		:geospatial_lat_max = 60. ;
		:geospatial_lon_max = -88. ;
		:extent_description = "Canada south of 60°N" ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:targetCrsWkt = "GEOGCRS[\"NAD83(Original)\",\n  DATUM[\"North American Datum 1983\",\n    ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		ggxfParameterType :parameters = 
    {{"latitudeOffset"}, {"offset"}, {"arc-second"}, 4.84813681109536e-06, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"longitudeOffset"}, {"offset"}, {"arc-second"}, 4.84813681109536e-06, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"latitudeOffsetUncertainty"}, {"offsetUncertainty"}, {"metre"}, 1, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"longitudeOffsetUncertainty"}, {"offsetUncertainty"}, {"metre"}, 1, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38} ;
		:operationAccuracy = 1.5 ;
		:uncertaintyMeasure = "2CEE" ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: national_transformation_v2_0 {
  dimensions:
  	offsetCount = 2 ;
  	offsetUncertaintyCount = 2 ;

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: CAeast {
    dimensions:
    	iNodeCount = 529 ;
    	jNodeCount = 241 ;
    variables:
    	float offset(jNodeCount, iNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.0833333333333333, -88., 0.0833333333333333, 0. ;
    		:iNodeCount = 529LL ;
    		:jNodeCount = 241LL ;
    		:gridPriority = 1LL ;

    group: NFstjohn {
      dimensions:
      	iNodeCount = 81 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 47.8333333333333, 0., -0.00833333333333333, -53., 0.00833333333333333, 0. ;
      		:iNodeCount = 81LL ;
      		:jNodeCount = 51LL ;
      		:gridPriority = 1LL ;
      } // group NFstjohn

    group: ONkinstn {
      dimensions:
      	iNodeCount = 321 ;
      	jNodeCount = 321 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.5, 0., -0.00833333333333333, -78.8333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 321LL ;
      		:jNodeCount = 321LL ;
      		:gridPriority = 2LL ;
      } // group ONkinstn

    group: ONottawa {
      dimensions:
      	iNodeCount = 221 ;
      	jNodeCount = 201 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 45.9166666666667, 0., -0.00833333333333333, -76.1666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 221LL ;
      		:jNodeCount = 201LL ;
      		:gridPriority = 3LL ;
      } // group ONottawa

    group: ONsarnia {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 121 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 43.4166666666667, 0., -0.00833333333333333, -82.5833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 101LL ;
      		:jNodeCount = 121LL ;
      		:gridPriority = 4LL ;
      } // group ONsarnia

    group: ONsault {
      dimensions:
      	iNodeCount = 351 ;
      	jNodeCount = 71 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.6666666666667, 0., -0.00833333333333333, -84.6666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 351LL ;
      		:jNodeCount = 71LL ;
      		:gridPriority = 5LL ;
      } // group ONsault

    group: ONtimins {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.6666666666667, 0., -0.00833333333333333, -81.6666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 101LL ;
      		:jNodeCount = 41LL ;
      		:gridPriority = 6LL ;
      } // group ONtimins

    group: ONtronto {
      dimensions:
      	iNodeCount = 351 ;
      	jNodeCount = 511 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.6666666666667, 0., -0.00833333333333333, -81.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 351LL ;
      		:jNodeCount = 511LL ;
      		:gridPriority = 7LL ;
      } // group ONtronto

    group: ONwinsor {
      dimensions:
      	iNodeCount = 171 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 42.4166666666667, 0., -0.00833333333333333, -83.1666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 171LL ;
      		:jNodeCount = 61LL ;
      		:gridPriority = 8LL ;
      } // group ONwinsor
    } // group CAeast

  group: CAwest {
    dimensions:
    	iNodeCount = 649 ;
    	jNodeCount = 157 ;
    variables:
    	float offset(jNodeCount, iNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.0833333333333333, -142., 0.0833333333333333, 0. ;
    		:iNodeCount = 649LL ;
    		:jNodeCount = 157LL ;
    		:gridPriority = 2LL ;

    group: ALbanff {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.25, 0., -0.00833333333333333, -115.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 1LL ;
      } // group ALbanff

    group: ALbarhed {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.1666666666667, 0., -0.00833333333333333, -114.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 2LL ;
      } // group ALbarhed

    group: ALbonvil {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.3333333333333, 0., -0.00833333333333333, -110.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 3LL ;
      } // group ALbonvil

    group: ALbowisl {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -111.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 4LL ;
      } // group ALbowisl

    group: ALbrooks {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.6666666666667, 0., -0.00833333333333333, -112., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 5LL ;
      } // group ALbrooks

    group: ALcalgry {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 101 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.3333333333333, 0., -0.00833333333333333, -114.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 101LL ;
      		:jNodeCount = 101LL ;
      		:gridPriority = 6LL ;
      } // group ALcalgry

    group: ALcamros {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.0833333333333, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 7LL ;
      } // group ALcamros

    group: ALcanmor {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.1666666666667, 0., -0.00833333333333333, -115.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 8LL ;
      } // group ALcanmor

    group: ALcardst {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -113.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 9LL ;
      } // group ALcardst

    group: ALcarsta {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.6666666666667, 0., -0.00833333333333333, -114.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 10LL ;
      } // group ALcarsta

    group: ALclarho {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -113.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 11LL ;
      } // group ALclarho

    group: ALcoldlk {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.5833333333333, 0., -0.00833333333333333, -110.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 12LL ;
      } // group ALcoldlk

    group: ALcrowps {
      dimensions:
      	iNodeCount = 71 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.75, 0., -0.00833333333333333, -114.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 71LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 13LL ;
      } // group ALcrowps

    group: ALdraytn {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -115.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 14LL ;
      } // group ALdraytn

    group: ALdrumhl {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.5833333333333, 0., -0.00833333333333333, -112.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 41LL ;
      		:gridPriority = 15LL ;
      } // group ALdrumhl

    group: ALedmntn {
      dimensions:
      	iNodeCount = 131 ;
      	jNodeCount = 91 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.9166666666667, 0., -0.00833333333333333, -114.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 131LL ;
      		:jNodeCount = 91LL ;
      		:gridPriority = 16LL ;
      } // group ALedmntn

    group: ALedson {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.6666666666667, 0., -0.00833333333333333, -116.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 17LL ;
      } // group ALedson

    group: ALfairvw {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.1666666666667, 0., -0.00833333333333333, -118.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 18LL ;
      } // group ALfairvw

    group: ALftmacl {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.8333333333333, 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 19LL ;
      } // group ALftmacl

    group: ALftmcmr {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.8333333333333, 0., -0.00833333333333333, -111.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 20LL ;
      } // group ALftmcmr

    group: ALgrcach {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54., 0., -0.00833333333333333, -119.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 21LL ;
      } // group ALgrcach

    group: ALgrimsh {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.25, 0., -0.00833333333333333, -117.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 22LL ;
      } // group ALgrimsh

    group: ALgrprar {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.25, 0., -0.00833333333333333, -118.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 23LL ;
      } // group ALgrprar

    group: ALhanna {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.75, 0., -0.00833333333333333, -112.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 24LL ;
      } // group ALhanna

    group: ALhilevl {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 58.5833333333333, 0., -0.00833333333333333, -117.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 25LL ;
      } // group ALhilevl

    group: ALhinton {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.5, 0., -0.00833333333333333, -117.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 26LL ;
      } // group ALhinton

    group: ALhiprai {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.5, 0., -0.00833333333333333, -116.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 27LL ;
      } // group ALhiprai

    group: ALinnsfl {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.1666666666667, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 28LL ;
      } // group ALinnsfl

    group: ALjasper {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -118.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 29LL ;
      } // group ALjasper

    group: ALlacbic {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.8333333333333, 0., -0.00833333333333333, -112.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 30LL ;
      } // group ALlacbic

    group: ALlacomb {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.5833333333333, 0., -0.00833333333333333, -113.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 31LL ;
      } // group ALlacomb

    group: ALletbrg {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 41LL ;
      		:gridPriority = 32LL ;
      } // group ALletbrg

    group: ALlkloui {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.5, 0., -0.00833333333333333, -116.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 33LL ;
      } // group ALlkloui

    group: ALlydmin {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -110.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 34LL ;
      } // group ALlydmin

    group: ALmedhat {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.1666666666667, 0., -0.00833333333333333, -110.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 35LL ;
      } // group ALmedhat

    group: ALolds {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.9166666666667, 0., -0.00833333333333333, -114.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 36LL ;
      } // group ALolds

    group: ALoyen {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.4166666666667, 0., -0.00833333333333333, -110.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 37LL ;
      } // group ALoyen

    group: ALpeacer {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.3333333333333, 0., -0.00833333333333333, -117.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 38LL ;
      } // group ALpeacer

    group: ALpinchr {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 39LL ;
      } // group ALpinchr

    group: ALponoka {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.75, 0., -0.00833333333333333, -113.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 40LL ;
      } // group ALponoka

    group: ALraymnd {
      dimensions:
      	iNodeCount = 51 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      		:iNodeCount = 51LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 41LL ;
      } // group ALraymnd

    group: ALredeer {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.4166666666667, 0., -0.00833333333333333, -113.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 42LL ;
      } // group ALredeer

    group: ALrockmt {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.5, 0., -0.00833333333333333, -115., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 43LL ;
      } // group ALrockmt

    group: ALslavlk {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.3333333333333, 0., -0.00833333333333333, -114.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 44LL ;
      } // group ALslavlk

    group: ALstetlr {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.4166666666667, 0., -0.00833333333333333, -112.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 45LL ;
      } // group ALstetlr

    group: ALstpaul {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.0833333333333, 0., -0.00833333333333333, -111.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 46LL ;
      } // group ALstpaul

    group: ALstramr {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.1666666666667, 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 47LL ;
      } // group ALstramr

    group: ALswanhi {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.8333333333333, 0., -0.00833333333333333, -115.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 48LL ;
      } // group ALswanhi

    group: ALtaber {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -112.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 49LL ;
      } // group ALtaber

    group: ALtrehil {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.75, 0., -0.00833333333333333, -113.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 50LL ;
      } // group ALtrehil

    group: ALvegvil {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.5833333333333, 0., -0.00833333333333333, -112.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 51LL ;
      } // group ALvegvil

    group: ALvermil {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.4166666666667, 0., -0.00833333333333333, -111., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 52LL ;
      } // group ALvermil

    group: ALwanwgt {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -111., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 53LL ;
      } // group ALwanwgt

    group: ALweslok {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.25, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 54LL ;
      } // group ALweslok

    group: ALwetask {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53., 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 55LL ;
      } // group ALwetask

    group: ALwhitec {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.1666666666667, 0., -0.00833333333333333, -115.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 56LL ;
      } // group ALwhitec

    group: BCcambel {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -125.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 57LL ;
      } // group BCcambel

    group: BCcranbk {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -115.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 58LL ;
      } // group BCcranbk

    group: BCdawson {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.8333333333333, 0., -0.00833333333333333, -120.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 59LL ;
      } // group BCdawson

    group: BCelkfrd {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -115., 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 60LL ;
      } // group BCelkfrd

    group: BCfield {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.4166666666667, 0., -0.00833333333333333, -116.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 61LL ;
      } // group BCfield

    group: BCgranil {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.9166666666667, 0., -0.00833333333333333, -126.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 62LL ;
      } // group BCgranil

    group: BCkamlop {
      dimensions:
      	iNodeCount = 51 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.75, 0., -0.00833333333333333, -120.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 51LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 63LL ;
      } // group BCkamlop

    group: BCkelwna {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -119.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 64LL ;
      } // group BCkelwna

    group: BClogan {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5, 0., -0.00833333333333333, -120.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 65LL ;
      } // group BClogan

    group: BCmacknz {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.4166666666667, 0., -0.00833333333333333, -123.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 66LL ;
      } // group BCmacknz

    group: BCnanimo {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -124.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 61LL ;
      		:gridPriority = 67LL ;
      } // group BCnanimo

    group: BCnelson {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -117.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 68LL ;
      } // group BCnelson

    group: BCparkvl {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.3333333333333, 0., -0.00833333333333333, -124.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 69LL ;
      } // group BCparkvl

    group: BCpentic {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -119.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 70LL ;
      } // group BCpentic

    group: BCportal {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.3333333333333, 0., -0.00833333333333333, -124.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 71LL ;
      } // group BCportal

    group: BCpowell {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -124.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 72LL ;
      } // group BCpowell

    group: BCprigeo {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.0833333333333, 0., -0.00833333333333333, -122.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 41LL ;
      		:gridPriority = 73LL ;
      } // group BCprigeo

    group: BCroslnd {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.0833333333333, 0., -0.00833333333333333, -117.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 74LL ;
      } // group BCroslnd

    group: BCtrail {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.1666666666667, 0., -0.00833333333333333, -117.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 75LL ;
      } // group BCtrail

    group: BCtumblr {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.1666666666667, 0., -0.00833333333333333, -121.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 76LL ;
      } // group BCtumblr

    group: BCvancvr {
      dimensions:
      	iNodeCount = 131 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.4166666666667, 0., -0.00833333333333333, -123.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 131LL ;
      		:jNodeCount = 51LL ;
      		:gridPriority = 77LL ;
      } // group BCvancvr

    group: BCvernon {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.3333333333333, 0., -0.00833333333333333, -119.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 78LL ;
      } // group BCvernon

    group: BCvictor {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.75, 0., -0.00833333333333333, -123.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 51LL ;
      		:gridPriority = 79LL ;
      } // group BCvictor

    group: ONthundr {
      dimensions:
      	iNodeCount = 71 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.5833333333333, 0., -0.00833333333333333, -89.5833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 71LL ;
      		:jNodeCount = 51LL ;
      		:gridPriority = 80LL ;
      } // group ONthundr

    group: SAestvan {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -103.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 81LL ;
      } // group SAestvan

    group: SAmelfrt {
      dimensions:
      	iNodeCount = 71 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -104.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 71LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 82LL ;
      } // group SAmelfrt

    group: SAmelvil {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51., 0., -0.00833333333333333, -102.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 83LL ;
      } // group SAmelvil

    group: SAmosjaw {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5, 0., -0.00833333333333333, -105.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 84LL ;
      } // group SAmosjaw

    group: SAnbatle {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.8333333333333, 0., -0.00833333333333333, -108.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 85LL ;
      } // group SAnbatle

    group: SApralbt {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -106., 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 86LL ;
      } // group SApralbt

    group: SAregina {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5833333333333, 0., -0.00833333333333333, -104.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 87LL ;
      } // group SAregina

    group: SAsatoon {
      dimensions:
      	iNodeCount = 51 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.25, 0., -0.00833333333333333, -106.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 51LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 88LL ;
      } // group SAsatoon

    group: SAswiftc {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.4166666666667, 0., -0.00833333333333333, -107.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 89LL ;
      } // group SAswiftc

    group: SAweybrn {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.75, 0., -0.00833333333333333, -103.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 90LL ;
      } // group SAweybrn

    group: SAyorktn {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.3333333333333, 0., -0.00833333333333333, -102.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 91LL ;
      } // group SAyorktn
    } // group CAwest

  group: CAnorth {
    dimensions:
    	iNodeCount = 589 ;
    	jNodeCount = 181 ;
    variables:
    	float offset(jNodeCount, iNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 75., 0., -0.0833333333333333, -142., 0.166666666666667, 0. ;
    		:iNodeCount = 589LL ;
    		:jNodeCount = 181LL ;
    		:gridPriority = 3LL ;

    group: NWclyder {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 70.5833333333333, 0., -0.00833333333333333, -68.8333333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      		:gridPriority = 1LL ;
      } // group NWclyder

    group: NWftgood {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 66.3333333333333, 0., -0.00833333333333333, -128.833333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 2LL ;
      } // group NWftgood

    group: NWhayriv {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 61., 0., -0.00833333333333333, -116.5, 0.0166666666666667, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 61LL ;
      		:gridPriority = 3LL ;
      } // group NWhayriv

    group: NWinuvik {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 68.5, 0., -0.00833333333333333, -133.833333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 41LL ;
      		:gridPriority = 4LL ;
      } // group NWinuvik

    group: NWiqulit {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 64., 0., -0.00833333333333333, -69., 0.0166666666666667, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 61LL ;
      		:gridPriority = 5LL ;
      } // group NWiqulit

    group: NWpondin {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 72.75, 0., -0.00833333333333333, -78.1666666666667, 0.0166666666666667, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 6LL ;
      } // group NWpondin

    group: NWrankin {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.9166666666667, 0., -0.00833333333333333, -92.1666666666667, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 7LL ;
      } // group NWrankin

    group: NWyellow {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.5, 0., -0.00833333333333333, -114.5, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 8LL ;
      } // group NWyellow

    group: YUdawson {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 64.1666666666667, 0., -0.00833333333333333, -139.5, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 9LL ;
      } // group YUdawson

    group: YUrossri {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.0833333333333, 0., -0.00833333333333333, -132.583333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      		:gridPriority = 10LL ;
      } // group YUrossri

    group: YUwhiteh {
      dimensions:
      	iNodeCount = 6 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(jNodeCount, iNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 60.75, 0., -0.00833333333333333, -135.083333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 6LL ;
      		:jNodeCount = 11LL ;
      		:gridPriority = 11LL ;
      } // group YUwhiteh
    } // group CAnorth

  group: CAarctic {
    dimensions:
    	iNodeCount = 295 ;
    	jNodeCount = 109 ;
    variables:
    	float offset(jNodeCount, iNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(jNodeCount, iNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 84., 0., -0.0833333333333333, -142., 0.333333333333333, 0. ;
    		:iNodeCount = 295LL ;
    		:jNodeCount = 109LL ;
    		:gridPriority = 4LL ;
    } // group CAarctic
  } // group national_transformation_v2_0
}

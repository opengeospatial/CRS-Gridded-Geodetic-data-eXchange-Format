netcdf def_packed {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "nz_linz_nzgd2000-20180701.yaml" ;
		:product_version = "20180701" ;
		:content = "deformationModel" ;
		:title = "New Zealand Deformation Model." ;
		:summary = "Defines the secular model (National Deformation Model)\nand patches for significant deformation events since 2000.\n" ;
		:institution = "Land Information New Zealand" ;
		:deliveryPoint = "Level 7, Radio New Zealand House\n155 The Terrace\nPO Box 5501\n" ;
		:city = "Wellington" ;
		:postalCode = "6145" ;
		:creator_email = "customersupport@linz.govt.nz" ;
		:publisher_url = "https://www.linz.govt.nz/nzgd2000" ;
		:date_issued = "2018-07-01" ;
		:extent_description = "New Zealand EEZ" ;
		:geospatial_lat_min = -55.94 ;
		:geospatial_lon_min = 160.62 ;
		:geospatial_lat_max = -25.89 ;
		:geospatial_lon_max = -171.23 ;
		:start_date = "1900-01-01" ;
		:end_date = "2050-01-01" ;
		:sourceCrsWkt = "GEOGCRS[\"NZGD2000\",DATUM[\"New Zealand Geodetic Datum 2000\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6167]],CS[ellipsoidal,3,ID[\"EPSG\",6423]],AXIS[\"Geodetic latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Geodetic longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],ID[\"EPSG\",4959]]" ;
		:targetCrsWkt = "GEOGCRS[\"ITRF96\", DYNAMIC[FRAMEEPOCH[1997.0]],DATUM[\"International Terrestrial Reference Frame 1996\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6654]],CS[ellipsoidal,3,ID[\"EPSG\",6423]],AXIS[\"Geodetic latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Geodetic longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],ID[\"EPSG\",7907]]" ;
		:interpolationCrsWkt = "GEOGCRS[\"NZGD2000\",DATUM[\"New Zealand Geodetic Datum 2000\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6167]],CS[ellipsoidal,2,ID[\"EPSG\",6422]],AXIS[\"Geodetic latitude (Lat)\",north],AXIS[\"Geodetic longitude (Lon)\",east],ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]],ID[\"EPSG\",4167]]" ;
		:parameters.count = 5LL ;
		:parameters.0.parameterName = "displacementEast" ;
		:parameters.0.parameterSet = "displacement" ;
		:parameters.0.unit = "metre" ;
		:parameters.0.unitSiRatio = 1. ;
		:parameters.0.sourceCrsAxis = 1LL ;
		:parameters.0.noDataFlag = 9999. ;
		:parameters.1.parameterName = "displacementNorth" ;
		:parameters.1.parameterSet = "displacement" ;
		:parameters.1.unit = "metre" ;
		:parameters.1.unitSiRatio = 1. ;
		:parameters.1.sourceCrsAxis = 0LL ;
		:parameters.1.noDataFlag = 9999. ;
		:parameters.2.parameterName = "displacementUp" ;
		:parameters.2.parameterSet = "displacement" ;
		:parameters.2.unit = "metre" ;
		:parameters.2.unitSiRatio = 1. ;
		:parameters.2.sourceCrsAxis = 2LL ;
		:parameters.2.noDataFlag = 9999. ;
		:parameters.3.parameterName = "displacementHorizontalUncertainty" ;
		:parameters.3.parameterSet = "displacementUncertainty" ;
		:parameters.3.unit = "metre" ;
		:parameters.3.unitSiRatio = 1. ;
		:parameters.3.uncertaintyMeasure = "2CEP" ;
		:parameters.3.defaultValue = 0.01 ;
		:parameters.3.noDataFlag = 999. ;
		:parameters.4.parameterName = "displacementUpUncertainty" ;
		:parameters.4.parameterSet = "displacementUncertainty" ;
		:parameters.4.unit = "metre" ;
		:parameters.4.unitSiRatio = 1. ;
		:parameters.4.uncertaintyMeasure = "2SE" ;
		:parameters.4.defaultValue = 0.02 ;
		:parameters.4.noDataFlag = 999. ;
		:operationAccuracy = 0.01 ;
		:_NCProperties = "version=2,netcdf=4.9.0,hdf5=1.12.2" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: secular-vertical-velocity {

  // group attributes:
  		:interpolationMethod = "bilinear" ;
  		:gridParameters = "displacementUp" ;
  		:constantParameters.count = 1LL ;
  		:constantParameters.0.parameterName = "displacementUpUncertainty" ;
  		:constantParameters.0.parameterValue = 0.001 ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "velocity" ;
  		:timeFunctions.0.functionReferenceDate = "2000-01-01T00:00:00Z" ;

  group: national-vertical-velocity-grid {
    dimensions:
    	iNodeCount = 3 ;
    	jNodeCount = 4 ;
    variables:
    	short displacement(jNodeCount, iNodeCount) ;
    		displacement:add_offset = 0.33 ;
    		displacement:scale_factor = 0.01 ;
    		displacement:missing_value = 32767s ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 172.6, 0.6, 0., -41.6, 0., 0.4 ;
    data:

     displacement =
  11, 41, 31,
  -21, 9, -1,
  -38, -8, -18,
  -41, -11, 32767 ;
    } // group national-vertical-velocity-grid
  } // group secular-vertical-velocity

group: co-and-post-seismic-deformation {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Hypothetical earthquake" ;
  		:interpolationMethod = "bilinear" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1.05 ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 0.29 ;

  group: far-field-deformation-grid {
    dimensions:
    	iNodeCount = 5 ;
    	jNodeCount = 6 ;
    variables:
    	short displacement(jNodeCount, iNodeCount, displacementCount) ;
    		displacement:add_offset = -0.44 ;
    		displacement:scale_factor = 0.01 ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 172.6, 0.6, 0., -41.6, 0., 0.4 ;
    data:

     displacement =
  168, -164, -196,
  228, -144, -178,
  248, -124, -161,
  228, -104, -143,
  168, -84, -126,
  150, -220, -86,
  210, -200, -68,
  230, -180, -51,
  210, -160, -33,
  150, -140, -16,
  132, -248, -14,
  192, -228, 3,
  212, -208, 21,
  192, -188, 38,
  132, -168, 56,
  114, -246, 19,
  174, -226, 37,
  194, -206, 54,
  174, -186, 72,
  114, -166, 89,
  96, -216, 14,
  156, -196, 31,
  176, -176, 49,
  156, -156, 66,
  96, -136, 84,
  78, -156, -30,
  138, -136, -12,
  158, -116, 5,
  138, -96, 23,
  78, -76, 40 ;

    group: near-field-deformation-grid {
      dimensions:
      	iNodeCount = 5 ;
      	jNodeCount = 3 ;
      variables:
      	short displacement(jNodeCount, iNodeCount, displacementCount) ;
      		displacement:add_offset = -0.53 ;
      		displacement:scale_factor = 0.01 ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 172.6, 0.3, 0., -41.2, 0., 0.2 ;
      data:

       displacement =
  201, -219, 12,
  216, -209, 21,
  221, -199, 30,
  216, -189, 39,
  201, -179, 47,
  192, -221, 34,
  207, -211, 42,
  212, -201, 51,
  207, -191, 60,
  192, -181, 69,
  183, -217, 45,
  198, -207, 54,
  203, -197, 63,
  198, -187, 72,
  183, -177, 80 ;
      } // group near-field-deformation-grid
    } // group far-field-deformation-grid
  } // group co-and-post-seismic-deformation
}

netcdf GGXFspec-E1_parameterSet-removed {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:title = "Catalino Canyon transformation version 2022-06" ;
		:summary = "Example transformation constructed for purposes of illustration." ;
		:source_file = "Catalano_Canyon.yaml" ;
		:content = "geographic2dOffsets" ;
		:extent_description = "Italy - Mediterranean Sea west of Sardinia - Catalano Canyon." ;
		:geospatial_lat_min = 39.9 ;
		:geospatial_lon_min = 7.6 ;
		:geospatial_lat_max = 40.15 ;
		:geospatial_lon_max = 7.87 ;
		:geospatial_bounds = "Polygon(( 40.09, 7.72, 40.12, 7.71, 39.92, 7.84, 39.93, 7.64, 40.05, 7.64, 40.09, 7.72 ))" ;
		:interpolationCrsWkt = "GEOGCRS[\"ED50\",\n  DATUM[\"European Datum 1950\",\n    ELLIPSOID[\"International 1924\",6378388,297,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"ED50\",\n  DATUM[\"European Datum 1950\",\n    ELLIPSOID[\"International 1924\",6378388,297,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:targetCrsWkt = "GEOGCRS[\"ETRF2000\",\n  DATUM[\"European Terrestrial Reference Frame 2000\",\n    ELLIPSOID[\"GRS 1980\",6378137,298.257222101,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:operationAccuracy = 2LL ;
		:parameters.count = 2LL ;
		:parameters.0.parameterName = "latitudeOffset" ;
		:parameters.0.sourceCrsAxis = 0LL ;
		:parameters.0.unit = "arc-second" ;
		:parameters.0.unitSiRatio = 4.84813681109536e-06 ;
		:parameters.1.parameterName = "longitudeOffset" ;
		:parameters.1.sourceCrsAxis = 1LL ;
		:parameters.1.unit = "arc-second" ;
		:parameters.1.unitSiRatio = 4.84813681109536e-06 ;
		:_NCProperties = "version=2,netcdf=4.9.0,hdf5=1.12.2" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: Catalano_Canyon {

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: South {
    dimensions:
    	iNodeCount = 5 ;
    	jNodeCount = 3 ;
    variables:
    	float latitudeOffset(jNodeCount, iNodeCount) ;
    		latitudeOffset:_Storage = "contiguous" ;
    		latitudeOffset:_Endianness = "little" ;
    	float longitudeOffset(jNodeCount, iNodeCount) ;
    		longitudeOffset:_Storage = "contiguous" ;
    		longitudeOffset:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 40., 0., -0.05, 7.6, 0.0666666666666667, 0. ;
    } // group South

  group: North {
    dimensions:
    	iNodeCount = 3 ;
    	jNodeCount = 4 ;
    variables:
    	float latitudeOffset(jNodeCount, iNodeCount) ;
    		latitudeOffset:_Storage = "contiguous" ;
    		latitudeOffset:_Endianness = "little" ;
    	float longitudeOffset(jNodeCount, iNodeCount) ;
    		longitudeOffset:_Storage = "contiguous" ;
    		longitudeOffset:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 40.15, 0., -0.05, 7.6, 0.1, 0. ;
    } // group North
  } // group Catalano_Canyon
}

netcdf test_geoid {
types:
  compound ggxfParameterType {
    char parameterName(32) ;
    char parameterSet(32) ;
    char unit(16) ;
    double unitSiRatio ;
    int sourceCrsAxis ;
    float parameterMinimumValue ;
    float parameterMaximumValue ;
    float noDataFlag ;
  }; // ggxfParameterType

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "tiny_geoid.gxt" ;
		:content = "geoidModel" ;
		:title = "hybrid geoid" ;
		:summary = "Tiny geoid for testing GGXF implementation" ;
		:geospatial_lat_min = 22.5 ;
		:geospatial_lon_min = -69. ;
		:geospatial_lat_max = 24.6 ;
		:geospatial_lon_max = -67. ;
		:extent_description = "Tiny example geoid." ;
		:interpolationCrsWkt = "GEOGCRS[\"WGS 84 (G2139)\", \n  DYNAMIC[FRAMEEPOCH[2016.0]],\n  DATUM[\"World Geodetic System 1984 (G2139)\",ELLIPSOID[\"WGS 84\",6378137,298.257223563,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7030]],ID[\"EPSG\",1309]],\n  CS[ellipsoidal,3,ID[\"EPSG\",6423]],\n    AXIS[\"latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],\n    AXIS[\"longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],\n    AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]]\n  ,ID[\"EPSG\",9754]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"WGS 84 (G2139)\", \n  DYNAMIC[FRAMEEPOCH[2016.0]],\n  DATUM[\"World Geodetic System 1984 (G2139)\",ELLIPSOID[\"WGS 84\",6378137,298.257223563,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7030]],ID[\"EPSG\",1309]],\n  CS[ellipsoidal,3,ID[\"EPSG\",6423]],\n    AXIS[\"latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],\n    AXIS[\"longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],\n    AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]]\n  ,ID[\"EPSG\",9754]]\n" ;
		:targetCrsWkt = "VERTCRS[\"Vertical datum height\",\n VDATUM[\"Imaginary vertical datum\",ID[\"EPSG\",1124]],\n CS[vertical,1,ID[\"EPSG\",6499]],\n   AXIS[\"Gravity-related height (H)\",up],LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]\n ,ID[\"EPSG\",6642]]    \n" ;
		ggxfParameterType :parameters = 
    {{"geoidHeight"}, {"geoidHeight"}, {"metre"}, 1, 2, -3.402823e+38, -3.402823e+38, -3.402823e+38} ;
		:operationAccuracy = 0.015 ;
		:organisationName = "A Hypothetical National Geodetic Survey." ;
		:deliveryPoint = "Somewhere" ;
		:city = "A city" ;
		:postalCode = "99999" ;
		:country = "United States of America" ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: default {

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: geoid_grid {
    dimensions:
    	iNodeCount = 3 ;
    	jNodeCount = 4 ;
    variables:
    	float geoidHeight(jNodeCount, iNodeCount) ;
    		geoidHeight:_Storage = "contiguous" ;
    		geoidHeight:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 22.5, 0., 0.7, -69., 1., 0. ;
    		:gridPriority = 1LL ;
    data:

     geoidHeight =
  -10.5, -20.5, -30.5,
  -11.5, -21.5, -31.5,
  -12.5, -22.5, -32.5,
  -13.5, -23.5, -33.5 ;
    } // group geoid_grid
  } // group default
}

netcdf nzgd2000-20180701 {
types:
  compound ggxfParameterType {
    char parameterName(32) ;
    char parameterSet(32) ;
    char unitName(16) ;
    float unitSiRatio ;
    int sourceCrsAxis ;
    float parameterMinimumValue ;
    float parameterMaximumValue ;
    float noDataFlag ;
  }; // ggxfParameterType

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "nzgd2000-20180701.yaml" ;
		:product_version = "20180701" ;
		:content = "deformationModel" ;
		:title = "New Zealand Deformation Model." ;
		:summary = "Defines the secular model (National Deformation Model)\nand patches for significant deformation events since 2000.\n" ;
		:publisher_institution = "Land Information New Zealand" ;
		:deliveryPoint = "Level 7, Radio New Zealand House\n155 The Terrace\nPO Box 5501\n" ;
		:city = "Wellington" ;
		:postalCode = "6145" ;
		:creator_email = "customersupport@linz.govt.nz" ;
		:publisher_url = "https://www.linz.govt.nz/nzgd2000" ;
		:date_issued = "2018-07-01" ;
		:extent_description = "New Zealand EEZ" ;
		:geospatial_lat_min = -55.94 ;
		:geospatial_lon_min = 160.62 ;
		:geospatial_lat_max = -25.89 ;
		:geospatial_lon_max = -171.23 ;
		:start_date = "1900-01-01" ;
		:end_date = "2050-01-01" ;
		:geospatial_bounds = "<gml:Polygon srsName=\"EPSG:4167\">\n  <gml:exterior>\n    <gml:LinearRing>\n      <gml:posList>-32.42 168.65 -34.98 168.10 -37.58 170.07 -40.60 167.30 -44.32 162.17 -51.17 160.62 -54.97 165.11 -55.94 168.78 -54.70 173.54 -53.26 174.64 -51.66 174.48 -53.04 178.46 -51.94 182.69 -50.45 183.84 -47.76 184.00 -46.81 187.31 -44.68 188.77 -42.93 188.53 -41.50 187.23 -40.26 182.07 -36.91 182.64 -34.59 180.22 -34.45 182.66 -33.12 184.50 -29.73 185.92 -27.47 185.34 -25.89 182.29 -27.22 179.01 -31.55 177.28 -34.32 179.37 -30.85 172.97 -30.88 171.22 -32.42 168.65</gml:posList>\n    </gml:LinearRing>\n  </gml:exterior>\n</gml:Polygon>\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NZGD2000\",DATUM[\"New Zealand Geodetic Datum 2000\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6167]],CS[ellipsoidal,3,ID[\"EPSG\",6423]],AXIS[\"Geodetic latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Geodetic longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],ID[\"EPSG\",4959]]" ;
		:targetCrsWkt = "GEOGCRS[\"ITRF96\", DYNAMIC[FRAMEEPOCH[1997.0]],DATUM[\"International Terrestrial Reference Frame 1996\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6654]],CS[ellipsoidal,3,ID[\"EPSG\",6423]],AXIS[\"Geodetic latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Geodetic longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],ID[\"EPSG\",7907]]" ;
		:interpolationCrsWkt = "GEOGCRS[\"NZGD2000\",DATUM[\"New Zealand Geodetic Datum 2000\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6167]],CS[ellipsoidal,2,ID[\"EPSG\",6422]],AXIS[\"Geodetic latitude (Lat)\",north],AXIS[\"Geodetic longitude (Lon)\",east],ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]],ID[\"EPSG\",4167]]" ;
		ggxfParameterType :parameters = 
    {{"displacementEast"}, {"displacement"}, {"metre"}, 1, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"displacementNorth"}, {"displacement"}, {"metre"}, 1, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"displacementUp"}, {"displacement"}, {"metre"}, 1, 2, -3.402823e+38, -3.402823e+38, -3.402823e+38} ;
		:operationAccuracy = 0.01 ;
		:uncertaintyMeasure = "2CEP 2SE" ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: nz_linz_nzgd2000-ndm-grid02 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Secular deformation model derived from NUVEL-1A rotation rates\nSecular deformation model derived from GNS model 2011 V4\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "velocity" ;
  		:timeFunctions.1.functionReferenceDate = "2000-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: ndm_grid_nuvel1a_eez {
    dimensions:
    	gridi = 73 ;
    	gridj = 67 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -25., 0., -0.5, 158., 0.5, 0. ;
    		:iNodeCount = 73LL ;
    		:jNodeCount = 67LL ;

    group: ndm_grid_igns2011_nz {
      dimensions:
      	gridi = 141 ;
      	gridj = 151 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -33., 0., -0.1, 165.5, 0.1, 0. ;
      		:iNodeCount = 141LL ;
      		:jNodeCount = 151LL ;
      } // group ndm_grid_igns2011_nz
    } // group ndm_grid_nuvel1a_eez
  } // group nz_linz_nzgd2000-ndm-grid02

group: nz_linz_nzgd2000-si20030821-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Secretary Island (Fiordland) earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2003-08-21T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2004-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_si_20030821_grid_si_l1 {
    dimensions:
    	gridi = 44 ;
    	gridj = 34 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -43.5, 0., -0.125, 165.85, 0.15, 0. ;
    		:iNodeCount = 44LL ;
    		:jNodeCount = 34LL ;

    group: patch_si_20030821_grid_si_l2 {
      dimensions:
      	gridi = 47 ;
      	gridj = 45 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -44.5, 0., -0.03125, 166.225, 0.0375, 0. ;
      		:iNodeCount = 47LL ;
      		:jNodeCount = 45LL ;

      group: patch_si_20030821_grid_si_l3 {
        dimensions:
        	gridi = 93 ;
        	gridj = 81 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -44.828125, 0., -0.0078125, 166.5625, 0.009375, 0. ;
        		:iNodeCount = 93LL ;
        		:jNodeCount = 81LL ;
        } // group patch_si_20030821_grid_si_l3
      } // group patch_si_20030821_grid_si_l2
    } // group patch_si_20030821_grid_si_l1
  } // group nz_linz_nzgd2000-si20030821-grid01

group: nz_linz_nzgd2000-mq20041223-grid011 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p0_l1 {
    dimensions:
    	gridi = 10 ;
    	gridj = 8 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -52.125, 0., -0.125, 168.4, 0.15, 0. ;
    		:iNodeCount = 10LL ;
    		:jNodeCount = 8LL ;
    } // group patch_mq_20041223_grid_mq_p0_l1
  } // group nz_linz_nzgd2000-mq20041223-grid011

group: nz_linz_nzgd2000-mq20041223-grid012 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p1_sl2 {
    dimensions:
    	gridi = 105 ;
    	gridj = 137 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -48.25, 0., -0.03125, 158.8, 0.0375, 0. ;
    		:iNodeCount = 105LL ;
    		:jNodeCount = 137LL ;
    } // group patch_mq_20041223_grid_mq_p1_sl2
  } // group nz_linz_nzgd2000-mq20041223-grid012

group: nz_linz_nzgd2000-mq20041223-grid013 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p2_l1 {
    dimensions:
    	gridi = 11 ;
    	gridj = 11 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -50.125, 0., -0.125, 165.4, 0.15, 0. ;
    		:iNodeCount = 11LL ;
    		:jNodeCount = 11LL ;
    } // group patch_mq_20041223_grid_mq_p2_l1
  } // group nz_linz_nzgd2000-mq20041223-grid013

group: nz_linz_nzgd2000-mq20041223-grid014 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p3_l1 {
    dimensions:
    	gridi = 9 ;
    	gridj = 8 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -49.25, 0., -0.125, 178.15, 0.15, 0. ;
    		:iNodeCount = 9LL ;
    		:jNodeCount = 8LL ;
    } // group patch_mq_20041223_grid_mq_p3_l1
  } // group nz_linz_nzgd2000-mq20041223-grid014

group: nz_linz_nzgd2000-mq20041223-grid015 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p4_l1 {
    dimensions:
    	gridi = 70 ;
    	gridj = 68 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.125, 0., -0.125, 165.85, 0.15, 0. ;
    		:iNodeCount = 70LL ;
    		:jNodeCount = 68LL ;
    } // group patch_mq_20041223_grid_mq_p4_l1
  } // group nz_linz_nzgd2000-mq20041223-grid015

group: nz_linz_nzgd2000-mq20041223-grid016 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p5_l1 {
    dimensions:
    	gridi = 8 ;
    	gridj = 7 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -47.375, 0., -0.125, 178.45, 0.15, 0. ;
    		:iNodeCount = 8LL ;
    		:jNodeCount = 7LL ;
    } // group patch_mq_20041223_grid_mq_p5_l1
  } // group nz_linz_nzgd2000-mq20041223-grid016

group: nz_linz_nzgd2000-gs20071016-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Fiordland (George Sound) earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2007-10-16T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2008-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_gs_20071016_grid_gs_l1 {
    dimensions:
    	gridi = 37 ;
    	gridj = 27 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -43.75, 0., -0.125, 165.85, 0.15, 0. ;
    		:iNodeCount = 37LL ;
    		:jNodeCount = 27LL ;

    group: patch_gs_20071016_grid_gs_l2 {
      dimensions:
      	gridi = 45 ;
      	gridj = 37 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -44.28125, 0., -0.03125, 166.6375, 0.0375, 0. ;
      		:iNodeCount = 45LL ;
      		:jNodeCount = 37LL ;

      group: patch_gs_20071016_grid_gs_l3 {
        dimensions:
        	gridi = 54 ;
        	gridj = 52 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -44.6171875, 0., -0.0078125, 167.0875, 0.009375, 0. ;
        		:iNodeCount = 54LL ;
        		:jNodeCount = 52LL ;
        } // group patch_gs_20071016_grid_gs_l3
      } // group patch_gs_20071016_grid_gs_l2
    } // group patch_gs_20071016_grid_gs_l1
  } // group nz_linz_nzgd2000-gs20071016-grid01

group: nz_linz_nzgd2000-ds20090715-grid011 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1.05 ;
  		:timeFunctions.2.functionType = "ramp" ;
  		:timeFunctions.2.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.2.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p0_l1 {
    dimensions:
    	gridi = 11 ;
    	gridj = 11 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -50.125, 0., -0.125, 165.4, 0.15, 0. ;
    		:iNodeCount = 11LL ;
    		:jNodeCount = 11LL ;
    } // group patch_ds_20090715_grid_ds_p0_l1
  } // group nz_linz_nzgd2000-ds20090715-grid011

group: nz_linz_nzgd2000-ds20090715-grid012 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1.05 ;
  		:timeFunctions.2.functionType = "ramp" ;
  		:timeFunctions.2.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.2.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p1_l1 {
    dimensions:
    	gridi = 6 ;
    	gridj = 7 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -49.25, 0., -0.125, 178.15, 0.15, 0. ;
    		:iNodeCount = 6LL ;
    		:jNodeCount = 7LL ;
    } // group patch_ds_20090715_grid_ds_p1_l1
  } // group nz_linz_nzgd2000-ds20090715-grid012

group: nz_linz_nzgd2000-ds20090715-grid013 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1.05 ;
  		:timeFunctions.2.functionType = "ramp" ;
  		:timeFunctions.2.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.2.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p2_l1 {
    dimensions:
    	gridi = 85 ;
    	gridj = 72 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39.625, 0., -0.125, 164.65, 0.15, 0. ;
    		:iNodeCount = 85LL ;
    		:jNodeCount = 72LL ;

    group: patch_ds_20090715_grid_ds_p2_l2 {
      dimensions:
      	gridi = 67 ;
      	gridj = 73 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -44.6875, 0., -0.03125, 165.2875, 0.0375, 0. ;
      		:iNodeCount = 67LL ;
      		:jNodeCount = 73LL ;

      group: patch_ds_20090715_grid_ds_p2_l3 {
        dimensions:
        	gridi = 83 ;
        	gridj = 138 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -45.28125, 0., -0.0078125, 166.075, 0.009375, 0. ;
        		:iNodeCount = 83LL ;
        		:jNodeCount = 138LL ;
        } // group patch_ds_20090715_grid_ds_p2_l3
      } // group patch_ds_20090715_grid_ds_p2_l2
    } // group patch_ds_20090715_grid_ds_p2_l1
  } // group nz_linz_nzgd2000-ds20090715-grid013

group: nz_linz_nzgd2000-ds20090715-grid014 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1.05 ;
  		:timeFunctions.2.functionType = "ramp" ;
  		:timeFunctions.2.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.2.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.2.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p3_l1 {
    dimensions:
    	gridi = 8 ;
    	gridj = 7 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -47.375, 0., -0.125, 178.45, 0.15, 0. ;
    		:iNodeCount = 8LL ;
    		:jNodeCount = 7LL ;
    } // group patch_ds_20090715_grid_ds_p3_l1
  } // group nz_linz_nzgd2000-ds20090715-grid014

group: nz_linz_nzgd2000-c120100904-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Darfield earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2010-09-04T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c1_20100904_grid_c1_l1 {
    dimensions:
    	gridi = 55 ;
    	gridj = 52 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.375, 0., -0.125, 168.1, 0.15, 0. ;
    		:iNodeCount = 55LL ;
    		:jNodeCount = 52LL ;

    group: patch_c1_20100904_grid_c1_l2 {
      dimensions:
      	gridi = 59 ;
      	gridj = 50 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.8125, 0., -0.03125, 171.1, 0.0375, 0. ;
      		:iNodeCount = 59LL ;
      		:jNodeCount = 50LL ;

      group: patch_c1_20100904_grid_c1_l3 {
        dimensions:
        	gridi = 118 ;
        	gridj = 84 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.25, 0., -0.0078125, 171.625, 0.009375, 0. ;
        		:iNodeCount = 118LL ;
        		:jNodeCount = 84LL ;

        group: patch_c1_20100904_grid_c1_l4 {
          dimensions:
          	gridi = 306 ;
          	gridj = 141 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.423828125, 0., -0.001953125, 171.8125, 0.00234375, 0. ;
          		:iNodeCount = 306LL ;
          		:jNodeCount = 141LL ;
          } // group patch_c1_20100904_grid_c1_l4
        } // group patch_c1_20100904_grid_c1_l3
      } // group patch_c1_20100904_grid_c1_l2
    } // group patch_c1_20100904_grid_c1_l1
  } // group nz_linz_nzgd2000-c120100904-grid01

group: nz_linz_nzgd2000-c220110222-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Christchurch February earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2011-02-22T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2012-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c2_20110222_grid_c2_l1 {
    dimensions:
    	gridi = 21 ;
    	gridj = 18 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.375, 0., -0.125, 170.8, 0.15, 0. ;
    		:iNodeCount = 21LL ;
    		:jNodeCount = 18LL ;

    group: patch_c2_20110222_grid_c2_l2 {
      dimensions:
      	gridi = 38 ;
      	gridj = 34 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.03125, 0., -0.03125, 172., 0.0375, 0. ;
      		:iNodeCount = 38LL ;
      		:jNodeCount = 34LL ;

      group: patch_c2_20110222_grid_c2_l3 {
        dimensions:
        	gridi = 62 ;
        	gridj = 52 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.3515625, 0., -0.0078125, 172.4125, 0.009375, 0. ;
        		:iNodeCount = 62LL ;
        		:jNodeCount = 52LL ;

        group: patch_c2_20110222_grid_c2_l4 {
          dimensions:
          	gridi = 118 ;
          	gridj = 81 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.474609375, 0., -0.001953125, 172.56015625, 0.00234375, 0. ;
          		:iNodeCount = 118LL ;
          		:jNodeCount = 81LL ;
          } // group patch_c2_20110222_grid_c2_l4
        } // group patch_c2_20110222_grid_c2_l3
      } // group patch_c2_20110222_grid_c2_l2
    } // group patch_c2_20110222_grid_c2_l1
  } // group nz_linz_nzgd2000-c220110222-grid01

group: nz_linz_nzgd2000-c320110613-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Christchurch June earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2011-06-13T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2012-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c3_20110613_grid_c3_l1 {
    dimensions:
    	gridi = 16 ;
    	gridj = 15 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.625, 0., -0.125, 171.4, 0.15, 0. ;
    		:iNodeCount = 16LL ;
    		:jNodeCount = 15LL ;

    group: patch_c3_20110613_grid_c3_l2 {
      dimensions:
      	gridi = 33 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.09375, 0., -0.03125, 172.15, 0.0375, 0. ;
      		:iNodeCount = 33LL ;
      		:jNodeCount = 31LL ;

      group: patch_c3_20110613_grid_c3_l3 {
        dimensions:
        	gridi = 51 ;
        	gridj = 48 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.375, 0., -0.0078125, 172.515625, 0.009375, 0. ;
        		:iNodeCount = 51LL ;
        		:jNodeCount = 48LL ;

        group: patch_c3_20110613_grid_c3_l4 {
          dimensions:
          	gridi = 88 ;
          	gridj = 84 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.484375, 0., -0.001953125, 172.65390625, 0.00234375, 0. ;
          		:iNodeCount = 88LL ;
          		:jNodeCount = 84LL ;
          } // group patch_c3_20110613_grid_c3_l4
        } // group patch_c3_20110613_grid_c3_l3
      } // group patch_c3_20110613_grid_c3_l2
    } // group patch_c3_20110613_grid_c3_l1
  } // group nz_linz_nzgd2000-c320110613-grid01

group: nz_linz_nzgd2000-c420111223-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Christchurch earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2011-12-23T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2012-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c4_20111223_grid_c4_l1 {
    dimensions:
    	gridi = 15 ;
    	gridj = 13 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.75, 0., -0.125, 171.55, 0.15, 0. ;
    		:iNodeCount = 15LL ;
    		:jNodeCount = 13LL ;

    group: patch_c4_20111223_grid_c4_l2 {
      dimensions:
      	gridi = 32 ;
      	gridj = 30 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.03125, 0., -0.03125, 172.1875, 0.0375, 0. ;
      		:iNodeCount = 32LL ;
      		:jNodeCount = 30LL ;

      group: patch_c4_20111223_grid_c4_l3 {
        dimensions:
        	gridi = 52 ;
        	gridj = 44 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.3125, 0., -0.0078125, 172.553125, 0.009375, 0. ;
        		:iNodeCount = 52LL ;
        		:jNodeCount = 44LL ;

        group: patch_c4_20111223_grid_c4_l4 {
          dimensions:
          	gridi = 87 ;
          	gridj = 61 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.421875, 0., -0.001953125, 172.67734375, 0.00234375, 0. ;
          		:iNodeCount = 87LL ;
          		:jNodeCount = 61LL ;
          } // group patch_c4_20111223_grid_c4_l4
        } // group patch_c4_20111223_grid_c4_l3
      } // group patch_c4_20111223_grid_c4_l2
    } // group patch_c4_20111223_grid_c4_l1
  } // group nz_linz_nzgd2000-c420111223-grid01

group: nz_linz_nzgd2000-cs20130721-grid02 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Mw 6.6 Cook Strait earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2013-07-21T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2014-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_cs_20130721_grid_cs_20130721_l1 {
    dimensions:
    	gridi = 34 ;
    	gridj = 32 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39.5, 0., -0.125, 171.55, 0.15, 0. ;
    		:iNodeCount = 34LL ;
    		:jNodeCount = 32LL ;

    group: patch_cs_20130721_grid_cs_20130721_l2 {
      dimensions:
      	gridi = 43 ;
      	gridj = 37 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.03125, 0., -0.03125, 173.5375, 0.0375, 0. ;
      		:iNodeCount = 43LL ;
      		:jNodeCount = 37LL ;

      group: patch_cs_20130721_grid_cs_20130721_l3 {
        dimensions:
        	gridi = 73 ;
        	gridj = 57 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.3828125, 0., -0.0078125, 173.9875, 0.009375, 0. ;
        		:iNodeCount = 73LL ;
        		:jNodeCount = 57LL ;

        group: patch_cs_20130721_grid_cs_20130721_l4 {
          dimensions:
          	gridi = 90 ;
          	gridj = 68 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.537109375, 0., -0.001953125, 174.28984375, 0.00234375, 0. ;
          		:iNodeCount = 90LL ;
          		:jNodeCount = 68LL ;
          } // group patch_cs_20130721_grid_cs_20130721_l4
        } // group patch_cs_20130721_grid_cs_20130721_l3
      } // group patch_cs_20130721_grid_cs_20130721_l2
    } // group patch_cs_20130721_grid_cs_20130721_l1
  } // group nz_linz_nzgd2000-cs20130721-grid02

group: nz_linz_nzgd2000-lg20130816-grid02 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Mw 6.6 Lake Grassmere earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2013-08-16T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2014-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_lg_20130816_grid_lg_20130816_l1 {
    dimensions:
    	gridi = 39 ;
    	gridj = 39 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39.25, 0., -0.125, 170.95, 0.15, 0. ;
    		:iNodeCount = 39LL ;
    		:jNodeCount = 39LL ;

    group: patch_lg_20130816_grid_lg_20130816_l2 {
      dimensions:
      	gridi = 44 ;
      	gridj = 40 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.09375, 0., -0.03125, 173.3875, 0.0375, 0. ;
      		:iNodeCount = 44LL ;
      		:jNodeCount = 40LL ;

      group: patch_lg_20130816_grid_lg_20130816_l3 {
        dimensions:
        	gridi = 79 ;
        	gridj = 63 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.4609375, 0., -0.0078125, 173.809375, 0.009375, 0. ;
        		:iNodeCount = 79LL ;
        		:jNodeCount = 63LL ;

        group: patch_lg_20130816_grid_lg_20130816_l4 {
          dimensions:
          	gridi = 134 ;
          	gridj = 104 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.60546875, 0., -0.001953125, 174.034375, 0.00234375, 0. ;
          		:iNodeCount = 134LL ;
          		:jNodeCount = 104LL ;
          } // group patch_lg_20130816_grid_lg_20130816_l4
        } // group patch_lg_20130816_grid_lg_20130816_l3
      } // group patch_lg_20130816_grid_lg_20130816_l2
    } // group patch_lg_20130816_grid_lg_20130816_l1
  } // group nz_linz_nzgd2000-lg20130816-grid02

group: nz_linz_nzgd2000-ch20160214-grid01 {
  dimensions:
  	parameter = 3 ;

  // group attributes:
  		:comment = "Christchurch Valentines Day earthquake" ;
  		string :groupParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-02-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ch_20160214_grid_ch_20160214_l1 {
    dimensions:
    	gridi = 14 ;
    	gridj = 11 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.875, 0., -0.125, 171.7, 0.15, 0. ;
    		:iNodeCount = 14LL ;
    		:jNodeCount = 11LL ;

    group: patch_ch_20160214_grid_ch_20160214_l2 {
      dimensions:
      	gridi = 29 ;
      	gridj = 27 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.0625, 0., -0.03125, 172.225, 0.0375, 0. ;
      		:iNodeCount = 29LL ;
      		:jNodeCount = 27LL ;

      group: patch_ch_20160214_grid_ch_20160214_l3 {
        dimensions:
        	gridi = 46 ;
        	gridj = 38 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.3203125, 0., -0.0078125, 172.553125, 0.009375, 0. ;
        		:iNodeCount = 46LL ;
        		:jNodeCount = 38LL ;

        group: patch_ch_20160214_grid_ch_20160214_l4 {
          dimensions:
          	gridi = 79 ;
          	gridj = 61 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.408203125, 0., -0.001953125, 172.67265625, 0.00234375, 0. ;
          		:iNodeCount = 79LL ;
          		:jNodeCount = 61LL ;
          } // group patch_ch_20160214_grid_ch_20160214_l4
        } // group patch_ch_20160214_grid_ch_20160214_l3
      } // group patch_ch_20160214_grid_ch_20160214_l2
    } // group patch_ch_20160214_grid_ch_20160214_l1
  } // group nz_linz_nzgd2000-ch20160214-grid01

group: nz_linz_nzgd2000-ka20161114-grid01 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-11-14T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114co_h_l1_f {
    dimensions:
    	gridi = 89 ;
    	gridj = 110 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -34., 0., -0.125, 165.85, 0.15, 0. ;
    		:iNodeCount = 89LL ;
    		:jNodeCount = 110LL ;

    group: patch_ka_20161114_grid_ka_20161114co_h_l2_f {
      dimensions:
      	gridi = 95 ;
      	gridj = 82 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -40.8125, 0., -0.03125, 171.925, 0.0375, 0. ;
      		:iNodeCount = 95LL ;
      		:jNodeCount = 82LL ;
      } // group patch_ka_20161114_grid_ka_20161114co_h_l2_f
    } // group patch_ka_20161114_grid_ka_20161114co_h_l1_f
  } // group nz_linz_nzgd2000-ka20161114-grid01

group: nz_linz_nzgd2000-ka20161114-grid02 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114co_h_l2_r {
    dimensions:
    	gridi = 65 ;
    	gridj = 53 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -41.28125, 0., -0.03125, 172.525, 0.0375, 0. ;
    		:iNodeCount = 65LL ;
    		:jNodeCount = 53LL ;

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_00 {
      dimensions:
      	gridi = 115 ;
      	gridj = 94 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.1484375, 0., -0.0078125, 172.571875, 0.009375, 0. ;
      		:iNodeCount = 115LL ;
      		:jNodeCount = 94LL ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_00 {
        dimensions:
        	gridi = 106 ;
        	gridj = 107 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 172.7828125, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 107LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_00

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_01 {
        dimensions:
        	gridi = 11 ;
        	gridj = 26 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.435546875, 0., -0.001953125, 173.00546875, 0.00234375, 0. ;
        		:iNodeCount = 11LL ;
        		:jNodeCount = 26LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_01

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_02 {
        dimensions:
        	gridi = 106 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.02890625, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_02

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_03 {
        dimensions:
        	gridi = 106 ;
        	gridj = 51 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.38671875, 0., -0.001953125, 173.02890625, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 51LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_03

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_04 {
        dimensions:
        	gridi = 106 ;
        	gridj = 88 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.275, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 88LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_04

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_05 {
        dimensions:
        	gridi = 106 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.275, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_05

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_060 {
        dimensions:
        	gridi = 21 ;
        	gridj = 63 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.47421875, 0.00234375, 0. ;
        		:iNodeCount = 21LL ;
        		:jNodeCount = 63LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_060

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_080 {
        dimensions:
        	gridi = 52 ;
        	gridj = 30 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        		:iNodeCount = 52LL ;
        		:jNodeCount = 30LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_080

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_090 {
        dimensions:
        	gridi = 52 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        		:iNodeCount = 52LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_090

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_100 {
        dimensions:
        	gridi = 52 ;
        	gridj = 63 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        		:iNodeCount = 52LL ;
        		:jNodeCount = 63LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_100
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_00

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_01 {
      dimensions:
      	gridi = 53 ;
      	gridj = 89 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.4609375, 0., -0.0078125, 173.153125, 0.009375, 0. ;
      		:iNodeCount = 53LL ;
      		:jNodeCount = 89LL ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_061 {
        dimensions:
        	gridi = 21 ;
        	gridj = 49 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.47421875, 0.00234375, 0. ;
        		:iNodeCount = 21LL ;
        		:jNodeCount = 49LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_061

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_07 {
        dimensions:
        	gridi = 9 ;
        	gridj = 6 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.044921875, 0., -0.001953125, 173.50234375, 0.0023437500000014, 0. ;
        		:iNodeCount = 9LL ;
        		:jNodeCount = 6LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_07

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_101 {
        dimensions:
        	gridi = 52 ;
        	gridj = 49 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        		:iNodeCount = 52LL ;
        		:jNodeCount = 49LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_101

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_110 {
        dimensions:
        	gridi = 52 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        		:iNodeCount = 52LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_110
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_01

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_02 {
      dimensions:
      	gridi = 73 ;
      	gridj = 63 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.1484375, 0., -0.0078125, 173.640625, 0.009375, 0. ;
      		:iNodeCount = 73LL ;
      		:jNodeCount = 63LL ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_081 {
        dimensions:
        	gridi = 28 ;
        	gridj = 30 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        		:iNodeCount = 28LL ;
        		:jNodeCount = 30LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_081

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_091 {
        dimensions:
        	gridi = 55 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        		:iNodeCount = 55LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_091

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_102 {
        dimensions:
        	gridi = 55 ;
        	gridj = 63 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        		:iNodeCount = 55LL ;
        		:jNodeCount = 63LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_102

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_13 {
        dimensions:
        	gridi = 87 ;
        	gridj = 95 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        		:iNodeCount = 87LL ;
        		:jNodeCount = 95LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_13

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_140 {
        dimensions:
        	gridi = 106 ;
        	gridj = 63 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 63LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_140

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_170 {
        dimensions:
        	gridi = 62 ;
        	gridj = 41 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        		:iNodeCount = 62LL ;
        		:jNodeCount = 41LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_170
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_02

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_03 {
      dimensions:
      	gridi = 114 ;
      	gridj = 94 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.421875, 0., -0.0078125, 173.640625, 0.009375, 0. ;
      		:iNodeCount = 114LL ;
      		:jNodeCount = 94LL ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_103 {
        dimensions:
        	gridi = 55 ;
        	gridj = 49 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        		:iNodeCount = 55LL ;
        		:jNodeCount = 49LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_103

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_111 {
        dimensions:
        	gridi = 55 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        		:iNodeCount = 55LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_111

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_12 {
        dimensions:
        	gridi = 15 ;
        	gridj = 10 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.822265625, 0., -0.001953125, 173.734375, 0.00234375, 0. ;
        		:iNodeCount = 15LL ;
        		:jNodeCount = 10LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_12

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_141 {
        dimensions:
        	gridi = 106 ;
        	gridj = 49 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 49LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_141

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_15 {
        dimensions:
        	gridi = 106 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_15

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_16 {
        dimensions:
        	gridi = 106 ;
        	gridj = 41 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.76171875, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 41LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_16

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_171 {
        dimensions:
        	gridi = 62 ;
        	gridj = 49 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        		:iNodeCount = 62LL ;
        		:jNodeCount = 49LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_171

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_18 {
        dimensions:
        	gridi = 106 ;
        	gridj = 111 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 111LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_18

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_19 {
        dimensions:
        	gridi = 106 ;
        	gridj = 93 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.66015625, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        		:iNodeCount = 106LL ;
        		:jNodeCount = 93LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_19

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_20 {
        dimensions:
        	gridi = 59 ;
        	gridj = 35 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 174.259375, 0.00234375, 0. ;
        		:iNodeCount = 59LL ;
        		:jNodeCount = 35LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_20

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_21 {
        dimensions:
        	gridi = 104 ;
        	gridj = 110 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.626953125, 0., -0.001953125, 174.259375, 0.00234375, 0. ;
        		:iNodeCount = 104LL ;
        		:jNodeCount = 110LL ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_21
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_03
    } // group patch_ka_20161114_grid_ka_20161114co_h_l2_r
  } // group nz_linz_nzgd2000-ka20161114-grid02

group: nz_linz_nzgd2000-ka20161114-grid03 {
  dimensions:
  	parameter = 1 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		:groupParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114co_v_l1 {
    dimensions:
    	gridi = 86 ;
    	gridj = 108 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -34.25, 0., -0.125, 166.3, 0.15, 0. ;
    		:iNodeCount = 86LL ;
    		:jNodeCount = 108LL ;

    group: patch_ka_20161114_grid_ka_20161114co_v_l2 {
      dimensions:
      	gridi = 74 ;
      	gridj = 67 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.0625, 0., -0.03125, 172.225, 0.0375, 0. ;
      		:iNodeCount = 74LL ;
      		:jNodeCount = 67LL ;

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_00 {
        dimensions:
        	gridi = 103 ;
        	gridj = 89 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1171875, 0., -0.0078125, 172.65625, 0.009375, 0. ;
        		:iNodeCount = 103LL ;
        		:jNodeCount = 89LL ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_00 {
          dimensions:
          	gridi = 103 ;
          	gridj = 88 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.490234375, 0., -0.001953125, 172.79921875, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 88LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_00

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_01 {
          dimensions:
          	gridi = 103 ;
          	gridj = 105 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.03828125, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 105LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_01

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_02 {
          dimensions:
          	gridi = 89 ;
          	gridj = 52 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.353515625, 0., -0.001953125, 173.07109375, 0.00234375, 0. ;
          		:iNodeCount = 89LL ;
          		:jNodeCount = 52LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_02

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_03 {
          dimensions:
          	gridi = 103 ;
          	gridj = 100 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.27734375, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 100LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_03

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_04 {
          dimensions:
          	gridi = 103 ;
          	gridj = 89 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.28125, 0., -0.001953125, 173.27734375, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 89LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_04

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_050 {
          dimensions:
          	gridi = 21 ;
          	gridj = 67 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.46953125, 0.00234375, 0. ;
          		:iNodeCount = 21LL ;
          		:jNodeCount = 67LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_050

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_060 {
          dimensions:
          	gridi = 42 ;
          	gridj = 34 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          		:iNodeCount = 42LL ;
          		:jNodeCount = 34LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_060

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_070 {
          dimensions:
          	gridi = 42 ;
          	gridj = 107 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.24609375, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          		:iNodeCount = 42LL ;
          		:jNodeCount = 107LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_070

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_080 {
          dimensions:
          	gridi = 42 ;
          	gridj = 67 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          		:iNodeCount = 42LL ;
          		:jNodeCount = 67LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_080
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_00

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_01 {
        dimensions:
        	gridi = 44 ;
        	gridj = 70 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.578125, 0., -0.0078125, 173.209375, 0.009375, 0. ;
        		:iNodeCount = 44LL ;
        		:jNodeCount = 70LL ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_051 {
          dimensions:
          	gridi = 21 ;
          	gridj = 33 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.46953125, 0.00234375, 0. ;
          		:iNodeCount = 21LL ;
          		:jNodeCount = 33LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_051

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_081 {
          dimensions:
          	gridi = 42 ;
          	gridj = 41 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          		:iNodeCount = 42LL ;
          		:jNodeCount = 41LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_081

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_090 {
          dimensions:
          	gridi = 12 ;
          	gridj = 66 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.912109375, 0., -0.001953125, 173.58671875, 0.00234375, 0. ;
          		:iNodeCount = 12LL ;
          		:jNodeCount = 66LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_090
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_01

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_02 {
        dimensions:
        	gridi = 79 ;
        	gridj = 60 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1171875, 0., -0.0078125, 173.6125, 0.009375, 0. ;
        		:iNodeCount = 79LL ;
        		:jNodeCount = 60LL ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_061 {
          dimensions:
          	gridi = 62 ;
          	gridj = 34 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          		:iNodeCount = 62LL ;
          		:jNodeCount = 34LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_061

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_071 {
          dimensions:
          	gridi = 62 ;
          	gridj = 107 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.24609375, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          		:iNodeCount = 62LL ;
          		:jNodeCount = 107LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_071

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_082 {
          dimensions:
          	gridi = 62 ;
          	gridj = 67 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          		:iNodeCount = 62LL ;
          		:jNodeCount = 67LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_082

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_10 {
          dimensions:
          	gridi = 7 ;
          	gridj = 4 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          		:iNodeCount = 7LL ;
          		:jNodeCount = 4LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_10

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_11 {
          dimensions:
          	gridi = 93 ;
          	gridj = 107 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.24609375, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          		:iNodeCount = 93LL ;
          		:jNodeCount = 107LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_11

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_120 {
          dimensions:
          	gridi = 103 ;
          	gridj = 67 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 67LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_120

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_140 {
          dimensions:
          	gridi = 40 ;
          	gridj = 59 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.99453125, 0.00234375, 0. ;
          		:iNodeCount = 40LL ;
          		:jNodeCount = 59LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_140
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_02

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_03 {
        dimensions:
        	gridi = 103 ;
        	gridj = 88 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.4375, 0., -0.0078125, 173.6125, 0.009375, 0. ;
        		:iNodeCount = 103LL ;
        		:jNodeCount = 88LL ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_083 {
          dimensions:
          	gridi = 62 ;
          	gridj = 41 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          		:iNodeCount = 62LL ;
          		:jNodeCount = 41LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_083

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_091 {
          dimensions:
          	gridi = 62 ;
          	gridj = 66 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.912109375, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          		:iNodeCount = 62LL ;
          		:jNodeCount = 66LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_091

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_121 {
          dimensions:
          	gridi = 103 ;
          	gridj = 41 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 41LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_121

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_13 {
          dimensions:
          	gridi = 103 ;
          	gridj = 93 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.859375, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 93LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_13

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_141 {
          dimensions:
          	gridi = 40 ;
          	gridj = 41 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.99453125, 0.00234375, 0. ;
          		:iNodeCount = 40LL ;
          		:jNodeCount = 41LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_141

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_15 {
          dimensions:
          	gridi = 103 ;
          	gridj = 107 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.83203125, 0., -0.001953125, 173.99453125, 0.00234375, 0. ;
          		:iNodeCount = 103LL ;
          		:jNodeCount = 107LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_15

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_16 {
          dimensions:
          	gridi = 64 ;
          	gridj = 78 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.681640625, 0., -0.001953125, 174.0859375, 0.00234375, 0. ;
          		:iNodeCount = 64LL ;
          		:jNodeCount = 78LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_16

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_17 {
          dimensions:
          	gridi = 56 ;
          	gridj = 45 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.83203125, 0., -0.001953125, 174.23359375, 0.00234375, 0. ;
          		:iNodeCount = 56LL ;
          		:jNodeCount = 45LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_17

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_18 {
          dimensions:
          	gridi = 101 ;
          	gridj = 106 ;
          variables:
          	float data(gridj, gridi, parameter) ;
          		data:_Storage = "contiguous" ;
          		data:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.626953125, 0., -0.001953125, 174.23359375, 0.00234375, 0. ;
          		:iNodeCount = 101LL ;
          		:jNodeCount = 106LL ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_18
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_03
      } // group patch_ka_20161114_grid_ka_20161114co_v_l2
    } // group patch_ka_20161114_grid_ka_20161114co_v_l1
  } // group nz_linz_nzgd2000-ka20161114-grid03

group: nz_linz_nzgd2000-ka20161114-grid04 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake postearthquake month 0-1,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe1_h_l1_f {
    dimensions:
    	gridi = 46 ;
    	gridj = 39 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39., 0., -0.125, 169.6, 0.15, 0. ;
    		:iNodeCount = 46LL ;
    		:jNodeCount = 39LL ;

    group: patch_ka_20161114_grid_ka_20161114pe1_h_l2_f {
      dimensions:
      	gridi = 74 ;
      	gridj = 59 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.125, 0., -0.03125, 172.6375, 0.0375, 0. ;
      		:iNodeCount = 74LL ;
      		:jNodeCount = 59LL ;
      } // group patch_ka_20161114_grid_ka_20161114pe1_h_l2_f
    } // group patch_ka_20161114_grid_ka_20161114pe1_h_l1_f
  } // group nz_linz_nzgd2000-ka20161114-grid04

group: nz_linz_nzgd2000-ka20161114-grid05 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake postearthquake month 0-1,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe1_h_l2_r {
    dimensions:
    	gridi = 67 ;
    	gridj = 56 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -41.28125, 0., -0.03125, 172.45, 0.0375, 0. ;
    		:iNodeCount = 67LL ;
    		:jNodeCount = 56LL ;

    group: patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_00 {
      dimensions:
      	gridi = 93 ;
      	gridj = 83 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.0546875, 0., -0.0078125, 172.834375, 0.009375, 0. ;
      		:iNodeCount = 93LL ;
      		:jNodeCount = 83LL ;
      } // group patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_00

    group: patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_01 {
      dimensions:
      	gridi = 92 ;
      	gridj = 125 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.5703125, 0., -0.0078125, 173.696875, 0.009375, 0. ;
      		:iNodeCount = 92LL ;
      		:jNodeCount = 125LL ;
      } // group patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_01
    } // group patch_ka_20161114_grid_ka_20161114pe1_h_l2_r
  } // group nz_linz_nzgd2000-ka20161114-grid05

group: nz_linz_nzgd2000-ka20161114-grid06 {
  dimensions:
  	parameter = 1 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake postearthquake month 0-1,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		:groupParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe1_v_l1 {
    dimensions:
    	gridi = 29 ;
    	gridj = 27 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.5, 0., -0.125, 171.85, 0.15, 0. ;
    		:iNodeCount = 29LL ;
    		:jNodeCount = 27LL ;

    group: patch_ka_20161114_grid_ka_20161114pe1_v_l2 {
      dimensions:
      	gridi = 72 ;
      	gridj = 74 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -40.75, 0., -0.03125, 172.675, 0.0375, 0. ;
      		:iNodeCount = 72LL ;
      		:jNodeCount = 74LL ;

      group: patch_ka_20161114_grid_ka_20161114pe1_v_l3_00 {
        dimensions:
        	gridi = 92 ;
        	gridj = 82 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.0078125, 172.84375, 0.009375, 0. ;
        		:iNodeCount = 92LL ;
        		:jNodeCount = 82LL ;
        } // group patch_ka_20161114_grid_ka_20161114pe1_v_l3_00

      group: patch_ka_20161114_grid_ka_20161114pe1_v_l3_01 {
        dimensions:
        	gridi = 91 ;
        	gridj = 119 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.609375, 0., -0.0078125, 173.696875, 0.009375, 0. ;
        		:iNodeCount = 91LL ;
        		:jNodeCount = 119LL ;
        } // group patch_ka_20161114_grid_ka_20161114pe1_v_l3_01
      } // group patch_ka_20161114_grid_ka_20161114pe1_v_l2
    } // group patch_ka_20161114_grid_ka_20161114pe1_v_l1
  } // group nz_linz_nzgd2000-ka20161114-grid06

group: nz_linz_nzgd2000-ka20161114-grid10 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\nRefinement for horizontal difference between observations and model\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-11-14T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_hor_refinement {
    dimensions:
    	gridi = 43 ;
    	gridj = 40 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -38.625, 0., -0.125, 171.1, 0.15, 0. ;
    		:iNodeCount = 43LL ;
    		:jNodeCount = 40LL ;
    } // group patch_ka_20161114_grid_hor_refinement
  } // group nz_linz_nzgd2000-ka20161114-grid10

group: nz_linz_nzgd2000-ka20161114-grid11 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Kaikoura earthquake second refinement grid - horizontal" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_hor_refinement2 {
    dimensions:
    	gridi = 214 ;
    	gridj = 192 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.56, 0., -0.015, 171.5, 0.02, 0. ;
    		:iNodeCount = 214LL ;
    		:jNodeCount = 192LL ;
    } // group patch_ka_20161114_grid_hor_refinement2
  } // group nz_linz_nzgd2000-ka20161114-grid11

group: nz_linz_nzgd2000-ka20161114-grid12 {
  dimensions:
  	parameter = 1 ;

  // group attributes:
  		:comment = "Kaikoura earthquake second refinement grid -vertical" ;
  		:groupParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "step" ;
  		:timeFunctions.1.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_vrt_refinement2 {
    dimensions:
    	gridi = 216 ;
    	gridj = 199 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.395, 0., -0.015, 171.9, 0.02, 0. ;
    		:iNodeCount = 216LL ;
    		:jNodeCount = 199LL ;
    } // group patch_ka_20161114_grid_vrt_refinement2
  } // group nz_linz_nzgd2000-ka20161114-grid12

group: nz_linz_nzgd2000-ka20161114-grid07 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake months1-3 post-earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe3_h_l1_f {
    dimensions:
    	gridi = 46 ;
    	gridj = 40 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -38.875, 0., -0.125, 169.6, 0.15, 0. ;
    		:iNodeCount = 46LL ;
    		:jNodeCount = 40LL ;

    group: patch_ka_20161114_grid_ka_20161114pe3_h_l2_f {
      dimensions:
      	gridi = 66 ;
      	gridj = 60 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.0625, 0., -0.03125, 172.525, 0.0375, 0. ;
      		:iNodeCount = 66LL ;
      		:jNodeCount = 60LL ;
      } // group patch_ka_20161114_grid_ka_20161114pe3_h_l2_f
    } // group patch_ka_20161114_grid_ka_20161114pe3_h_l1_f
  } // group nz_linz_nzgd2000-ka20161114-grid07

group: nz_linz_nzgd2000-ka20161114-grid08 {
  dimensions:
  	parameter = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake months1-3 post-earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :groupParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe3_h_l2_r {
    dimensions:
    	gridi = 67 ;
    	gridj = 56 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -41.28125, 0., -0.03125, 172.45, 0.0375, 0. ;
    		:iNodeCount = 67LL ;
    		:jNodeCount = 56LL ;

    group: patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_00 {
      dimensions:
      	gridi = 88 ;
      	gridj = 91 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42., 0., -0.0078125, 172.91875, 0.009375, 0. ;
      		:iNodeCount = 88LL ;
      		:jNodeCount = 91LL ;
      } // group patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_00

    group: patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_01 {
      dimensions:
      	gridi = 88 ;
      	gridj = 122 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.5546875, 0., -0.0078125, 173.734375, 0.009375, 0. ;
      		:iNodeCount = 88LL ;
      		:jNodeCount = 122LL ;
      } // group patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_01
    } // group patch_ka_20161114_grid_ka_20161114pe3_h_l2_r
  } // group nz_linz_nzgd2000-ka20161114-grid08

group: nz_linz_nzgd2000-ka20161114-grid09 {
  dimensions:
  	parameter = 1 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake months1-3 post-earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		:groupParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe3_v_l1 {
    dimensions:
    	gridi = 31 ;
    	gridj = 28 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.25, 0., -0.125, 171.4, 0.15, 0. ;
    		:iNodeCount = 31LL ;
    		:jNodeCount = 28LL ;

    group: patch_ka_20161114_grid_ka_20161114pe3_v_l2 {
      dimensions:
      	gridi = 82 ;
      	gridj = 76 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -40.65625, 0., -0.03125, 172.1875, 0.0375, 0. ;
      		:iNodeCount = 82LL ;
      		:jNodeCount = 76LL ;

      group: patch_ka_20161114_grid_ka_20161114pe3_v_l3_00 {
        dimensions:
        	gridi = 92 ;
        	gridj = 80 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0703125, 0., -0.0078125, 172.825, 0.009375, 0. ;
        		:iNodeCount = 92LL ;
        		:jNodeCount = 80LL ;
        } // group patch_ka_20161114_grid_ka_20161114pe3_v_l3_00

      group: patch_ka_20161114_grid_ka_20161114pe3_v_l3_01 {
        dimensions:
        	gridi = 92 ;
        	gridj = 121 ;
        variables:
        	float data(gridj, gridi, parameter) ;
        		data:_Storage = "contiguous" ;
        		data:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.5859375, 0., -0.0078125, 173.678125, 0.009375, 0. ;
        		:iNodeCount = 92LL ;
        		:jNodeCount = 121LL ;
        } // group patch_ka_20161114_grid_ka_20161114pe3_v_l3_01
      } // group patch_ka_20161114_grid_ka_20161114pe3_v_l2
    } // group patch_ka_20161114_grid_ka_20161114pe3_v_l1
  } // group nz_linz_nzgd2000-ka20161114-grid09
}

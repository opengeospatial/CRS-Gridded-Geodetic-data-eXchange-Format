netcdf test_geoid {

// global attributes:
		:ggxfVersion = "1.0" ;
		:filename = "g2018vi.gxt" ;
		:content = "heightCorrectionModel" ;
		:remark = "hybrid geoid" ;
		:contentApplicability.boundingBox.southBoundLatitude = 17.67 ;
		:contentApplicability.boundingBox.westBoundLongitude = -65.09 ;
		:contentApplicability.boundingBox.northBoundLatitude = 18.42 ;
		:contentApplicability.boundingBox.eastBoundLongitude = -64.6 ;
		:contentApplicability.description = "US Virgin Islands - onshore." ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,3],\n  AXIS[\"Geodetic latitude (Lat)\",north,\n    ANGLEUNIT[\"degree\\\",0.0174532925199433]],\n  AXIS[\"Geodetic longitude (Lon)\",east,\n    ANGLEUNIT[\"degree\\\",0.0174532925199433]],\n  AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1]]]\n" ;
		:targetCrsWkt = "VERTCRS[\"VIVD09 - NOHt\",\n  VDATUM[\"Virgin Islands Vertical Datum of 2009\"],\n  CS[vertical,1],\n  AXIS[\"Gravity-related height (H)\",up],\n  LENGTHUNIT[\"metre\",1]]\n" ;
		:operationAccuracy = 0.015 ;
		:organisationName = "National Geodetic Survey, National Oceanic and Atmospheric Administration." ;
		:deliveryPoint = "1315 East West Hwy" ;
		:city = "Silver Spring" ;
		:postalCode = "20910" ;
		:country = "United States of America" ;
		:onlineResourceLinkage = "https://geodesy.noaa.gov/PC_PROD/GEOID18/Format_ascii/g2018p0.asc.zip" ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: Puerto\ Rico\ Virgin\ Islands\ GEOID18 {
  dimensions:
  	nParam = 1 ;

  // group attributes:
  		:remark = "" ;
  		:parameters.count = 1LL ;
  		:parameters.0.parameterName = "geoidHeight" ;
  		:parameters.0.lengthUnit = "metre" ;
  		:parameters.0.unitSiRatio = 1. ;
  		:interpolationMethod = "biquadratic" ;

  group: Puerto\ Rico\ Virgin\ Islands\ GEOID18 {
    dimensions:
    	nCol = 3 ;
    	nRow = 4 ;
    variables:
    	double data(nRow, nCol, nParam) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 15., 0., 1.66667, -69., 1.5, 0. ;
    		:iNodeMaximum = 2LL ;
    		:jNodeMaximum = 3LL ;
    data:

     data =
  -29.2936,
  -29.3314,
  -29.371,
  -29.4121,
  -29.454,
  -29.4965,
  -29.5382,
  -29.5807,
  -29.6233,
  -29.666,
  -29.709,
  -29.7522 ;
    } // group Puerto\ Rico\ Virgin\ Islands\ GEOID18
  } // group Puerto\ Rico\ Virgin\ Islands\ GEOID18
}

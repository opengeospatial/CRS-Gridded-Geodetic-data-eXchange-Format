netcdf alaska_velocity {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:content = "velocityGrid" ;
		:source_file = "alaska_velocity.ggxf" ;
		:title = "Alaska velocity grid" ;
		:summary = "Alaska velocity model" ;
		:product_version = "Test_1.0" ;
		:date_issued = "2022-09" ;
		:institution = "Test developer" ;
		:geospatial_lat_min = 53.25 ;
		:geospatial_lon_min = -170. ;
		:geospatial_lat_max = 73. ;
		:geospatial_lon_max = -130. ;
		:extent_description = "Alaska" ;
		:interpolationCrsWkt = "GEOGCRS[\"ITRF2008\",DYNAMIC[FRAMEEPOCH[2005]],DATUM[\"International Terrestrial Reference Frame 2008\",ELLIPSOID[\"GRS 1980\",6378137,298.257222101,LENGTHUNIT[\"metre\",1]]],PRIMEM[\"Greenwich\",0,ANGLEUNIT[\"degree\",0.0174532925199433]],CS[ellipsoidal,3],AXIS[\"geodetic latitude (Lat)\",north,ORDER[1],ANGLEUNIT[\"degree\",0.0174532925199433]],AXIS[\"geodetic longitude (Lon)\",east,ORDER[2],ANGLEUNIT[\"degree\",0.0174532925199433]],AXIS[\"ellipsoidal height (h)\",up,ORDER[3],LENGTHUNIT[\"metre\",1]],USAGE[SCOPE[\"Geodesy.\"],AREA[\"World.\"],BBOX[-90,-180,90,180]],ID[\"EPSG\",7911]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"ITRF2008\",DYNAMIC[FRAMEEPOCH[2005]],DATUM[\"International Terrestrial Reference Frame 2008\",ELLIPSOID[\"GRS 1980\",6378137,298.257222101,LENGTHUNIT[\"metre\",1]]],PRIMEM[\"Greenwich\",0,ANGLEUNIT[\"degree\",0.0174532925199433]],CS[ellipsoidal,3],AXIS[\"geodetic latitude (Lat)\",north,ORDER[1],ANGLEUNIT[\"degree\",0.0174532925199433]],AXIS[\"geodetic longitude (Lon)\",east,ORDER[2],ANGLEUNIT[\"degree\",0.0174532925199433]],AXIS[\"ellipsoidal height (h)\",up,ORDER[3],LENGTHUNIT[\"metre\",1]],USAGE[SCOPE[\"Geodesy.\"],AREA[\"World.\"],BBOX[-90,-180,90,180]],ID[\"EPSG\",7911]]\n" ;
		:targetCrsWkt = "GEOGCRS[\"ITRF2008\",DYNAMIC[FRAMEEPOCH[2005]],DATUM[\"International Terrestrial Reference Frame 2008\",ELLIPSOID[\"GRS 1980\",6378137,298.257222101,LENGTHUNIT[\"metre\",1]]],PRIMEM[\"Greenwich\",0,ANGLEUNIT[\"degree\",0.0174532925199433]],CS[ellipsoidal,3],AXIS[\"geodetic latitude (Lat)\",north,ORDER[1],ANGLEUNIT[\"degree\",0.0174532925199433]],AXIS[\"geodetic longitude (Lon)\",east,ORDER[2],ANGLEUNIT[\"degree\",0.0174532925199433]],AXIS[\"ellipsoidal height (h)\",up,ORDER[3],LENGTHUNIT[\"metre\",1]],USAGE[SCOPE[\"Geodesy.\"],AREA[\"World.\"],BBOX[-90,-180,90,180]],ID[\"EPSG\",7911]]\n" ;
		:parameters.count = 3LL ;
		:parameters.0.parameterName = "velocityEast" ;
		:parameters.0.parameterSet = "velocity" ;
		:parameters.0.sourceCrsAxis = 1LL ;
		:parameters.0.unitName = "m/yr" ;
		:parameters.0.unitSiRatio = 3.16887651727315e-08 ;
		:parameters.1.parameterName = "velocityNorth" ;
		:parameters.1.parameterSet = "velocity" ;
		:parameters.1.sourceCrsAxis = 0LL ;
		:parameters.1.unitName = "m/yr" ;
		:parameters.1.unitSiRatio = 3.16887651727315e-08 ;
		:parameters.2.parameterName = "velocityUp" ;
		:parameters.2.parameterSet = "velocity" ;
		:parameters.2.sourceCrsAxis = 2LL ;
		:parameters.2.unitName = "m/yr" ;
		:parameters.2.unitSiRatio = 3.16887651727315e-08 ;
		:operationAccuracy = 0.001 ;
		:_NCProperties = "version=2,netcdf=4.9.0,hdf5=1.12.2" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: alaska-grids {
  dimensions:
  	velocityCount = 3 ;

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: Alaska-mainland {
    dimensions:
    	iNodeCount = 69 ;
    	jNodeCount = 161 ;
    variables:
    	float velocity(iNodeCount, jNodeCount, velocityCount) ;
    		velocity:_Storage = "contiguous" ;
    		velocity:_Endianness = "little" ;

    // group attributes:
    		:gridPriority = 1LL ;
    		:affineCoeffs = 56., 0.25, 0., -170., 0., 0.25 ;
    } // group Alaska-mainland

  group: Alaska-south-central {
    dimensions:
    	iNodeCount = 51 ;
    	jNodeCount = 76 ;
    variables:
    	float velocity(iNodeCount, jNodeCount, velocityCount) ;
    		velocity:_Storage = "contiguous" ;
    		velocity:_Endianness = "little" ;

    // group attributes:
    		:gridPriority = 2LL ;
    		:affineCoeffs = 53.25, 0.25, 0., -162., 0., 0.25 ;
    } // group Alaska-south-central

  group: Alaska-south-east {
    dimensions:
    	iNodeCount = 41 ;
    	jNodeCount = 49 ;
    variables:
    	float velocity(iNodeCount, jNodeCount, velocityCount) ;
    		velocity:_Storage = "contiguous" ;
    		velocity:_Endianness = "little" ;

    // group attributes:
    		:gridPriority = 3LL ;
    		:affineCoeffs = 54., 0.25, 0., -142., 0., 0.25 ;
    } // group Alaska-south-east

  group: Alaska-st-elias {
    dimensions:
    	iNodeCount = 27 ;
    	jNodeCount = 41 ;
    variables:
    	float velocity(iNodeCount, jNodeCount, velocityCount) ;
    		velocity:_Storage = "contiguous" ;
    		velocity:_Endianness = "little" ;

    // group attributes:
    		:gridPriority = 4LL ;
    		:affineCoeffs = 56.5, 0.25, 0., -150., 0., 0.25 ;
    } // group Alaska-st-elias
  } // group alaska-grids
}

netcdf test_geoid {

// global attributes:
		:ggxfVersion = "GGXF-1.0" ;
		:filename = "tiny_geoid.gxt" ;
		:content = "geoidModel" ;
		:title = "hybrid geoid" ;
		:abstract = "Tiny geoid for testing GGXF implementation" ;
		:contentApplicabilityExtent.boundingBox.southBoundLatitude = 22.5 ;
		:contentApplicabilityExtent.boundingBox.westBoundLongitude = -69. ;
		:contentApplicabilityExtent.boundingBox.northBoundLatitude = 24.6 ;
		:contentApplicabilityExtent.boundingBox.eastBoundLongitude = -67. ;
		:contentApplicabilityExtent.extentDescription = "Tiny example geoid." ;
		:interpolationCrsWkt = "GEOGCS[\"WGS 84\",\n  DATUM[\"WGS_1984\",\n    SPHEROID[\"WGS 84\",6378137,298.257223563,AUTHORITY[\"EPSG\",\"7030\"]],\n    AUTHORITY[\"EPSG\",\"6326\"]],\n  PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],\n  UNIT[\"degree\",0.01745329251994328,AUTHORITY[\"EPSG\",\"9122\"]],\n  AUTHORITY[\"EPSG\",\"4326\"]]\n" ;
		:sourceCrsWkt = "GEOGCS[\"WGS 84\",\n  DATUM[\"WGS_1984\",\n    SPHEROID[\"WGS 84\",6378137,298.257223563,AUTHORITY[\"EPSG\",\"7030\"]],\n    AUTHORITY[\"EPSG\",\"6326\"]],\n  PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],\n  UNIT[\"degree\",0.01745329251994328,AUTHORITY[\"EPSG\",\"9122\"]],\n  AUTHORITY[\"EPSG\",\"4326\"]]\n" ;
		:targetCrsWkt = "VERTCRS[\"VRTDTM2000\",\n  VDATUM[\"A vertical datum\"],\n  CS[vertical,1],\n  AXIS[\"Gravity-related height (H)\",up],\n  LENGTHUNIT[\"metre\",1]]\n" ;
		:parameters.count = 1LL ;
		:parameters.0.parameterName = "geoidHeight" ;
		:parameters.0.lengthUnit = "metre" ;
		:parameters.0.unitSiRatio = 1. ;
		:operationAccuracy = 0.015 ;
		:organisationName = "A Hypothetical National Geodetic Survey." ;
		:deliveryPoint = "Somewhere" ;
		:city = "A city" ;
		:postalCode = "99999" ;
		:country = "United States of America" ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: default {
  dimensions:
  	parameter = 1 ;

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: geoid_grid {
    dimensions:
    	gridi = 3 ;
    	gridj = 4 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:iNodeCount = 3LL ;
    		:jNodeCount = 4LL ;
    		:affineCoeffs = 22.5, 0., 0.7, -69., 1., 0. ;
    data:

     data =
  -10.5,
  -20.5,
  -30.5,
  -11.5,
  -21.5,
  -31.5,
  -12.5,
  -22.5,
  -32.5,
  -13.5,
  -23.5,
  -33.5 ;
    } // group geoid_grid
  } // group default
}

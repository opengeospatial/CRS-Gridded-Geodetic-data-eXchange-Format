netcdf ca_ntv2 {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "ca_ntv2.ggxf" ;
		:title = "Canadian National NAD27-NAD83(Original) NTV2 transformation" ;
		:summary = "Canadian National NAD27-NAD83(Original) NTV2 transformation" ;
		:content = "geographic2dOffsets" ;
		:product_version = "National Transformation v2_0" ;
		:date_issued = "1995-02" ;
		:institution = "Geodetic Survey Division, Natural Resources Canada" ;
		:publisher_url = "https://webapp.geod.nrcan.gc.ca/geod/data-donnees/transformations.php" ;
		:license = "https://open.canada.ca/en/open-government-licence-canada" ;
		:geospatial_lat_min = 40. ;
		:geospatial_lon_min = -141. ;
		:geospatial_lat_max = 84. ;
		:geospatial_lon_max = -44. ;
		:extent_description = "Canada south of 84°N" ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:targetCrsWkt = "GEOGCRS[\"NAD83(Original)\",\n  DATUM[\"North American Datum 1983\",\n    ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:parameters.count = 4LL ;
		:parameters.0.parameterName = "latitudeOffset" ;
		:parameters.0.parameterSet = "offset" ;
		:parameters.0.sourceCrsAxis = 0LL ;
		:parameters.0.unitName = "arc-second" ;
		:parameters.0.unitSiRatio = 4.84813681109536e-06 ;
		:parameters.1.parameterName = "longitudeOffset" ;
		:parameters.1.parameterSet = "offset" ;
		:parameters.1.sourceCrsAxis = 1LL ;
		:parameters.1.unitName = "arc-second" ;
		:parameters.1.unitSiRatio = 4.84813681109536e-06 ;
		:parameters.2.parameterName = "latitudeOffsetUncertainty" ;
		:parameters.2.parameterSet = "offsetUncertainty" ;
		:parameters.2.sourceCrsAxis = 0LL ;
		:parameters.2.unitName = "metre" ;
		:parameters.2.unitSiRatio = 1. ;
		:parameters.2.uncertaintyMeasure = "2SE" ;
		:parameters.3.parameterName = "longitudeOffsetUncertainty" ;
		:parameters.3.parameterSet = "offsetUncertainty" ;
		:parameters.3.sourceCrsAxis = 1LL ;
		:parameters.3.unitName = "metre" ;
		:parameters.3.unitSiRatio = 1. ;
		:parameters.3.uncertaintyMeasure = "2SE" ;
		:operationAccuracy = 1.5 ;
		:_NCProperties = "version=2,netcdf=4.9.0,hdf5=1.12.2" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: national_transformation_v2_0 {
  dimensions:
  	offsetCount = 2 ;
  	offsetUncertaintyCount = 2 ;

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: CAeast {
    dimensions:
    	iNodeCount = 529 ;
    	jNodeCount = 241 ;
    variables:
    	float offset(iNodeCount, jNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.0833333333333333, -88., 0.0833333333333333, 0. ;

    group: NFstjohn {
      dimensions:
      	iNodeCount = 81 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 47.8333333333333, 0., -0.00833333333333333, -53., 0.00833333333333333, 0. ;
      } // group NFstjohn

    group: ONkinstn {
      dimensions:
      	iNodeCount = 321 ;
      	jNodeCount = 321 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.5, 0., -0.00833333333333333, -78.8333333333333, 0.00833333333333333, 0. ;
      } // group ONkinstn

    group: ONottawa {
      dimensions:
      	iNodeCount = 221 ;
      	jNodeCount = 201 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 45.9166666666667, 0., -0.00833333333333333, -76.1666666666667, 0.00833333333333333, 0. ;
      } // group ONottawa

    group: ONsarnia {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 121 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 43.4166666666667, 0., -0.00833333333333333, -82.5833333333333, 0.00833333333333333, 0. ;
      } // group ONsarnia

    group: ONsault {
      dimensions:
      	iNodeCount = 351 ;
      	jNodeCount = 71 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.6666666666667, 0., -0.00833333333333333, -84.6666666666667, 0.00833333333333333, 0. ;
      } // group ONsault

    group: ONtimins {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.6666666666667, 0., -0.00833333333333333, -81.6666666666667, 0.00833333333333333, 0. ;
      } // group ONtimins

    group: ONtronto {
      dimensions:
      	iNodeCount = 351 ;
      	jNodeCount = 511 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.6666666666667, 0., -0.00833333333333333, -81.75, 0.00833333333333333, 0. ;
      } // group ONtronto

    group: ONwinsor {
      dimensions:
      	iNodeCount = 171 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 42.4166666666667, 0., -0.00833333333333333, -83.1666666666667, 0.00833333333333333, 0. ;
      } // group ONwinsor
    } // group CAeast

  group: CAwest {
    dimensions:
    	iNodeCount = 649 ;
    	jNodeCount = 157 ;
    variables:
    	float offset(iNodeCount, jNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.0833333333333333, -142., 0.0833333333333333, 0. ;

    group: ALbanff {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.25, 0., -0.00833333333333333, -115.583333333333, 0.00833333333333333, 0. ;
      } // group ALbanff

    group: ALbarhed {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.1666666666667, 0., -0.00833333333333333, -114.5, 0.00833333333333333, 0. ;
      } // group ALbarhed

    group: ALbonvil {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.3333333333333, 0., -0.00833333333333333, -110.833333333333, 0.00833333333333333, 0. ;
      } // group ALbonvil

    group: ALbowisl {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -111.5, 0.00833333333333333, 0. ;
      } // group ALbowisl

    group: ALbrooks {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.6666666666667, 0., -0.00833333333333333, -112., 0.00833333333333333, 0. ;
      } // group ALbrooks

    group: ALcalgry {
      dimensions:
      	iNodeCount = 101 ;
      	jNodeCount = 101 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.3333333333333, 0., -0.00833333333333333, -114.583333333333, 0.00833333333333333, 0. ;
      } // group ALcalgry

    group: ALcamros {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.0833333333333, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      } // group ALcamros

    group: ALcanmor {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.1666666666667, 0., -0.00833333333333333, -115.5, 0.00833333333333333, 0. ;
      } // group ALcanmor

    group: ALcardst {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -113.416666666667, 0.00833333333333333, 0. ;
      } // group ALcardst

    group: ALcarsta {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.6666666666667, 0., -0.00833333333333333, -114.25, 0.00833333333333333, 0. ;
      } // group ALcarsta

    group: ALclarho {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -113.666666666667, 0.00833333333333333, 0. ;
      } // group ALclarho

    group: ALcoldlk {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.5833333333333, 0., -0.00833333333333333, -110.333333333333, 0.00833333333333333, 0. ;
      } // group ALcoldlk

    group: ALcrowps {
      dimensions:
      	iNodeCount = 71 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.75, 0., -0.00833333333333333, -114.75, 0.00833333333333333, 0. ;
      } // group ALcrowps

    group: ALdraytn {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -115.083333333333, 0.00833333333333333, 0. ;
      } // group ALdraytn

    group: ALdrumhl {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.5833333333333, 0., -0.00833333333333333, -112.916666666667, 0.00833333333333333, 0. ;
      } // group ALdrumhl

    group: ALedmntn {
      dimensions:
      	iNodeCount = 131 ;
      	jNodeCount = 91 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.9166666666667, 0., -0.00833333333333333, -114.166666666667, 0.00833333333333333, 0. ;
      } // group ALedmntn

    group: ALedson {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.6666666666667, 0., -0.00833333333333333, -116.583333333333, 0.00833333333333333, 0. ;
      } // group ALedson

    group: ALfairvw {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.1666666666667, 0., -0.00833333333333333, -118.5, 0.00833333333333333, 0. ;
      } // group ALfairvw

    group: ALftmacl {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.8333333333333, 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      } // group ALftmacl

    group: ALftmcmr {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.8333333333333, 0., -0.00833333333333333, -111.583333333333, 0.00833333333333333, 0. ;
      } // group ALftmcmr

    group: ALgrcach {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54., 0., -0.00833333333333333, -119.25, 0.00833333333333333, 0. ;
      } // group ALgrcach

    group: ALgrimsh {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.25, 0., -0.00833333333333333, -117.666666666667, 0.00833333333333333, 0. ;
      } // group ALgrimsh

    group: ALgrprar {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.25, 0., -0.00833333333333333, -118.916666666667, 0.00833333333333333, 0. ;
      } // group ALgrprar

    group: ALhanna {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.75, 0., -0.00833333333333333, -112.083333333333, 0.00833333333333333, 0. ;
      } // group ALhanna

    group: ALhilevl {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 58.5833333333333, 0., -0.00833333333333333, -117.25, 0.00833333333333333, 0. ;
      } // group ALhilevl

    group: ALhinton {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.5, 0., -0.00833333333333333, -117.666666666667, 0.00833333333333333, 0. ;
      } // group ALhinton

    group: ALhiprai {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.5, 0., -0.00833333333333333, -116.666666666667, 0.00833333333333333, 0. ;
      } // group ALhiprai

    group: ALinnsfl {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.1666666666667, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      } // group ALinnsfl

    group: ALjasper {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -118.166666666667, 0.00833333333333333, 0. ;
      } // group ALjasper

    group: ALlacbic {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.8333333333333, 0., -0.00833333333333333, -112.083333333333, 0.00833333333333333, 0. ;
      } // group ALlacbic

    group: ALlacomb {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.5833333333333, 0., -0.00833333333333333, -113.833333333333, 0.00833333333333333, 0. ;
      } // group ALlacomb

    group: ALletbrg {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      } // group ALletbrg

    group: ALlkloui {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.5, 0., -0.00833333333333333, -116.25, 0.00833333333333333, 0. ;
      } // group ALlkloui

    group: ALlydmin {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -110.166666666667, 0.00833333333333333, 0. ;
      } // group ALlydmin

    group: ALmedhat {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.1666666666667, 0., -0.00833333333333333, -110.833333333333, 0.00833333333333333, 0. ;
      } // group ALmedhat

    group: ALolds {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.9166666666667, 0., -0.00833333333333333, -114.25, 0.00833333333333333, 0. ;
      } // group ALolds

    group: ALoyen {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.4166666666667, 0., -0.00833333333333333, -110.583333333333, 0.00833333333333333, 0. ;
      } // group ALoyen

    group: ALpeacer {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.3333333333333, 0., -0.00833333333333333, -117.416666666667, 0.00833333333333333, 0. ;
      } // group ALpeacer

    group: ALpinchr {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      } // group ALpinchr

    group: ALponoka {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.75, 0., -0.00833333333333333, -113.666666666667, 0.00833333333333333, 0. ;
      } // group ALponoka

    group: ALraymnd {
      dimensions:
      	iNodeCount = 51 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      } // group ALraymnd

    group: ALredeer {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.4166666666667, 0., -0.00833333333333333, -113.916666666667, 0.00833333333333333, 0. ;
      } // group ALredeer

    group: ALrockmt {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.5, 0., -0.00833333333333333, -115., 0.00833333333333333, 0. ;
      } // group ALrockmt

    group: ALslavlk {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.3333333333333, 0., -0.00833333333333333, -114.916666666667, 0.00833333333333333, 0. ;
      } // group ALslavlk

    group: ALstetlr {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.4166666666667, 0., -0.00833333333333333, -112.833333333333, 0.00833333333333333, 0. ;
      } // group ALstetlr

    group: ALstpaul {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.0833333333333, 0., -0.00833333333333333, -111.416666666667, 0.00833333333333333, 0. ;
      } // group ALstpaul

    group: ALstramr {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.1666666666667, 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      } // group ALstramr

    group: ALswanhi {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.8333333333333, 0., -0.00833333333333333, -115.583333333333, 0.00833333333333333, 0. ;
      } // group ALswanhi

    group: ALtaber {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -112.25, 0.00833333333333333, 0. ;
      } // group ALtaber

    group: ALtrehil {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.75, 0., -0.00833333333333333, -113.333333333333, 0.00833333333333333, 0. ;
      } // group ALtrehil

    group: ALvegvil {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.5833333333333, 0., -0.00833333333333333, -112.166666666667, 0.00833333333333333, 0. ;
      } // group ALvegvil

    group: ALvermil {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.4166666666667, 0., -0.00833333333333333, -111., 0.00833333333333333, 0. ;
      } // group ALvermil

    group: ALwanwgt {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -111., 0.00833333333333333, 0. ;
      } // group ALwanwgt

    group: ALweslok {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.25, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      } // group ALweslok

    group: ALwetask {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53., 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      } // group ALwetask

    group: ALwhitec {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.1666666666667, 0., -0.00833333333333333, -115.833333333333, 0.00833333333333333, 0. ;
      } // group ALwhitec

    group: BCcambel {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -125.333333333333, 0.00833333333333333, 0. ;
      } // group BCcambel

    group: BCcranbk {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -115.833333333333, 0.00833333333333333, 0. ;
      } // group BCcranbk

    group: BCdawson {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.8333333333333, 0., -0.00833333333333333, -120.333333333333, 0.00833333333333333, 0. ;
      } // group BCdawson

    group: BCelkfrd {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -115., 0.00833333333333333, 0. ;
      } // group BCelkfrd

    group: BCfield {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.4166666666667, 0., -0.00833333333333333, -116.583333333333, 0.00833333333333333, 0. ;
      } // group BCfield

    group: BCgranil {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.9166666666667, 0., -0.00833333333333333, -126.25, 0.00833333333333333, 0. ;
      } // group BCgranil

    group: BCkamlop {
      dimensions:
      	iNodeCount = 51 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.75, 0., -0.00833333333333333, -120.5, 0.00833333333333333, 0. ;
      } // group BCkamlop

    group: BCkelwna {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -119.583333333333, 0.00833333333333333, 0. ;
      } // group BCkelwna

    group: BClogan {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5, 0., -0.00833333333333333, -120.833333333333, 0.00833333333333333, 0. ;
      } // group BClogan

    group: BCmacknz {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.4166666666667, 0., -0.00833333333333333, -123.166666666667, 0.00833333333333333, 0. ;
      } // group BCmacknz

    group: BCnanimo {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -124.083333333333, 0.00833333333333333, 0. ;
      } // group BCnanimo

    group: BCnelson {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -117.333333333333, 0.00833333333333333, 0. ;
      } // group BCnelson

    group: BCparkvl {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.3333333333333, 0., -0.00833333333333333, -124.416666666667, 0.00833333333333333, 0. ;
      } // group BCparkvl

    group: BCpentic {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -119.666666666667, 0.00833333333333333, 0. ;
      } // group BCpentic

    group: BCportal {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.3333333333333, 0., -0.00833333333333333, -124.833333333333, 0.00833333333333333, 0. ;
      } // group BCportal

    group: BCpowell {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -124.583333333333, 0.00833333333333333, 0. ;
      } // group BCpowell

    group: BCprigeo {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.0833333333333, 0., -0.00833333333333333, -122.916666666667, 0.00833333333333333, 0. ;
      } // group BCprigeo

    group: BCroslnd {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.0833333333333, 0., -0.00833333333333333, -117.833333333333, 0.00833333333333333, 0. ;
      } // group BCroslnd

    group: BCtrail {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.1666666666667, 0., -0.00833333333333333, -117.75, 0.00833333333333333, 0. ;
      } // group BCtrail

    group: BCtumblr {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.1666666666667, 0., -0.00833333333333333, -121.083333333333, 0.00833333333333333, 0. ;
      } // group BCtumblr

    group: BCvancvr {
      dimensions:
      	iNodeCount = 131 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.4166666666667, 0., -0.00833333333333333, -123.25, 0.00833333333333333, 0. ;
      } // group BCvancvr

    group: BCvernon {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.3333333333333, 0., -0.00833333333333333, -119.333333333333, 0.00833333333333333, 0. ;
      } // group BCvernon

    group: BCvictor {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.75, 0., -0.00833333333333333, -123.583333333333, 0.00833333333333333, 0. ;
      } // group BCvictor

    group: ONthundr {
      dimensions:
      	iNodeCount = 71 ;
      	jNodeCount = 51 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.5833333333333, 0., -0.00833333333333333, -89.5833333333333, 0.00833333333333333, 0. ;
      } // group ONthundr

    group: SAestvan {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -103.083333333333, 0.00833333333333333, 0. ;
      } // group SAestvan

    group: SAmelfrt {
      dimensions:
      	iNodeCount = 71 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -104.666666666667, 0.00833333333333333, 0. ;
      } // group SAmelfrt

    group: SAmelvil {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51., 0., -0.00833333333333333, -102.916666666667, 0.00833333333333333, 0. ;
      } // group SAmelvil

    group: SAmosjaw {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5, 0., -0.00833333333333333, -105.75, 0.00833333333333333, 0. ;
      } // group SAmosjaw

    group: SAnbatle {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.8333333333333, 0., -0.00833333333333333, -108.416666666667, 0.00833333333333333, 0. ;
      } // group SAnbatle

    group: SApralbt {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -106., 0.00833333333333333, 0. ;
      } // group SApralbt

    group: SAregina {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5833333333333, 0., -0.00833333333333333, -104.75, 0.00833333333333333, 0. ;
      } // group SAregina

    group: SAsatoon {
      dimensions:
      	iNodeCount = 51 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.25, 0., -0.00833333333333333, -106.833333333333, 0.00833333333333333, 0. ;
      } // group SAsatoon

    group: SAswiftc {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.4166666666667, 0., -0.00833333333333333, -107.916666666667, 0.00833333333333333, 0. ;
      } // group SAswiftc

    group: SAweybrn {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.75, 0., -0.00833333333333333, -103.916666666667, 0.00833333333333333, 0. ;
      } // group SAweybrn

    group: SAyorktn {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.3333333333333, 0., -0.00833333333333333, -102.583333333333, 0.00833333333333333, 0. ;
      } // group SAyorktn
    } // group CAwest

  group: CAnorth {
    dimensions:
    	iNodeCount = 589 ;
    	jNodeCount = 181 ;
    variables:
    	float offset(iNodeCount, jNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 75., 0., -0.0833333333333333, -142., 0.166666666666667, 0. ;

    group: NWclyder {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 31 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 70.5833333333333, 0., -0.00833333333333333, -68.8333333333333, 0.0166666666666667, 0. ;
      } // group NWclyder

    group: NWftgood {
      dimensions:
      	iNodeCount = 21 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 66.3333333333333, 0., -0.00833333333333333, -128.833333333333, 0.0166666666666667, 0. ;
      } // group NWftgood

    group: NWhayriv {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 61., 0., -0.00833333333333333, -116.5, 0.0166666666666667, 0. ;
      } // group NWhayriv

    group: NWinuvik {
      dimensions:
      	iNodeCount = 31 ;
      	jNodeCount = 41 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 68.5, 0., -0.00833333333333333, -133.833333333333, 0.0166666666666667, 0. ;
      } // group NWinuvik

    group: NWiqulit {
      dimensions:
      	iNodeCount = 61 ;
      	jNodeCount = 61 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 64., 0., -0.00833333333333333, -69., 0.0166666666666667, 0. ;
      } // group NWiqulit

    group: NWpondin {
      dimensions:
      	iNodeCount = 41 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 72.75, 0., -0.00833333333333333, -78.1666666666667, 0.0166666666666667, 0. ;
      } // group NWpondin

    group: NWrankin {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.9166666666667, 0., -0.00833333333333333, -92.1666666666667, 0.0166666666666667, 0. ;
      } // group NWrankin

    group: NWyellow {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.5, 0., -0.00833333333333333, -114.5, 0.0166666666666667, 0. ;
      } // group NWyellow

    group: YUdawson {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 64.1666666666667, 0., -0.00833333333333333, -139.5, 0.0166666666666667, 0. ;
      } // group YUdawson

    group: YUrossri {
      dimensions:
      	iNodeCount = 11 ;
      	jNodeCount = 21 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.0833333333333, 0., -0.00833333333333333, -132.583333333333, 0.0166666666666667, 0. ;
      } // group YUrossri

    group: YUwhiteh {
      dimensions:
      	iNodeCount = 6 ;
      	jNodeCount = 11 ;
      variables:
      	float offset(iNodeCount, jNodeCount, offsetCount) ;
      		offset:_Storage = "contiguous" ;
      		offset:_Endianness = "little" ;
      	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
      		offsetUncertainty:_Storage = "contiguous" ;
      		offsetUncertainty:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 60.75, 0., -0.00833333333333333, -135.083333333333, 0.0166666666666667, 0. ;
      } // group YUwhiteh
    } // group CAnorth

  group: CAarctic {
    dimensions:
    	iNodeCount = 295 ;
    	jNodeCount = 109 ;
    variables:
    	float offset(iNodeCount, jNodeCount, offsetCount) ;
    		offset:_Storage = "contiguous" ;
    		offset:_Endianness = "little" ;
    	float offsetUncertainty(iNodeCount, jNodeCount, offsetUncertaintyCount) ;
    		offsetUncertainty:_Storage = "contiguous" ;
    		offsetUncertainty:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 84., 0., -0.0833333333333333, -142., 0.333333333333333, 0. ;
    } // group CAarctic
  } // group national_transformation_v2_0
}

netcdf ca_ntv2 {
types:
  compound ggxfParameterType {
    char parameterName(32) ;
    char parameterSet(32) ;
    char unit(16) ;
    double unitSiRatio ;
    int sourceCrsAxis ;
    float parameterMinimumValue ;
    float parameterMaximumValue ;
    float noDataFlag ;
  }; // ggxfParameterType

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "27to83.gxt" ;
		:title = "Canadian National NAD27-NAD83(Original) NTV2 transformation" ;
		:summary = "Canadian National NAD27-NAD83(Original) NTV2 transformation" ;
		:content = "geographic2dOffsets" ;
		:product_version = "National Transformation v2_0" ;
		:date_issued = "1995-02" ;
		:publisher_institution = "Geodetic Survey Division, Natural Resources Canada" ;
		:publisher_url = "https://webapp.geod.nrcan.gc.ca/geod/data-donnees/transformations.php" ;
		:license = "https://open.canada.ca/en/open-government-licence-canada" ;
		:geospatial_lat_min = 40. ;
		:geospatial_lon_min = -141. ;
		:geospatial_lat_max = 60. ;
		:geospatial_lon_max = -88. ;
		:extent_description = "Canada south of 60°N" ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD27\",\n  DATUM[\"North American Datum 1927\",\n    ELLIPSOID[\"Clarke 1866\",6378206.4,294.9786982,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:targetCrsWkt = "GEOGCRS[\"NAD83(Original)\",\n  DATUM[\"North American Datum 1983\",\n    ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		ggxfParameterType :parameters = 
    {{"latitudeOffset"}, {"offset"}, {"arc-second"}, 4.84813681109536e-06, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"longitudeOffset"}, {"offset"}, {"arc-second"}, 4.84813681109536e-06, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"latitudeOffsetUncertainty"}, {"offsetUncertainty"}, {"metre"}, 1, 0, -3.402823e+38, -3.402823e+38, -3.402823e+38}, 
    {{"longitudeOffsetUncertainty"}, {"offsetUncertainty"}, {"metre"}, 1, 1, -3.402823e+38, -3.402823e+38, -3.402823e+38} ;
		:operationAccuracy = 1.5 ;
		:uncertaintyMeasure = "2CEE" ;
		:_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.12.0," ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;

group: national_transformation_v2_0 {
  dimensions:
  	parameter = 4 ;

  // group attributes:
  		:interpolationMethod = "bilinear" ;

  group: CAeast {
    dimensions:
    	gridi = 529 ;
    	gridj = 241 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.0833333333333333, -88., 0.0833333333333333, 0. ;
    		:iNodeCount = 529LL ;
    		:jNodeCount = 241LL ;

    group: NFstjohn {
      dimensions:
      	gridi = 81 ;
      	gridj = 51 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 47.8333333333333, 0., -0.00833333333333333, -53., 0.00833333333333333, 0. ;
      		:iNodeCount = 81LL ;
      		:jNodeCount = 51LL ;
      } // group NFstjohn

    group: ONkinstn {
      dimensions:
      	gridi = 321 ;
      	gridj = 321 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.5, 0., -0.00833333333333333, -78.8333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 321LL ;
      		:jNodeCount = 321LL ;
      } // group ONkinstn

    group: ONottawa {
      dimensions:
      	gridi = 221 ;
      	gridj = 201 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 45.9166666666667, 0., -0.00833333333333333, -76.1666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 221LL ;
      		:jNodeCount = 201LL ;
      } // group ONottawa

    group: ONsarnia {
      dimensions:
      	gridi = 101 ;
      	gridj = 121 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 43.4166666666667, 0., -0.00833333333333333, -82.5833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 101LL ;
      		:jNodeCount = 121LL ;
      } // group ONsarnia

    group: ONsault {
      dimensions:
      	gridi = 351 ;
      	gridj = 71 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.6666666666667, 0., -0.00833333333333333, -84.6666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 351LL ;
      		:jNodeCount = 71LL ;
      } // group ONsault

    group: ONtimins {
      dimensions:
      	gridi = 101 ;
      	gridj = 41 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.6666666666667, 0., -0.00833333333333333, -81.6666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 101LL ;
      		:jNodeCount = 41LL ;
      } // group ONtimins

    group: ONtronto {
      dimensions:
      	gridi = 351 ;
      	gridj = 511 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 46.6666666666667, 0., -0.00833333333333333, -81.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 351LL ;
      		:jNodeCount = 511LL ;
      } // group ONtronto

    group: ONwinsor {
      dimensions:
      	gridi = 171 ;
      	gridj = 61 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 42.4166666666667, 0., -0.00833333333333333, -83.1666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 171LL ;
      		:jNodeCount = 61LL ;
      } // group ONwinsor
    } // group CAeast

  group: CAwest {
    dimensions:
    	gridi = 649 ;
    	gridj = 157 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 60., 0., -0.0833333333333333, -142., 0.0833333333333333, 0. ;
    		:iNodeCount = 649LL ;
    		:jNodeCount = 157LL ;

    group: ALbanff {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.25, 0., -0.00833333333333333, -115.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group ALbanff

    group: ALbarhed {
      dimensions:
      	gridi = 21 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.1666666666667, 0., -0.00833333333333333, -114.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      } // group ALbarhed

    group: ALbonvil {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.3333333333333, 0., -0.00833333333333333, -110.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALbonvil

    group: ALbowisl {
      dimensions:
      	gridi = 31 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -111.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 11LL ;
      } // group ALbowisl

    group: ALbrooks {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.6666666666667, 0., -0.00833333333333333, -112., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALbrooks

    group: ALcalgry {
      dimensions:
      	gridi = 101 ;
      	gridj = 101 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.3333333333333, 0., -0.00833333333333333, -114.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 101LL ;
      		:jNodeCount = 101LL ;
      } // group ALcalgry

    group: ALcamros {
      dimensions:
      	gridi = 41 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.0833333333333, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 31LL ;
      } // group ALcamros

    group: ALcanmor {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.1666666666667, 0., -0.00833333333333333, -115.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALcanmor

    group: ALcardst {
      dimensions:
      	gridi = 31 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -113.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 11LL ;
      } // group ALcardst

    group: ALcarsta {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.6666666666667, 0., -0.00833333333333333, -114.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALcarsta

    group: ALclarho {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -113.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALclarho

    group: ALcoldlk {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.5833333333333, 0., -0.00833333333333333, -110.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group ALcoldlk

    group: ALcrowps {
      dimensions:
      	gridi = 71 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.75, 0., -0.00833333333333333, -114.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 71LL ;
      		:jNodeCount = 31LL ;
      } // group ALcrowps

    group: ALdraytn {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -115.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group ALdraytn

    group: ALdrumhl {
      dimensions:
      	gridi = 61 ;
      	gridj = 41 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.5833333333333, 0., -0.00833333333333333, -112.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 41LL ;
      } // group ALdrumhl

    group: ALedmntn {
      dimensions:
      	gridi = 131 ;
      	gridj = 91 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.9166666666667, 0., -0.00833333333333333, -114.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 131LL ;
      		:jNodeCount = 91LL ;
      } // group ALedmntn

    group: ALedson {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.6666666666667, 0., -0.00833333333333333, -116.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group ALedson

    group: ALfairvw {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.1666666666667, 0., -0.00833333333333333, -118.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group ALfairvw

    group: ALftmacl {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.8333333333333, 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALftmacl

    group: ALftmcmr {
      dimensions:
      	gridi = 61 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.8333333333333, 0., -0.00833333333333333, -111.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 31LL ;
      } // group ALftmcmr

    group: ALgrcach {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54., 0., -0.00833333333333333, -119.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALgrcach

    group: ALgrimsh {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.25, 0., -0.00833333333333333, -117.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group ALgrimsh

    group: ALgrprar {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.25, 0., -0.00833333333333333, -118.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group ALgrprar

    group: ALhanna {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.75, 0., -0.00833333333333333, -112.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALhanna

    group: ALhilevl {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 58.5833333333333, 0., -0.00833333333333333, -117.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALhilevl

    group: ALhinton {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.5, 0., -0.00833333333333333, -117.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALhinton

    group: ALhiprai {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.5, 0., -0.00833333333333333, -116.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group ALhiprai

    group: ALinnsfl {
      dimensions:
      	gridi = 21 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.1666666666667, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 31LL ;
      } // group ALinnsfl

    group: ALjasper {
      dimensions:
      	gridi = 21 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -118.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      } // group ALjasper

    group: ALlacbic {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.8333333333333, 0., -0.00833333333333333, -112.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALlacbic

    group: ALlacomb {
      dimensions:
      	gridi = 31 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.5833333333333, 0., -0.00833333333333333, -113.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 11LL ;
      } // group ALlacomb

    group: ALletbrg {
      dimensions:
      	gridi = 61 ;
      	gridj = 41 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 41LL ;
      } // group ALletbrg

    group: ALlkloui {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.5, 0., -0.00833333333333333, -116.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group ALlkloui

    group: ALlydmin {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -110.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALlydmin

    group: ALmedhat {
      dimensions:
      	gridi = 41 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.1666666666667, 0., -0.00833333333333333, -110.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 31LL ;
      } // group ALmedhat

    group: ALolds {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.9166666666667, 0., -0.00833333333333333, -114.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALolds

    group: ALoyen {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.4166666666667, 0., -0.00833333333333333, -110.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALoyen

    group: ALpeacer {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 56.3333333333333, 0., -0.00833333333333333, -117.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group ALpeacer

    group: ALpinchr {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group ALpinchr

    group: ALponoka {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.75, 0., -0.00833333333333333, -113.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group ALponoka

    group: ALraymnd {
      dimensions:
      	gridi = 51 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5, 0., -0.00833333333333333, -113., 0.00833333333333333, 0. ;
      		:iNodeCount = 51LL ;
      		:jNodeCount = 21LL ;
      } // group ALraymnd

    group: ALredeer {
      dimensions:
      	gridi = 41 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.4166666666667, 0., -0.00833333333333333, -113.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 31LL ;
      } // group ALredeer

    group: ALrockmt {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.5, 0., -0.00833333333333333, -115., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group ALrockmt

    group: ALslavlk {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.3333333333333, 0., -0.00833333333333333, -114.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALslavlk

    group: ALstetlr {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.4166666666667, 0., -0.00833333333333333, -112.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALstetlr

    group: ALstpaul {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.0833333333333, 0., -0.00833333333333333, -111.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALstpaul

    group: ALstramr {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.1666666666667, 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALstramr

    group: ALswanhi {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.8333333333333, 0., -0.00833333333333333, -115.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group ALswanhi

    group: ALtaber {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -112.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALtaber

    group: ALtrehil {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.75, 0., -0.00833333333333333, -113.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group ALtrehil

    group: ALvegvil {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.5833333333333, 0., -0.00833333333333333, -112.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALvegvil

    group: ALvermil {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.4166666666667, 0., -0.00833333333333333, -111., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALvermil

    group: ALwanwgt {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -111., 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALwanwgt

    group: ALweslok {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.25, 0., -0.00833333333333333, -114., 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group ALweslok

    group: ALwetask {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53., 0., -0.00833333333333333, -113.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group ALwetask

    group: ALwhitec {
      dimensions:
      	gridi = 41 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.1666666666667, 0., -0.00833333333333333, -115.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 11LL ;
      } // group ALwhitec

    group: BCcambel {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -125.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCcambel

    group: BCcranbk {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -115.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCcranbk

    group: BCdawson {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.8333333333333, 0., -0.00833333333333333, -120.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCdawson

    group: BCelkfrd {
      dimensions:
      	gridi = 21 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -115., 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      } // group BCelkfrd

    group: BCfield {
      dimensions:
      	gridi = 21 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.4166666666667, 0., -0.00833333333333333, -116.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      } // group BCfield

    group: BCgranil {
      dimensions:
      	gridi = 11 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.9166666666667, 0., -0.00833333333333333, -126.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      } // group BCgranil

    group: BCkamlop {
      dimensions:
      	gridi = 51 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.75, 0., -0.00833333333333333, -120.5, 0.00833333333333333, 0. ;
      		:iNodeCount = 51LL ;
      		:jNodeCount = 21LL ;
      } // group BCkamlop

    group: BCkelwna {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.0833333333333, 0., -0.00833333333333333, -119.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group BCkelwna

    group: BClogan {
      dimensions:
      	gridi = 11 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5, 0., -0.00833333333333333, -120.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      } // group BClogan

    group: BCmacknz {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.4166666666667, 0., -0.00833333333333333, -123.166666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCmacknz

    group: BCnanimo {
      dimensions:
      	gridi = 61 ;
      	gridj = 61 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -124.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 61LL ;
      } // group BCnanimo

    group: BCnelson {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -117.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group BCnelson

    group: BCparkvl {
      dimensions:
      	gridi = 21 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.3333333333333, 0., -0.00833333333333333, -124.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      } // group BCparkvl

    group: BCpentic {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.5833333333333, 0., -0.00833333333333333, -119.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCpentic

    group: BCportal {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.3333333333333, 0., -0.00833333333333333, -124.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group BCportal

    group: BCpowell {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.9166666666667, 0., -0.00833333333333333, -124.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCpowell

    group: BCprigeo {
      dimensions:
      	gridi = 41 ;
      	gridj = 41 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 54.0833333333333, 0., -0.00833333333333333, -122.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 41LL ;
      } // group BCprigeo

    group: BCroslnd {
      dimensions:
      	gridi = 11 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.0833333333333, 0., -0.00833333333333333, -117.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      } // group BCroslnd

    group: BCtrail {
      dimensions:
      	gridi = 11 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.1666666666667, 0., -0.00833333333333333, -117.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      } // group BCtrail

    group: BCtumblr {
      dimensions:
      	gridi = 21 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 55.1666666666667, 0., -0.00833333333333333, -121.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 11LL ;
      } // group BCtumblr

    group: BCvancvr {
      dimensions:
      	gridi = 131 ;
      	gridj = 51 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.4166666666667, 0., -0.00833333333333333, -123.25, 0.00833333333333333, 0. ;
      		:iNodeCount = 131LL ;
      		:jNodeCount = 51LL ;
      } // group BCvancvr

    group: BCvernon {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.3333333333333, 0., -0.00833333333333333, -119.333333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group BCvernon

    group: BCvictor {
      dimensions:
      	gridi = 41 ;
      	gridj = 51 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.75, 0., -0.00833333333333333, -123.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 51LL ;
      } // group BCvictor

    group: ONthundr {
      dimensions:
      	gridi = 71 ;
      	gridj = 51 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 48.5833333333333, 0., -0.00833333333333333, -89.5833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 71LL ;
      		:jNodeCount = 51LL ;
      } // group ONthundr

    group: SAestvan {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.25, 0., -0.00833333333333333, -103.083333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group SAestvan

    group: SAmelfrt {
      dimensions:
      	gridi = 71 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.9166666666667, 0., -0.00833333333333333, -104.666666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 71LL ;
      		:jNodeCount = 21LL ;
      } // group SAmelfrt

    group: SAmelvil {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51., 0., -0.00833333333333333, -102.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group SAmelvil

    group: SAmosjaw {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5, 0., -0.00833333333333333, -105.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group SAmosjaw

    group: SAnbatle {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.8333333333333, 0., -0.00833333333333333, -108.416666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group SAnbatle

    group: SApralbt {
      dimensions:
      	gridi = 61 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 53.3333333333333, 0., -0.00833333333333333, -106., 0.00833333333333333, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 31LL ;
      } // group SApralbt

    group: SAregina {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.5833333333333, 0., -0.00833333333333333, -104.75, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group SAregina

    group: SAsatoon {
      dimensions:
      	gridi = 51 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 52.25, 0., -0.00833333333333333, -106.833333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 51LL ;
      		:jNodeCount = 31LL ;
      } // group SAsatoon

    group: SAswiftc {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 50.4166666666667, 0., -0.00833333333333333, -107.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group SAswiftc

    group: SAweybrn {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 49.75, 0., -0.00833333333333333, -103.916666666667, 0.00833333333333333, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group SAweybrn

    group: SAyorktn {
      dimensions:
      	gridi = 31 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 51.3333333333333, 0., -0.00833333333333333, -102.583333333333, 0.00833333333333333, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 21LL ;
      } // group SAyorktn
    } // group CAwest

  group: CAnorth {
    dimensions:
    	gridi = 589 ;
    	gridj = 181 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 75., 0., -0.0833333333333333, -142., 0.166666666666667, 0. ;
    		:iNodeCount = 589LL ;
    		:jNodeCount = 181LL ;

    group: NWclyder {
      dimensions:
      	gridi = 31 ;
      	gridj = 31 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 70.5833333333333, 0., -0.00833333333333333, -68.8333333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 31LL ;
      } // group NWclyder

    group: NWftgood {
      dimensions:
      	gridi = 21 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 66.3333333333333, 0., -0.00833333333333333, -128.833333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 21LL ;
      		:jNodeCount = 21LL ;
      } // group NWftgood

    group: NWhayriv {
      dimensions:
      	gridi = 61 ;
      	gridj = 61 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 61., 0., -0.00833333333333333, -116.5, 0.0166666666666667, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 61LL ;
      } // group NWhayriv

    group: NWinuvik {
      dimensions:
      	gridi = 31 ;
      	gridj = 41 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 68.5, 0., -0.00833333333333333, -133.833333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 31LL ;
      		:jNodeCount = 41LL ;
      } // group NWinuvik

    group: NWiqulit {
      dimensions:
      	gridi = 61 ;
      	gridj = 61 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 64., 0., -0.00833333333333333, -69., 0.0166666666666667, 0. ;
      		:iNodeCount = 61LL ;
      		:jNodeCount = 61LL ;
      } // group NWiqulit

    group: NWpondin {
      dimensions:
      	gridi = 41 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 72.75, 0., -0.00833333333333333, -78.1666666666667, 0.0166666666666667, 0. ;
      		:iNodeCount = 41LL ;
      		:jNodeCount = 21LL ;
      } // group NWpondin

    group: NWrankin {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.9166666666667, 0., -0.00833333333333333, -92.1666666666667, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group NWrankin

    group: NWyellow {
      dimensions:
      	gridi = 11 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.5, 0., -0.00833333333333333, -114.5, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 11LL ;
      } // group NWyellow

    group: YUdawson {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 64.1666666666667, 0., -0.00833333333333333, -139.5, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group YUdawson

    group: YUrossri {
      dimensions:
      	gridi = 11 ;
      	gridj = 21 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 62.0833333333333, 0., -0.00833333333333333, -132.583333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 11LL ;
      		:jNodeCount = 21LL ;
      } // group YUrossri

    group: YUwhiteh {
      dimensions:
      	gridi = 6 ;
      	gridj = 11 ;
      variables:
      	float data(gridj, gridi, parameter) ;
      		data:_Storage = "contiguous" ;
      		data:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = 60.75, 0., -0.00833333333333333, -135.083333333333, 0.0166666666666667, 0. ;
      		:iNodeCount = 6LL ;
      		:jNodeCount = 11LL ;
      } // group YUwhiteh
    } // group CAnorth

  group: CAarctic {
    dimensions:
    	gridi = 295 ;
    	gridj = 109 ;
    variables:
    	float data(gridj, gridi, parameter) ;
    		data:_Storage = "contiguous" ;
    		data:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = 84., 0., -0.0833333333333333, -142., 0.333333333333333, 0. ;
    		:iNodeCount = 295LL ;
    		:jNodeCount = 109LL ;
    } // group CAarctic
  } // group national_transformation_v2_0
}

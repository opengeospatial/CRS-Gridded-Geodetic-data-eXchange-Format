netcdf PRGEOID18b {

// global attributes:
		:ggxfVersion = "1.0" ;
		:filename = "g2018pr.yaml" ;
		:content = "geoidModel" ;
		:remark = "hybrid geoid" ;
		:contentApplicabilityExtent.boundingBox.southBoundLatitude = 17.87 ;
		:contentApplicabilityExtent.boundingBox.westBoundLongitude = -68. ;
		:contentApplicabilityExtent.boundingBox.northBoundLatitude = 18.53 ;
		:contentApplicabilityExtent.boundingBox.eastBoundLongitude = -65. ;
		:contentApplicabilityExtent.extentDescription = "Puerto Rico - onshore." ;
		:interpolationCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,2],\n  AXIS[\"Geodetic latitude (Lat)\",north],\n  AXIS[\"Geodetic longitude (Lon)\",east],\n  ANGLEUNIT[\"degree\",0.0174532925199433]]\n" ;
		:sourceCrsWkt = "GEOGCRS[\"NAD83 (2011)\",\n  DATUM[\"North American Datum 1983 (2011) epoch 2010.00\",\n      ELLIPSOID[\"GRS 1980\",6378137.0,298.2572221,LENGTHUNIT[\"metre\",1]]],\n  CS[ellipsoidal,3],\n  AXIS[\"Geodetic latitude (Lat)\",north,\n    ANGLEUNIT[\"degree\",0.0174532925199433]],\n  AXIS[\"Geodetic longitude (Lon)\",east,\n    ANGLEUNIT[\"degree\",0.0174532925199433]],\n  AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1]]]\n" ;
		:targetCrsWkt = "VERTCRS[\"PRVD02 - NOHt\",\n  VDATUM[\"Puerto Rico Vertical Datum of 2002\"],\n  CS[vertical,1],\n  AXIS[\"Gravity-related height (H)\",up],\n  LENGTHUNIT[\"metre\",1]]\n" ;
		:operationAccuracy = 0.015 ;
		:organisationName = "National Geodetic Survey, National Oceanic and Atmospheric Administration." ;
		:deliveryPoint = "1315 East West Hwy" ;
		:city = "Silver Spring" ;
		:postalCode = "20910" ;
		:country = "United States of America" ;
		:onlineResourceLinkage = "https://geodesy.noaa.gov/PC_PROD/GEOID18/Format_ascii/g2018p0.asc.zip" ;

group: puerto_rico_virgin_islands_geoid18 {
  dimensions:
  	parameter = 1 ;

  // group attributes:
  		:parameters.count = 1LL ;
  		:parameters.0.parameterName = "geoidHeight" ;
  		:parameters.0.lengthUnit = "metre" ;
  		:parameters.0.unitSiRatio = 1. ;
  		:interpolationMethod = "biquadratic" ;

  group: puerto_rico_virgin_islands_geoid18 {
    dimensions:
    	gridi = 301 ;
    	gridj = 361 ;
    variables:
    	float data(gridj, gridi, parameter) ;

    // group attributes:
    		:iNodeCount = 301LL ;
    		:jNodeCount = 361LL ;
    		:remark = "grid starts in the top left (northwest) corner and works across (east) and down (south)" ;
    		:affineCoeffs = 21., 0., -0.01666666667, -69., 0.01666666667, 0. ;
    data:

     data =
  -48.7831,
  -48.8003,
  -48.8168,
  -48.8321,
  -48.8453,
  -48.8568,
  -48.8663,
  -48.8735,
  -48.8791,
  -48.8833,
  -48.8862,
  -48.8886,
  -48.8907,
  -48.8923,
  -48.8933,
  -48.8938,
  -48.8931,
  -48.8929,
  -48.8926,
  -48.8919,
  -48.8922,
  -48.8922,
  -48.8917,
  -48.8903,
  -48.8879,
  -48.8844,
  -48.8798,
  -48.8743,
  -48.8683,
  -48.8624,
  -48.8573,
  -48.8537,
  -48.8525,
  -48.8542,
  -48.8584,
  -48.8667,
  -48.8774,
  -48.8898,
  -48.9028,
  -48.9162,
  -48.9298,
  -48.9438,
  -48.9584,
  -48.9733,
  -48.9883,
  -49.003,
  -49.0166,
  -49.0286,
  -49.0385,
  -49.047,
  -49.0526,
  -49.0582,
  -49.0629,
  -49.0676,
  -49.0728,
  -49.0791,
  -49.0865,
  -49.0948,
  -49.1037,
  -49.1125,
  -49.1201,
  -49.126,
  -49.1295,
  -49.1306,
  -49.1294,
  -49.1257,
  -49.1197,
  -49.1104,
  -49.1,
  -49.088,
  -49.0744,
  -49.0592,
  -49.0424,
  -49.0245,
  -49.0059,
  -48.9872,
  -48.969,
  -48.9515,
  -48.9355,
  -48.9211,
  -48.9088,
  -48.8982,
  -48.8893,
  -48.8817,
  -48.8752,
  -48.8685,
  -48.864,
  -48.8602,
  -48.8571,
  -48.8542,
  -48.851,
  -48.8469,
  -48.8416,
  -48.8352,
  -48.8278,
  -48.8201,
  -48.8127,
  -48.8062,
  -48.8011,
  -48.7974,
  -48.7952,
  -48.7944,
  -48.7946,
  -48.7957,
  -48.7962,
  -48.7978,
  -48.7996,
  -48.8018,
  -48.8044,
  -48.8072,
  -48.8099,
  -48.8123,
  -48.8144,
  -48.8158,
  -48.8165,
  -48.817,
  -48.8177,
  -48.8191,
  -48.8218,
  -48.8264,
  -48.8333,
  -48.8423,
  -48.8531,
  -48.8651,
  -48.8769,
  -48.8904,
  -48.9049,
  -48.9207,
  -48.9382,
  -48.9576,
  -48.979,
  -49.0022,
  -49.0266,
  -49.0516,
  -49.0764,
  -49.1003,
  -49.1225,
  -49.1429,
  -49.1616,
  -49.1785,
  -49.1941,
  -49.2086,
  -49.2226,
  -49.2367,
  -49.2512,
  -49.2662,
  -49.2806,
  -49.2963,
  -49.3121,
  -49.3283,
  -49.3447,
  -49.3618,
  -49.3792,
  -49.3975,
  -49.4166,
  -49.4365,
  -49.457,
  -49.4778,
  -49.4989,
  -49.5199,
  -49.5403,
  -49.5597,
  -49.5778,
  -49.5944,
  -49.6098,
  -49.6242,
  -49.6375,
  -49.6505,
  -49.6636,
  -49.6772,
  -49.6905,
  -49.7054,
  -49.7207,
  -49.7362,
  -49.7518,
  -49.7676,
  -49.7838,
  -49.8003,
  -49.8166,
  -49.8324,
  -49.8472,
  -49.8609,
  -49.8736,
  -49.8857,
  -49.8975,
  -49.9091,
  -49.921,
  -49.9331,
  -49.9454,
  -49.9577,
  -49.9694,
  -49.9805,
  -49.9906,
  -49.9999,
  -50.0085,
  -50.017,
  -50.0243,
  -50.0326,
  -50.0403,
  -50.0468,
  -50.0516,
  -50.0544,
  -50.0554,
  -50.0546,
  -50.0523,
  -50.0488,
  -50.0443,
  -50.0393,
  -50.0345,
  -50.0305,
  -50.0279,
  -50.0267,
  -50.0266,
  -50.0271,
  -50.0277,
  -50.0282,
  -50.0289,
  -50.0299,
  -50.0311,
  -50.0324,
  -50.0331,
  -50.0328,
  -50.0313,
  -50.0287,
  -50.025,
  -50.0204,
  -50.014,
  -50.0079,
  -50.001,
  -49.9933,
  -49.9849,
  -49.9757,
  -49.9656,
  -49.9547,
  -49.9429,
  -49.93,
  -49.9157,
  -49.9002,
  -49.8832,
  -49.865,
  -49.8457,
  -49.8257,
  -49.8056,
  -49.7857,
  -49.7662,
  -49.7472,
  -49.7284,
  -49.7099,
  -49.6913,
  -49.6722,
  -49.6525,
  -49.6324,
  -49.6121,
  -49.5918,
  -49.5716,
  -49.5512,
  -49.531,
  -49.511,
  -49.4917,
  -49.4732,
  -49.4557,
  -49.4392,
  -49.4221,
  -49.4063,
  -49.3904,
  -49.3748,
  -49.3595,
  -49.3451,
  -49.3314,
  -49.3184,
  -49.306,
  -49.2939,
  -49.2823,
  -49.271,
  -49.2598,
  -49.2488,
  -49.238,
  -49.2276,
  -49.2176,
  -49.2077,
  -49.198,
  -49.1884,
  -49.179,
  -49.1701,
  -49.1616,
  -49.1536,
  -49.1463,
  -49.1394,
  -49.1333,
  -49.1271,
  -49.1206,
  -49.114,
  -49.1069,
  -49.0992,
  -49.0912,
  -49.0827,
  -49.0736,
  -49.064,
  -49.0544,
  -49.0447,
  -49.0349,
  -48.7783,
  -48.7972,
  -48.8158,
  -48.8328,
  -48.8485,
  -48.8619,
  -48.873,
  -48.8819,
  -48.8889,
  -48.8943,
  -48.8983,
  -48.9016,
  -48.9045,
  -48.9056,
  -48.9068,
  -48.9073,
  -48.9073,
  -48.9072,
  -48.9072,
  -48.9077,
  -48.9081,
  -48.9083,
  -48.9079,
  -48.907,
  -48.9052,
  -48.9024,
  -48.8985,
  -48.8935,
  -48.8867,
  -48.8807,
  -48.8751,
  -48.8707,
  -48.8685,
  -48.8691,
  -48.873,
  -48.8798,
  -48.8893,
  -48.9006,
  -48.9127,
  -48.9256,
  -48.9391,
  -48.9533,
  -48.9685,
  -48.9843,
  -48.9994,
  -49.0152,
  -49.0298,
  -49.0425,
  -49.053,
  -49.0612,
  -49.0675,
  -49.0725,
  -49.0766,
  -49.0805,
  -49.0851,
  -49.0907,
  -49.0975,
  -49.1055,
  -49.1143,
  -49.1234,
  -49.1319,
  -49.138,
  -49.1432,
  -49.1464,
  -49.1473,
  -49.146,
  -49.1422,
  -49.1359,
  -49.1275,
  -49.1172,
  -49.1053,
  -49.0918,
  -49.0767,
  -49.0602,
  -49.0432,
  -49.0261,
  -49.0093,
  -48.9931,
  -48.978,
  -48.9633,
  -48.9512,
  -48.9406,
  -48.9318,
  -48.9241,
  -48.9175,
  -48.9119,
  -48.9077,
  -48.9047,
  -48.9024,
  -48.9006,
  -48.8988,
  -48.8963,
  -48.8927,
  -48.8878,
  -48.8821,
  -48.8758,
  -48.8699,
  -48.8638,
  -48.8598,
  -48.8569,
  -48.8551,
  -48.8543,
  -48.854,
  -48.8543,
  -48.8549,
  -48.8555,
  -48.8564,
  -48.8575,
  -48.859,
  -48.8607,
  -48.8622,
  -48.8634,
  -48.8643,
  -48.8645,
  -48.8644,
  -48.8641,
  -48.8641,
  -48.864,
  -48.8663,
  -48.8707,
  -48.8772,
  -48.886,
  -48.8967,
  -48.9089,
  -48.9221,
  -48.9361,
  -48.951,
  -48.9672,
  -48.9849,
  -49.0046,
  -49.0265,
  -49.05,
  -49.0748,
  -49.1002,
  -49.1254,
  -49.1496,
  -49.1722,
  -49.193,
  -49.211,
  -49.2284,
  -49.2441,
  -49.2587,
  -49.2727,
  -49.2864,
  -49.3004,
  -49.3145,
  -49.3291,
  -49.3441,
  -49.3592,
  -49.3748,
  -49.3909,
  -49.4076,
  -49.4253,
  -49.4441,
  -49.4641,
  -49.4851,
  -49.5068,
  -49.5288,
  -49.5508,
  -49.5725,
  -49.5933,
  -49.6117,
  -49.6294,
  -49.6453,
  -49.6597,
  -49.6729,
  -49.6854,
  -49.6976,
  -49.7102,
  -49.7235,
  -49.7378,
  -49.7531,
  -49.7691,
  -49.7857,
  -49.8026,
  -49.8201,
  -49.8378,
  -49.8556,
  -49.8731,
  -49.8897,
  -49.905,
  -49.9188,
  -49.9313,
  -49.9431,
  -49.9544,
  -49.966,
  -49.9769,
  -49.9892,
  -50.0019,
  -50.0145,
  -50.027,
  -50.0387,
  -50.0495,
  -50.0594,
  -50.0686,
  -50.0774,
  -50.0859,
  -50.0942,
  -50.1018,
  -50.1083,
  -50.1129,
  -50.1154,
  -50.116,
  -50.1151,
  -50.1127,
  -50.1092,
  -50.1047,
  -50.0995,
  -50.0944,
  -50.09,
  -50.0867,
  -50.0846,
  -50.0834,
  -50.0824,
  -50.0802,
  -50.0788,
  -50.0774,
  -50.0766,
  -50.0762,
  -50.0762,
  -50.076,
  -50.0752,
  -50.0735,
  -50.0709,
  -50.0674,
  -50.0629,
  -50.0573,
  -50.0508,
  -50.0433,
  -50.0348,
  -50.0253,
  -50.0151,
  -50.0041,
  -49.9924,
  -49.9798,
  -49.9665,
  -49.9519,
  -49.9365,
  -49.9198,
  -49.9024,
  -49.8841,
  -49.8652,
  -49.8461,
  -49.8269,
  -49.8078,
  -49.7888,
  -49.7698,
  -49.7507,
  -49.7302,
  -49.7107,
  -49.6906,
  -49.6702,
  -49.6497,
  -49.6292,
  -49.6084,
  -49.5874,
  -49.5665,
  -49.5459,
  -49.5259,
  -49.5068,
  -49.4886,
  -49.4714,
  -49.4546,
  -49.4381,
  -49.4216,
  -49.4054,
  -49.3894,
  -49.3742,
  -49.3599,
  -49.3461,
  -49.3328,
  -49.3198,
  -49.3069,
  -49.2942,
  -49.2817,
  -49.2694,
  -49.2577,
  -49.2466,
  -49.236,
  -49.2259,
  -49.216,
  -49.2063,
  -49.1967,
  -49.1876,
  -49.1788,
  -49.1704,
  -49.1624,
  -49.1552,
  -49.1485,
  -49.142,
  -49.1359,
  -49.1283,
  -49.1215,
  -49.1141,
  -49.1062,
  -49.0977,
  -49.089,
  -49.08,
  -49.0709,
  -49.0618,
  -49.0528,
  -48.7724,
  -48.794,
  -48.8148,
  -48.834,
  -48.8511,
  -48.8663,
  -48.879,
  -48.8894,
  -48.8971,
  -48.9039,
  -48.9093,
  -48.9135,
  -48.9169,
  -48.9196,
  -48.9211,
  -48.9216,
  -48.9221,
  -48.9224,
  -48.9229,
  -48.9233,
  -48.9237,
  -48.9238,
  -48.9238,
  -48.9224,
  -48.9214,
  -48.9196,
  -48.9167,
  -48.9125,
  -48.9074,
  -48.9018,
  -48.8963,
  -48.8918,
  -48.8891,
  -48.8888,
  -48.8916,
  -48.8972,
  -48.9054,
  -48.9154,
  -48.9257,
  -48.938,
  -48.9511,
  -48.9652,
  -48.9806,
  -48.9969,
  -49.0137,
  -49.0304,
  -49.0458,
  -49.0591,
  -49.0699,
  -49.0783,
  -49.0846,
  -49.0894,
  -49.0932,
  -49.0967,
  -49.1005,
  -49.1044,
  -49.1104,
  -49.1176,
  -49.1258,
  -49.1346,
  -49.1433,
  -49.1512,
  -49.1577,
  -49.1625,
  -49.1654,
  -49.1661,
  -49.1643,
  -49.16,
  -49.1534,
  -49.1448,
  -49.1345,
  -49.1228,
  -49.1086,
  -49.094,
  -49.0788,
  -49.0635,
  -49.0484,
  -49.0337,
  -49.0194,
  -49.0066,
  -48.995,
  -48.9847,
  -48.9754,
  -48.9678,
  -48.9611,
  -48.9555,
  -48.9511,
  -48.9484,
  -48.9473,
  -48.9467,
  -48.9452,
  -48.9446,
  -48.9428,
  -48.9398,
  -48.9358,
  -48.9314,
  -48.9269,
  -48.9231,
  -48.9202,
  -48.9181,
  -48.9167,
  -48.9158,
  -48.9152,
  -48.9149,
  -48.9149,
  -48.9151,
  -48.9153,
  -48.9158,
  -48.9165,
  -48.9163,
  -48.9169,
  -48.9172,
  -48.9172,
  -48.9168,
  -48.916,
  -48.9152,
  -48.9148,
  -48.9152,
  -48.9171,
  -48.921,
  -48.927,
  -48.935,
  -48.9451,
  -48.957,
  -48.9701,
  -48.9842,
  -48.9993,
  -49.0157,
  -49.0336,
  -49.054,
  -49.0752,
  -49.0993,
  -49.1245,
  -49.1505,
  -49.1763,
  -49.201,
  -49.2241,
  -49.2452,
  -49.2645,
  -49.2821,
  -49.2983,
  -49.3134,
  -49.3275,
  -49.3411,
  -49.3545,
  -49.3682,
  -49.3821,
  -49.3962,
  -49.4108,
  -49.4259,
  -49.4417,
  -49.4584,
  -49.4753,
  -49.4947,
  -49.5157,
  -49.5379,
  -49.5608,
  -49.5837,
  -49.6064,
  -49.6285,
  -49.6493,
  -49.6684,
  -49.6854,
  -49.7004,
  -49.7137,
  -49.7259,
  -49.7375,
  -49.7492,
  -49.7614,
  -49.7747,
  -49.7891,
  -49.8047,
  -49.8214,
  -49.8391,
  -49.8574,
  -49.8763,
  -49.8945,
  -49.9137,
  -49.9322,
  -49.9497,
  -49.9654,
  -49.9793,
  -49.9916,
  -50.003,
  -50.0141,
  -50.0256,
  -50.0376,
  -50.0501,
  -50.0631,
  -50.0763,
  -50.0893,
  -50.1017,
  -50.1133,
  -50.1239,
  -50.1336,
  -50.1427,
  -50.1513,
  -50.1596,
  -50.1671,
  -50.1733,
  -50.1777,
  -50.1801,
  -50.1808,
  -50.179,
  -50.1769,
  -50.1736,
  -50.1692,
  -50.164,
  -50.1587,
  -50.1537,
  -50.1496,
  -50.1465,
  -50.1439,
  -50.1411,
  -50.1379,
  -50.1345,
  -50.1311,
  -50.1285,
  -50.1266,
  -50.1252,
  -50.124,
  -50.1226,
  -50.1206,
  -50.118,
  -50.1146,
  -50.1101,
  -50.1043,
  -50.097,
  -50.0884,
  -50.0785,
  -50.0676,
  -50.056,
  -50.0438,
  -50.0311,
  -50.0179,
  -50.0029,
  -49.9881,
  -49.9725,
  -49.9562,
  -49.9394,
  -49.9222,
  -49.9044,
  -49.8863,
  -49.8678,
  -49.8492,
  -49.8303,
  -49.8111,
  -49.7916,
  -49.7715,
  -49.7515,
  -49.7314,
  -49.7111,
  -49.6908,
  -49.6703,
  -49.6493,
  -49.628,
  -49.6065,
  -49.5854,
  -49.5649,
  -49.5451,
  -49.5263,
  -49.5086,
  -49.4911,
  -49.4741,
  -49.4566,
  -49.4395,
  -49.4229,
  -49.4066,
  -49.3911,
  -49.3762,
  -49.3616,
  -49.3471,
  -49.3329,
  -49.3179,
  -49.3041,
  -49.2908,
  -49.2781,
  -49.2662,
  -49.255,
  -49.2444,
  -49.2343,
  -49.2246,
  -49.215,
  -49.2057,
  -49.1966,
  -49.1876,
  -49.179,
  -49.1711,
  -49.1639,
  -49.1573,
  -49.1507,
  -49.1442,
  -49.1373,
  -49.1302,
  -49.1225,
  -49.1144,
  -49.106,
  -49.0974,
  -49.0889,
  -49.0806,
  -49.0724,
  -48.7638,
  -48.7889,
  -48.8115,
  -48.8331,
  -48.8524,
  -48.8692,
  -48.8835,
  -48.8957,
  -48.9058,
  -48.914,
  -48.9207,
  -48.926,
  -48.9302,
  -48.9335,
  -48.9355,
  -48.9365,
  -48.937,
  -48.9363,
  -48.9366,
  -48.9369,
  -48.9371,
  -48.9374,
  -48.9376,
  -48.9378,
  -48.9379,
  -48.9375,
  -48.9358,
  -48.9328,
  -48.9287,
  -48.9239,
  -48.9192,
  -48.915,
  -48.9122,
  -48.9105,
  -48.9125,
  -48.9171,
  -48.9241,
  -48.933,
  -48.9434,
  -48.9551,
  -48.9676,
  -48.9815,
  -48.9966,
  -49.0128,
  -49.0299,
  -49.0469,
  -49.0627,
  -49.0764,
  -49.0876,
  -49.0956,
  -49.1024,
  -49.1075,
  -49.1114,
  -49.1149,
  -49.1184,
  -49.1225,
  -49.1276,
  -49.1339,
  -49.1412,
  -49.1493,
  -49.1577,
  -49.1658,
  -49.1731,
  -49.179,
  -49.1832,
  -49.1854,
  -49.1844,
  -49.1818,
  -49.1768,
  -49.1698,
  -49.1612,
  -49.1512,
  -49.1402,
  -49.128,
  -49.1151,
  -49.102,
  -49.0888,
  -49.0757,
  -49.063,
  -49.0509,
  -49.0397,
  -49.0295,
  -49.0203,
  -49.0113,
  -49.0044,
  -48.9986,
  -48.9945,
  -48.992,
  -48.9913,
  -48.9918,
  -48.9929,
  -48.9937,
  -48.9939,
  -48.9928,
  -48.9907,
  -48.988,
  -48.985,
  -48.9824,
  -48.9806,
  -48.9793,
  -48.9782,
  -48.9775,
  -48.9757,
  -48.9753,
  -48.9751,
  -48.9752,
  -48.9754,
  -48.9756,
  -48.9759,
  -48.976,
  -48.976,
  -48.9758,
  -48.9753,
  -48.9746,
  -48.9736,
  -48.9726,
  -48.9719,
  -48.9721,
  -48.9733,
  -48.9763,
  -48.9812,
  -48.9882,
  -48.9962,
  -49.0072,
  -49.0198,
  -49.0337,
  -49.049,
  -49.0657,
  -49.0841,
  -49.1049,
  -49.1277,
  -49.1526,
  -49.1787,
  -49.2054,
  -49.2318,
  -49.2571,
  -49.2805,
  -49.302,
  -49.3217,
  -49.3396,
  -49.3562,
  -49.3718,
  -49.3863,
  -49.399,
  -49.4123,
  -49.4253,
  -49.4386,
  -49.452,
  -49.466,
  -49.4807,
  -49.4963,
  -49.5132,
  -49.5316,
  -49.5519,
  -49.5739,
  -49.5971,
  -49.6208,
  -49.6444,
  -49.6675,
  -49.6896,
  -49.7102,
  -49.7287,
  -49.7448,
  -49.7588,
  -49.7711,
  -49.7825,
  -49.7936,
  -49.8041,
  -49.8163,
  -49.8296,
  -49.8443,
  -49.8604,
  -49.8777,
  -49.8962,
  -49.9157,
  -49.9358,
  -49.9563,
  -49.9766,
  -49.9962,
  -50.0142,
  -50.0303,
  -50.0444,
  -50.0563,
  -50.0675,
  -50.0785,
  -50.0899,
  -50.102,
  -50.1148,
  -50.1281,
  -50.1417,
  -50.1553,
  -50.1685,
  -50.1809,
  -50.1913,
  -50.2016,
  -50.2109,
  -50.2195,
  -50.2275,
  -50.2346,
  -50.2406,
  -50.2449,
  -50.2475,
  -50.2483,
  -50.248,
  -50.2464,
  -50.2434,
  -50.2392,
  -50.2339,
  -50.2283,
  -50.2229,
  -50.2181,
  -50.2137,
  -50.2094,
  -50.2047,
  -50.1995,
  -50.1941,
  -50.189,
  -50.1847,
  -50.1813,
  -50.1787,
  -50.1764,
  -50.1743,
  -50.171,
  -50.1682,
  -50.1647,
  -50.16,
  -50.1537,
  -50.1456,
  -50.1353,
  -50.1236,
  -50.1109,
  -50.0976,
  -50.084,
  -50.0703,
  -50.0563,
  -50.0416,
  -50.0263,
  -50.0105,
  -49.9944,
  -49.9782,
  -49.9618,
  -49.9451,
  -49.9279,
  -49.9103,
  -49.8921,
  -49.8733,
  -49.8543,
  -49.8348,
  -49.8148,
  -49.7945,
  -49.7744,
  -49.7544,
  -49.7344,
  -49.714,
  -49.6931,
  -49.6715,
  -49.6497,
  -49.6281,
  -49.6059,
  -49.5855,
  -49.5661,
  -49.5476,
  -49.5296,
  -49.5117,
  -49.4941,
  -49.4761,
  -49.4584,
  -49.441,
  -49.4243,
  -49.4078,
  -49.3916,
  -49.3757,
  -49.3601,
  -49.3447,
  -49.3296,
  -49.3154,
  -49.3018,
  -49.2891,
  -49.2771,
  -49.266,
  -49.2555,
  -49.2455,
  -49.2359,
  -49.2265,
  -49.2172,
  -49.2077,
  -49.1985,
  -49.19,
  -49.1822,
  -49.175,
  -49.1683,
  -49.1616,
  -49.1548,
  -49.1478,
  -49.1403,
  -49.1325,
  -49.1245,
  -49.1163,
  -49.1082,
  -49.1002,
  -49.0924,
  -48.7508,
  -48.7803,
  -48.8075,
  -48.8321,
  -48.8539,
  -48.8726,
  -48.8886,
  -48.9024,
  -48.9141,
  -48.9236,
  -48.9314,
  -48.9376,
  -48.9418,
  -48.9456,
  -48.9482,
  -48.9494,
  -48.9499,
  -48.95,
  -48.95,
  -48.9499,
  -48.95,
  -48.9504,
  -48.9511,
  -48.9521,
  -48.9534,
  -48.9543,
  -48.9541,
  -48.9516,
  -48.949,
  -48.9455,
  -48.9417,
  -48.9383,
  -48.9359,
  -48.9352,
  -48.9367,
  -48.9406,
  -48.9468,
  -48.955,
  -48.9647,
  -48.9757,
  -48.9878,
  -49.0011,
  -49.0158,
  -49.0307,
  -49.0472,
  -49.0638,
  -49.0794,
  -49.0932,
  -49.1048,
  -49.1146,
  -49.1223,
  -49.1284,
  -49.133,
  -49.1369,
  -49.1405,
  -49.1443,
  -49.1487,
  -49.154,
  -49.1602,
  -49.1664,
  -49.1741,
  -49.1819,
  -49.1892,
  -49.1956,
  -49.2005,
  -49.2038,
  -49.2049,
  -49.2035,
  -49.1999,
  -49.1943,
  -49.1874,
  -49.1795,
  -49.1705,
  -49.161,
  -49.1507,
  -49.1401,
  -49.1292,
  -49.1171,
  -49.1061,
  -49.0952,
  -49.0848,
  -49.0749,
  -49.0659,
  -49.0576,
  -49.0505,
  -49.0446,
  -49.0404,
  -49.038,
  -49.0376,
  -49.0385,
  -49.041,
  -49.0433,
  -49.045,
  -49.0455,
  -49.0451,
  -49.043,
  -49.0416,
  -49.0403,
  -49.0392,
  -49.0386,
  -49.0382,
  -49.0378,
  -49.0375,
  -49.0373,
  -49.0374,
  -49.0378,
  -49.0383,
  -49.0385,
  -49.0386,
  -49.0385,
  -49.0382,
  -49.0378,
  -49.0374,
  -49.0368,
  -49.0349,
  -49.0338,
  -49.0329,
  -49.0327,
  -49.0335,
  -49.0352,
  -49.0387,
  -49.0442,
  -49.0519,
  -49.0617,
  -49.0735,
  -49.0872,
  -49.1027,
  -49.1199,
  -49.1391,
  -49.1607,
  -49.1845,
  -49.21,
  -49.237,
  -49.2644,
  -49.2915,
  -49.3164,
  -49.34,
  -49.3617,
  -49.3815,
  -49.3998,
  -49.4169,
  -49.433,
  -49.4479,
  -49.4618,
  -49.4749,
  -49.4876,
  -49.5003,
  -49.5132,
  -49.5267,
  -49.5412,
  -49.557,
  -49.5743,
  -49.5935,
  -49.6147,
  -49.6376,
  -49.6616,
  -49.6859,
  -49.7098,
  -49.7318,
  -49.7536,
  -49.7735,
  -49.7912,
  -49.8064,
  -49.8195,
  -49.831,
  -49.8419,
  -49.8529,
  -49.8645,
  -49.8771,
  -49.8909,
  -49.9063,
  -49.9227,
  -49.9406,
  -49.9597,
  -49.98,
  -50.0011,
  -50.0225,
  -50.0437,
  -50.0639,
  -50.0825,
  -50.0987,
  -50.1127,
  -50.1246,
  -50.1345,
  -50.1454,
  -50.157,
  -50.1693,
  -50.1824,
  -50.1961,
  -50.2102,
  -50.2244,
  -50.2383,
  -50.2515,
  -50.2635,
  -50.2743,
  -50.2837,
  -50.2922,
  -50.3,
  -50.3068,
  -50.3126,
  -50.3169,
  -50.3198,
  -50.3212,
  -50.3214,
  -50.3201,
  -50.3172,
  -50.313,
  -50.3077,
  -50.3019,
  -50.2959,
  -50.2903,
  -50.2835,
  -50.2773,
  -50.2706,
  -50.2635,
  -50.2563,
  -50.2496,
  -50.2437,
  -50.2393,
  -50.2358,
  -50.2326,
  -50.2297,
  -50.2268,
  -50.2235,
  -50.2196,
  -50.2143,
  -50.2072,
  -50.1978,
  -50.186,
  -50.1724,
  -50.1577,
  -50.1426,
  -50.1273,
  -50.1124,
  -50.0974,
  -50.0821,
  -50.0663,
  -50.0502,
  -50.0342,
  -50.0184,
  -50.0028,
  -49.9868,
  -49.9704,
  -49.9533,
  -49.9347,
  -49.9164,
  -49.8977,
  -49.8784,
  -49.8588,
  -49.8389,
  -49.8191,
  -49.7992,
  -49.7793,
  -49.759,
  -49.7381,
  -49.7164,
  -49.6943,
  -49.6721,
  -49.6504,
  -49.6295,
  -49.6095,
  -49.5903,
  -49.5716,
  -49.5533,
  -49.535,
  -49.5165,
  -49.4979,
  -49.4794,
  -49.4611,
  -49.4431,
  -49.4253,
  -49.4077,
  -49.3905,
  -49.3739,
  -49.3578,
  -49.3424,
  -49.328,
  -49.3145,
  -49.3019,
  -49.29,
  -49.2791,
  -49.2689,
  -49.2591,
  -49.2494,
  -49.2398,
  -49.229,
  -49.2193,
  -49.2103,
  -49.2019,
  -49.1942,
  -49.1872,
  -49.1805,
  -49.1735,
  -49.1665,
  -49.1592,
  -49.1517,
  -49.144,
  -49.1359,
  -49.1279,
  -49.1201,
  -49.1129,
  -48.7357,
  -48.7702,
  -48.8017,
  -48.8299,
  -48.8547,
  -48.8756,
  -48.8925,
  -48.9079,
  -48.921,
  -48.9319,
  -48.9407,
  -48.9479,
  -48.9539,
  -48.9584,
  -48.9611,
  -48.9626,
  -48.963,
  -48.9626,
  -48.962,
  -48.9616,
  -48.9615,
  -48.961,
  -48.9623,
  -48.9644,
  -48.967,
  -48.9691,
  -48.9705,
  -48.9708,
  -48.9698,
  -48.9679,
  -48.9654,
  -48.963,
  -48.9612,
  -48.9609,
  -48.9624,
  -48.9662,
  -48.9721,
  -48.9788,
  -48.9881,
  -48.9986,
  -49.0103,
  -49.0233,
  -49.0373,
  -49.0524,
  -49.068,
  -49.0834,
  -49.0983,
  -49.1119,
  -49.1241,
  -49.1348,
  -49.1437,
  -49.1509,
  -49.1567,
  -49.1605,
  -49.1646,
  -49.1685,
  -49.1726,
  -49.1771,
  -49.1824,
  -49.1884,
  -49.1953,
  -49.2023,
  -49.2091,
  -49.2152,
  -49.2201,
  -49.2236,
  -49.2252,
  -49.2246,
  -49.222,
  -49.2177,
  -49.2114,
  -49.2055,
  -49.1991,
  -49.1922,
  -49.1847,
  -49.1768,
  -49.1685,
  -49.16,
  -49.1512,
  -49.1422,
  -49.1326,
  -49.1233,
  -49.1144,
  -49.1063,
  -49.099,
  -49.0931,
  -49.0889,
  -49.0865,
  -49.0851,
  -49.0865,
  -49.0893,
  -49.0923,
  -49.0952,
  -49.0972,
  -49.0981,
  -49.0984,
  -49.0983,
  -49.098,
  -49.0979,
  -49.0981,
  -49.0985,
  -49.099,
  -49.0995,
  -49.1001,
  -49.1007,
  -49.1016,
  -49.1025,
  -49.1021,
  -49.1023,
  -49.1022,
  -49.1021,
  -49.102,
  -49.1019,
  -49.1016,
  -49.101,
  -49.1001,
  -49.0992,
  -49.0986,
  -49.0985,
  -49.0992,
  -49.1012,
  -49.1051,
  -49.1113,
  -49.1199,
  -49.131,
  -49.1445,
  -49.1602,
  -49.1771,
  -49.1973,
  -49.2199,
  -49.2447,
  -49.2712,
  -49.2988,
  -49.327,
  -49.3545,
  -49.3806,
  -49.4046,
  -49.4265,
  -49.4465,
  -49.4651,
  -49.4825,
  -49.4991,
  -49.5144,
  -49.5285,
  -49.5415,
  -49.5539,
  -49.5662,
  -49.579,
  -49.5923,
  -49.606,
  -49.6221,
  -49.6401,
  -49.6601,
  -49.6822,
  -49.7058,
  -49.7303,
  -49.7548,
  -49.7787,
  -49.8012,
  -49.8222,
  -49.8412,
  -49.8578,
  -49.8721,
  -49.8844,
  -49.8956,
  -49.9064,
  -49.9177,
  -49.9298,
  -49.9431,
  -49.9576,
  -49.9735,
  -49.9907,
  -50.0091,
  -50.0279,
  -50.0486,
  -50.0703,
  -50.0924,
  -50.1141,
  -50.1347,
  -50.1535,
  -50.1698,
  -50.1836,
  -50.1955,
  -50.2065,
  -50.2176,
  -50.2293,
  -50.242,
  -50.2554,
  -50.2696,
  -50.2841,
  -50.2989,
  -50.3134,
  -50.3273,
  -50.3398,
  -50.3509,
  -50.3604,
  -50.3687,
  -50.3761,
  -50.3828,
  -50.3884,
  -50.392,
  -50.3954,
  -50.3973,
  -50.3978,
  -50.3966,
  -50.3937,
  -50.3894,
  -50.3839,
  -50.3776,
  -50.3711,
  -50.3642,
  -50.357,
  -50.3492,
  -50.3407,
  -50.3318,
  -50.3231,
  -50.3153,
  -50.3085,
  -50.3031,
  -50.2986,
  -50.2947,
  -50.2909,
  -50.2871,
  -50.283,
  -50.2781,
  -50.2719,
  -50.2636,
  -50.2528,
  -50.2395,
  -50.2242,
  -50.2077,
  -50.1897,
  -50.1729,
  -50.1567,
  -50.1406,
  -50.1245,
  -50.1082,
  -50.0919,
  -50.0759,
  -50.0603,
  -50.0449,
  -50.0294,
  -50.0134,
  -49.997,
  -49.9797,
  -49.9618,
  -49.9435,
  -49.9248,
  -49.9057,
  -49.8864,
  -49.867,
  -49.8474,
  -49.8276,
  -49.807,
  -49.7858,
  -49.7638,
  -49.7413,
  -49.7187,
  -49.6967,
  -49.6753,
  -49.6549,
  -49.6352,
  -49.6161,
  -49.5973,
  -49.5784,
  -49.5594,
  -49.5401,
  -49.5206,
  -49.5009,
  -49.4802,
  -49.4608,
  -49.4415,
  -49.4228,
  -49.4049,
  -49.3879,
  -49.3715,
  -49.3562,
  -49.342,
  -49.3287,
  -49.3162,
  -49.3048,
  -49.2939,
  -49.2837,
  -49.2737,
  -49.2636,
  -49.2535,
  -49.2436,
  -49.2341,
  -49.2253,
  -49.2173,
  -49.2099,
  -49.203,
  -49.1962,
  -49.1888,
  -49.1815,
  -49.174,
  -49.1663,
  -49.1583,
  -49.1503,
  -49.1426,
  -49.1353,
  -48.7162,
  -48.7556,
  -48.7925,
  -48.8249,
  -48.8534,
  -48.8773,
  -48.8974,
  -48.9145,
  -48.9291,
  -48.9412,
  -48.951,
  -48.9591,
  -48.9654,
  -48.9702,
  -48.9735,
  -48.9749,
  -48.9742,
  -48.9734,
  -48.9723,
  -48.9715,
  -48.9713,
  -48.9723,
  -48.9742,
  -48.9771,
  -48.9809,
  -48.9842,
  -48.9871,
  -48.9891,
  -48.9898,
  -48.9896,
  -48.9887,
  -48.9864,
  -48.9856,
  -48.9859,
  -48.9879,
  -48.992,
  -48.998,
  -49.0057,
  -49.015,
  -49.0253,
  -49.0369,
  -49.0495,
  -49.0629,
  -49.077,
  -49.0913,
  -49.1056,
  -49.1193,
  -49.1313,
  -49.1439,
  -49.1552,
  -49.1651,
  -49.1737,
  -49.1809,
  -49.1869,
  -49.1921,
  -49.1967,
  -49.2009,
  -49.2051,
  -49.2096,
  -49.2147,
  -49.2205,
  -49.2264,
  -49.2323,
  -49.2374,
  -49.2407,
  -49.2436,
  -49.2449,
  -49.2446,
  -49.2426,
  -49.2394,
  -49.2357,
  -49.2317,
  -49.2277,
  -49.2235,
  -49.219,
  -49.2141,
  -49.2089,
  -49.2032,
  -49.1969,
  -49.19,
  -49.1821,
  -49.1725,
  -49.1642,
  -49.1564,
  -49.1495,
  -49.1438,
  -49.1396,
  -49.1372,
  -49.1368,
  -49.1381,
  -49.1408,
  -49.144,
  -49.1471,
  -49.1499,
  -49.152,
  -49.1534,
  -49.1544,
  -49.1552,
  -49.1561,
  -49.1572,
  -49.1576,
  -49.1593,
  -49.1609,
  -49.1626,
  -49.1642,
  -49.1657,
  -49.1671,
  -49.1682,
  -49.1688,
  -49.169,
  -49.1692,
  -49.1696,
  -49.1701,
  -49.1704,
  -49.1703,
  -49.1697,
  -49.1689,
  -49.1678,
  -49.167,
  -49.1667,
  -49.1665,
  -49.1691,
  -49.1739,
  -49.1815,
  -49.1921,
  -49.2054,
  -49.2216,
  -49.2403,
  -49.2615,
  -49.2851,
  -49.3107,
  -49.3381,
  -49.3664,
  -49.3949,
  -49.4227,
  -49.449,
  -49.4732,
  -49.4952,
  -49.5154,
  -49.5344,
  -49.5522,
  -49.5681,
  -49.5838,
  -49.5982,
  -49.6114,
  -49.6237,
  -49.6359,
  -49.6485,
  -49.6619,
  -49.6769,
  -49.6936,
  -49.7125,
  -49.7335,
  -49.7563,
  -49.7805,
  -49.8051,
  -49.8295,
  -49.8528,
  -49.8746,
  -49.8944,
  -49.9121,
  -49.9275,
  -49.941,
  -49.9529,
  -49.963,
  -49.9742,
  -49.9861,
  -49.9992,
  -50.0134,
  -50.0288,
  -50.0454,
  -50.0633,
  -50.0823,
  -50.1023,
  -50.1234,
  -50.1454,
  -50.1678,
  -50.1898,
  -50.2106,
  -50.2293,
  -50.2455,
  -50.2593,
  -50.2715,
  -50.2829,
  -50.2944,
  -50.3065,
  -50.3196,
  -50.3335,
  -50.3482,
  -50.3632,
  -50.3774,
  -50.3924,
  -50.4066,
  -50.4194,
  -50.4305,
  -50.44,
  -50.4481,
  -50.4553,
  -50.4618,
  -50.4675,
  -50.4724,
  -50.4761,
  -50.4784,
  -50.479,
  -50.4778,
  -50.4748,
  -50.4702,
  -50.4642,
  -50.4574,
  -50.4499,
  -50.4419,
  -50.4332,
  -50.4237,
  -50.4139,
  -50.4039,
  -50.3943,
  -50.3856,
  -50.378,
  -50.3716,
  -50.3653,
  -50.3605,
  -50.3559,
  -50.351,
  -50.3456,
  -50.3394,
  -50.3318,
  -50.3221,
  -50.3098,
  -50.2952,
  -50.2785,
  -50.2605,
  -50.2421,
  -50.2239,
  -50.2063,
  -50.1891,
  -50.1721,
  -50.1553,
  -50.1388,
  -50.1227,
  -50.1072,
  -50.0918,
  -50.0761,
  -50.0602,
  -50.0438,
  -50.0268,
  -50.0093,
  -49.9915,
  -49.9733,
  -49.9549,
  -49.9362,
  -49.917,
  -49.8973,
  -49.8772,
  -49.8564,
  -49.8337,
  -49.8113,
  -49.7884,
  -49.7658,
  -49.7435,
  -49.7219,
  -49.7012,
  -49.6811,
  -49.6614,
  -49.6421,
  -49.6229,
  -49.6034,
  -49.5835,
  -49.5632,
  -49.5423,
  -49.5214,
  -49.5005,
  -49.4798,
  -49.4597,
  -49.4404,
  -49.4221,
  -49.405,
  -49.3889,
  -49.3736,
  -49.3598,
  -49.3469,
  -49.3348,
  -49.3234,
  -49.3125,
  -49.3018,
  -49.2911,
  -49.2808,
  -49.2705,
  -49.2607,
  -49.2515,
  -49.2432,
  -49.2352,
  -49.2279,
  -49.2208,
  -49.2133,
  -49.2059,
  -49.1982,
  -49.1903,
  -49.1823,
  -49.1743,
  -49.1655,
  -49.1583,
  -48.694,
  -48.7403,
  -48.7825,
  -48.8204,
  -48.8528,
  -48.8799,
  -48.9025,
  -48.9215,
  -48.9374,
  -48.9506,
  -48.9604,
  -48.9691,
  -48.976,
  -48.9812,
  -48.9844,
  -48.986,
  -48.986,
  -48.985,
  -48.9834,
  -48.9827,
  -48.9825,
  -48.984,
  -48.9865,
  -48.9903,
  -48.9949,
  -48.9983,
  -49.0023,
  -49.0057,
  -49.0082,
  -49.0097,
  -49.0103,
  -49.0104,
  -49.0106,
  -49.0118,
  -49.0146,
  -49.0193,
  -49.026,
  -49.0342,
  -49.0437,
  -49.0542,
  -49.0658,
  -49.0771,
  -49.09,
  -49.1031,
  -49.1161,
  -49.1289,
  -49.1415,
  -49.154,
  -49.1663,
  -49.178,
  -49.1888,
  -49.1984,
  -49.2069,
  -49.2144,
  -49.2209,
  -49.2266,
  -49.2316,
  -49.2352,
  -49.2395,
  -49.244,
  -49.2487,
  -49.2533,
  -49.2578,
  -49.2617,
  -49.2646,
  -49.2665,
  -49.2669,
  -49.2663,
  -49.2646,
  -49.2623,
  -49.2598,
  -49.2576,
  -49.2558,
  -49.2543,
  -49.2528,
  -49.2501,
  -49.2481,
  -49.2457,
  -49.2423,
  -49.2375,
  -49.2313,
  -49.2241,
  -49.2166,
  -49.2096,
  -49.2035,
  -49.1985,
  -49.1948,
  -49.1926,
  -49.192,
  -49.1929,
  -49.1948,
  -49.1974,
  -49.2004,
  -49.2023,
  -49.2051,
  -49.2075,
  -49.2096,
  -49.2114,
  -49.2133,
  -49.2155,
  -49.2182,
  -49.2212,
  -49.2242,
  -49.2271,
  -49.2298,
  -49.2321,
  -49.2341,
  -49.2357,
  -49.2367,
  -49.2374,
  -49.2383,
  -49.2393,
  -49.2396,
  -49.2407,
  -49.2412,
  -49.241,
  -49.2402,
  -49.239,
  -49.2377,
  -49.2367,
  -49.2366,
  -49.2383,
  -49.2422,
  -49.2492,
  -49.2593,
  -49.2727,
  -49.2895,
  -49.3089,
  -49.3311,
  -49.3556,
  -49.382,
  -49.4098,
  -49.4384,
  -49.466,
  -49.4938,
  -49.5201,
  -49.5444,
  -49.5667,
  -49.5874,
  -49.6066,
  -49.6249,
  -49.6422,
  -49.6584,
  -49.6731,
  -49.6866,
  -49.6992,
  -49.7113,
  -49.7239,
  -49.7376,
  -49.7531,
  -49.7708,
  -49.7906,
  -49.8125,
  -49.836,
  -49.8603,
  -49.8838,
  -49.9076,
  -49.9301,
  -49.9506,
  -49.9691,
  -49.9854,
  -49.9998,
  -50.0126,
  -50.0243,
  -50.0359,
  -50.0478,
  -50.0607,
  -50.0749,
  -50.0901,
  -50.1065,
  -50.124,
  -50.1424,
  -50.1617,
  -50.1821,
  -50.2034,
  -50.2256,
  -50.248,
  -50.2701,
  -50.2907,
  -50.3091,
  -50.3241,
  -50.3381,
  -50.3506,
  -50.3626,
  -50.3747,
  -50.3875,
  -50.4011,
  -50.4155,
  -50.4308,
  -50.4464,
  -50.4621,
  -50.4771,
  -50.4913,
  -50.504,
  -50.515,
  -50.5243,
  -50.5323,
  -50.5394,
  -50.5458,
  -50.5517,
  -50.5568,
  -50.5609,
  -50.5632,
  -50.5637,
  -50.5622,
  -50.5589,
  -50.554,
  -50.5477,
  -50.5392,
  -50.5306,
  -50.5213,
  -50.5113,
  -50.5008,
  -50.4899,
  -50.4792,
  -50.4689,
  -50.4594,
  -50.4509,
  -50.4437,
  -50.4375,
  -50.4318,
  -50.4262,
  -50.4202,
  -50.4134,
  -50.4057,
  -50.3965,
  -50.3852,
  -50.3718,
  -50.3557,
  -50.3379,
  -50.319,
  -50.2996,
  -50.2803,
  -50.2612,
  -50.2428,
  -50.225,
  -50.2078,
  -50.1909,
  -50.1745,
  -50.1586,
  -50.1416,
  -50.1255,
  -50.1092,
  -50.0926,
  -50.0757,
  -50.0584,
  -50.0408,
  -50.0233,
  -50.0053,
  -49.9866,
  -49.9677,
  -49.9479,
  -49.9274,
  -49.9059,
  -49.8836,
  -49.8606,
  -49.8376,
  -49.8148,
  -49.7927,
  -49.7712,
  -49.7502,
  -49.7298,
  -49.7096,
  -49.6899,
  -49.6704,
  -49.6505,
  -49.6301,
  -49.6091,
  -49.5875,
  -49.5655,
  -49.5435,
  -49.5216,
  -49.5003,
  -49.4797,
  -49.4601,
  -49.4418,
  -49.4247,
  -49.4091,
  -49.3947,
  -49.3813,
  -49.3677,
  -49.3556,
  -49.3439,
  -49.3324,
  -49.3212,
  -49.3101,
  -49.2994,
  -49.2891,
  -49.2794,
  -49.2704,
  -49.2621,
  -49.2544,
  -49.2467,
  -49.2389,
  -49.231,
  -49.223,
  -49.2148,
  -49.2066,
  -49.1985,
  -49.1907,
  -49.1833,
  -48.6722,
  -48.7242,
  -48.7722,
  -48.815,
  -48.8519,
  -48.8817,
  -48.907,
  -48.9281,
  -48.9454,
  -48.96,
  -48.9716,
  -48.9808,
  -48.9879,
  -48.9933,
  -48.9966,
  -48.9979,
  -48.9976,
  -48.9964,
  -48.995,
  -48.9942,
  -48.9934,
  -48.995,
  -48.9984,
  -49.0031,
  -49.0084,
  -49.0136,
  -49.0187,
  -49.0234,
  -49.0273,
  -49.0302,
  -49.0322,
  -49.0337,
  -49.0352,
  -49.0375,
  -49.0414,
  -49.0462,
  -49.0538,
  -49.0628,
  -49.0728,
  -49.0836,
  -49.0952,
  -49.1073,
  -49.1197,
  -49.1319,
  -49.1438,
  -49.1554,
  -49.167,
  -49.1787,
  -49.1905,
  -49.2022,
  -49.2134,
  -49.2228,
  -49.2324,
  -49.2412,
  -49.2493,
  -49.2565,
  -49.263,
  -49.2685,
  -49.2734,
  -49.2777,
  -49.2817,
  -49.2853,
  -49.2884,
  -49.2907,
  -49.2919,
  -49.2921,
  -49.2914,
  -49.29,
  -49.2871,
  -49.2852,
  -49.2837,
  -49.2829,
  -49.2831,
  -49.284,
  -49.2853,
  -49.2866,
  -49.2877,
  -49.2884,
  -49.2876,
  -49.2851,
  -49.2809,
  -49.2754,
  -49.2695,
  -49.2638,
  -49.259,
  -49.2552,
  -49.2515,
  -49.25,
  -49.2491,
  -49.2495,
  -49.2506,
  -49.2523,
  -49.2547,
  -49.2574,
  -49.2604,
  -49.2635,
  -49.2665,
  -49.2694,
  -49.2724,
  -49.2758,
  -49.2797,
  -49.284,
  -49.2884,
  -49.2926,
  -49.2963,
  -49.2986,
  -49.3013,
  -49.3035,
  -49.3052,
  -49.3067,
  -49.3082,
  -49.31,
  -49.3121,
  -49.3139,
  -49.3152,
  -49.3156,
  -49.3153,
  -49.3143,
  -49.3128,
  -49.3115,
  -49.3113,
  -49.3126,
  -49.3161,
  -49.3226,
  -49.3325,
  -49.3452,
  -49.3622,
  -49.3823,
  -49.4052,
  -49.4304,
  -49.4572,
  -49.4853,
  -49.5139,
  -49.5423,
  -49.5699,
  -49.596,
  -49.6204,
  -49.6429,
  -49.664,
  -49.6839,
  -49.7029,
  -49.7208,
  -49.7374,
  -49.7527,
  -49.7666,
  -49.7795,
  -49.792,
  -49.8039,
  -49.8181,
  -49.8342,
  -49.8525,
  -49.873,
  -49.8956,
  -49.9192,
  -49.9435,
  -49.9678,
  -49.9907,
  -50.0121,
  -50.0315,
  -50.0488,
  -50.0641,
  -50.0777,
  -50.09,
  -50.1018,
  -50.1138,
  -50.1265,
  -50.1405,
  -50.1557,
  -50.1722,
  -50.1897,
  -50.208,
  -50.2261,
  -50.2458,
  -50.2665,
  -50.2879,
  -50.3101,
  -50.3324,
  -50.3542,
  -50.3744,
  -50.3925,
  -50.4085,
  -50.4226,
  -50.4355,
  -50.448,
  -50.4607,
  -50.4741,
  -50.4883,
  -50.5033,
  -50.5192,
  -50.5353,
  -50.5511,
  -50.5662,
  -50.5801,
  -50.5925,
  -50.6032,
  -50.6123,
  -50.6201,
  -50.6261,
  -50.6325,
  -50.6386,
  -50.644,
  -50.648,
  -50.6502,
  -50.6505,
  -50.6487,
  -50.645,
  -50.6397,
  -50.6329,
  -50.6247,
  -50.6153,
  -50.6049,
  -50.5939,
  -50.5825,
  -50.5711,
  -50.5599,
  -50.549,
  -50.5388,
  -50.5296,
  -50.5213,
  -50.514,
  -50.5075,
  -50.5008,
  -50.4936,
  -50.4855,
  -50.4762,
  -50.4655,
  -50.4529,
  -50.4371,
  -50.4201,
  -50.4017,
  -50.3821,
  -50.3619,
  -50.3416,
  -50.3215,
  -50.302,
  -50.2833,
  -50.2652,
  -50.2477,
  -50.2306,
  -50.2138,
  -50.197,
  -50.18,
  -50.163,
  -50.1459,
  -50.1286,
  -50.1112,
  -50.0938,
  -50.0761,
  -50.0581,
  -50.0396,
  -50.0204,
  -50.0003,
  -49.9792,
  -49.9572,
  -49.9344,
  -49.9111,
  -49.888,
  -49.8653,
  -49.8433,
  -49.822,
  -49.8011,
  -49.7804,
  -49.76,
  -49.7398,
  -49.719,
  -49.6988,
  -49.678,
  -49.6565,
  -49.6343,
  -49.6117,
  -49.5888,
  -49.566,
  -49.5435,
  -49.5218,
  -49.5011,
  -49.4817,
  -49.4638,
  -49.4476,
  -49.4328,
  -49.419,
  -49.4061,
  -49.3935,
  -49.3811,
  -49.3688,
  -49.3566,
  -49.3446,
  -49.333,
  -49.3219,
  -49.3113,
  -49.3016,
  -49.2926,
  -49.2841,
  -49.2758,
  -49.2674,
  -49.2589,
  -49.2501,
  -49.2415,
  -49.233,
  -49.2247,
  -49.2167,
  -49.2092,
  -48.6512,
  -48.7084,
  -48.7618,
  -48.8094,
  -48.8505,
  -48.8849,
  -48.9131,
  -48.9365,
  -48.9558,
  -48.9715,
  -48.984,
  -48.9938,
  -49.0012,
  -49.0064,
  -49.0085,
  -49.0096,
  -49.0092,
  -49.0079,
  -49.0066,
  -49.0058,
  -49.0064,
  -49.0087,
  -49.0126,
  -49.0179,
  -49.0237,
  -49.0297,
  -49.0356,
  -49.0412,
  -49.0462,
  -49.0493,
  -49.0527,
  -49.0555,
  -49.0583,
  -49.0619,
  -49.0671,
  -49.0742,
  -49.0829,
  -49.0928,
  -49.1035,
  -49.1148,
  -49.1265,
  -49.1386,
  -49.1506,
  -49.1622,
  -49.1733,
  -49.183,
  -49.1935,
  -49.2044,
  -49.2155,
  -49.2268,
  -49.238,
  -49.2488,
  -49.2592,
  -49.2691,
  -49.2786,
  -49.2876,
  -49.2959,
  -49.3031,
  -49.3092,
  -49.3141,
  -49.3179,
  -49.3206,
  -49.3214,
  -49.322,
  -49.3216,
  -49.3201,
  -49.3179,
  -49.3155,
  -49.3131,
  -49.3112,
  -49.3103,
  -49.3106,
  -49.3124,
  -49.3153,
  -49.319,
  -49.323,
  -49.3269,
  -49.3301,
  -49.332,
  -49.331,
  -49.3291,
  -49.3256,
  -49.3214,
  -49.3176,
  -49.3145,
  -49.3123,
  -49.3109,
  -49.3101,
  -49.3095,
  -49.3093,
  -49.3094,
  -49.3102,
  -49.3117,
  -49.3141,
  -49.3172,
  -49.3208,
  -49.3246,
  -49.3286,
  -49.3318,
  -49.3364,
  -49.3416,
  -49.3471,
  -49.3526,
  -49.3578,
  -49.3626,
  -49.3668,
  -49.3704,
  -49.3735,
  -49.376,
  -49.3783,
  -49.3807,
  -49.3834,
  -49.3862,
  -49.389,
  -49.3912,
  -49.3925,
  -49.3929,
  -49.3924,
  -49.3905,
  -49.3896,
  -49.3895,
  -49.3908,
  -49.3944,
  -49.401,
  -49.411,
  -49.4246,
  -49.4419,
  -49.4625,
  -49.486,
  -49.5116,
  -49.5387,
  -49.5667,
  -49.5949,
  -49.6228,
  -49.6497,
  -49.6754,
  -49.6996,
  -49.7224,
  -49.7441,
  -49.7637,
  -49.7835,
  -49.8021,
  -49.8194,
  -49.8352,
  -49.8497,
  -49.8632,
  -49.8763,
  -49.8898,
  -49.9045,
  -49.9213,
  -49.9402,
  -49.9613,
  -49.9841,
  -50.0079,
  -50.032,
  -50.0556,
  -50.0778,
  -50.0982,
  -50.1166,
  -50.1329,
  -50.1474,
  -50.1605,
  -50.1718,
  -50.1838,
  -50.1962,
  -50.2097,
  -50.2247,
  -50.241,
  -50.2586,
  -50.2773,
  -50.2966,
  -50.3165,
  -50.3368,
  -50.3577,
  -50.3792,
  -50.4012,
  -50.4232,
  -50.4445,
  -50.4643,
  -50.482,
  -50.4977,
  -50.5119,
  -50.5251,
  -50.538,
  -50.5512,
  -50.5651,
  -50.5799,
  -50.5947,
  -50.611,
  -50.6274,
  -50.6434,
  -50.6583,
  -50.6719,
  -50.6837,
  -50.6939,
  -50.7026,
  -50.7103,
  -50.7172,
  -50.7237,
  -50.7299,
  -50.7352,
  -50.7392,
  -50.7412,
  -50.7411,
  -50.7389,
  -50.735,
  -50.7294,
  -50.7222,
  -50.7134,
  -50.7033,
  -50.6921,
  -50.6804,
  -50.6684,
  -50.6564,
  -50.6448,
  -50.6335,
  -50.6217,
  -50.6115,
  -50.6023,
  -50.594,
  -50.5863,
  -50.5786,
  -50.5703,
  -50.561,
  -50.5505,
  -50.5385,
  -50.5246,
  -50.5089,
  -50.4912,
  -50.4722,
  -50.4521,
  -50.4314,
  -50.4103,
  -50.3892,
  -50.3686,
  -50.3487,
  -50.3296,
  -50.3112,
  -50.2932,
  -50.2754,
  -50.2574,
  -50.2393,
  -50.2212,
  -50.2032,
  -50.1854,
  -50.1675,
  -50.1497,
  -50.1316,
  -50.1132,
  -50.0933,
  -50.0736,
  -50.0529,
  -50.0311,
  -50.0084,
  -49.985,
  -49.9614,
  -49.9383,
  -49.9158,
  -49.8942,
  -49.8731,
  -49.8524,
  -49.8317,
  -49.8111,
  -49.7907,
  -49.7705,
  -49.7502,
  -49.7292,
  -49.7075,
  -49.6849,
  -49.6618,
  -49.6383,
  -49.6149,
  -49.5916,
  -49.5689,
  -49.5471,
  -49.5267,
  -49.508,
  -49.4912,
  -49.4761,
  -49.4622,
  -49.4491,
  -49.4362,
  -49.4232,
  -49.4101,
  -49.3969,
  -49.3839,
  -49.3711,
  -49.3588,
  -49.3473,
  -49.3366,
  -49.3267,
  -49.3173,
  -49.3081,
  -49.2977,
  -49.2882,
  -49.2786,
  -49.2691,
  -49.2599,
  -49.2512,
  -49.2429,
  -49.2351,
  -48.6346,
  -48.6962,
  -48.7541,
  -48.8061,
  -48.8511,
  -48.8888,
  -48.9199,
  -48.9457,
  -48.9658,
  -48.9831,
  -48.9967,
  -49.0071,
  -49.0147,
  -49.0197,
  -49.0225,
  -49.0235,
  -49.0231,
  -49.022,
  -49.0208,
  -49.0203,
  -49.0212,
  -49.0238,
  -49.0283,
  -49.034,
  -49.0393,
  -49.0458,
  -49.0521,
  -49.0582,
  -49.0639,
  -49.069,
  -49.0736,
  -49.0777,
  -49.0819,
  -49.087,
  -49.0936,
  -49.1019,
  -49.1118,
  -49.1228,
  -49.1344,
  -49.1453,
  -49.1574,
  -49.1695,
  -49.1813,
  -49.1926,
  -49.2033,
  -49.2133,
  -49.2231,
  -49.233,
  -49.2434,
  -49.254,
  -49.2649,
  -49.2757,
  -49.2865,
  -49.2973,
  -49.308,
  -49.3187,
  -49.328,
  -49.3373,
  -49.3451,
  -49.3512,
  -49.3554,
  -49.3579,
  -49.3587,
  -49.358,
  -49.356,
  -49.3529,
  -49.3491,
  -49.3454,
  -49.3422,
  -49.3401,
  -49.3395,
  -49.3405,
  -49.3434,
  -49.3468,
  -49.3524,
  -49.3585,
  -49.3646,
  -49.3701,
  -49.3744,
  -49.3768,
  -49.3772,
  -49.376,
  -49.3741,
  -49.3724,
  -49.3713,
  -49.371,
  -49.3711,
  -49.3712,
  -49.371,
  -49.3705,
  -49.37,
  -49.3689,
  -49.3697,
  -49.3717,
  -49.3748,
  -49.3788,
  -49.3835,
  -49.3886,
  -49.394,
  -49.3999,
  -49.4061,
  -49.4125,
  -49.4188,
  -49.4249,
  -49.4305,
  -49.4356,
  -49.4402,
  -49.4441,
  -49.4477,
  -49.4509,
  -49.4533,
  -49.4568,
  -49.4606,
  -49.4644,
  -49.4678,
  -49.4704,
  -49.472,
  -49.4726,
  -49.4726,
  -49.4726,
  -49.4732,
  -49.4753,
  -49.4795,
  -49.4864,
  -49.4966,
  -49.5104,
  -49.5278,
  -49.5487,
  -49.5724,
  -49.5983,
  -49.6255,
  -49.6521,
  -49.6797,
  -49.7066,
  -49.7326,
  -49.7575,
  -49.7814,
  -49.8043,
  -49.8264,
  -49.8478,
  -49.8683,
  -49.8877,
  -49.9057,
  -49.9222,
  -49.9374,
  -49.9517,
  -49.9656,
  -49.9799,
  -49.9955,
  -50.0129,
  -50.0324,
  -50.0538,
  -50.0768,
  -50.0996,
  -50.1234,
  -50.1464,
  -50.1679,
  -50.1875,
  -50.2052,
  -50.2209,
  -50.2351,
  -50.2481,
  -50.2604,
  -50.2727,
  -50.2856,
  -50.2998,
  -50.3155,
  -50.3328,
  -50.3515,
  -50.3713,
  -50.3917,
  -50.4125,
  -50.4336,
  -50.4549,
  -50.4764,
  -50.4982,
  -50.5198,
  -50.5395,
  -50.5586,
  -50.5758,
  -50.5912,
  -50.6053,
  -50.6186,
  -50.6318,
  -50.6452,
  -50.6595,
  -50.6747,
  -50.6909,
  -50.7077,
  -50.7243,
  -50.7403,
  -50.755,
  -50.7681,
  -50.7794,
  -50.789,
  -50.7973,
  -50.8047,
  -50.8115,
  -50.8181,
  -50.8243,
  -50.8296,
  -50.8334,
  -50.8352,
  -50.8347,
  -50.8312,
  -50.8271,
  -50.8214,
  -50.814,
  -50.8048,
  -50.7941,
  -50.7823,
  -50.77,
  -50.7575,
  -50.7451,
  -50.7331,
  -50.7213,
  -50.7099,
  -50.699,
  -50.6888,
  -50.6795,
  -50.6707,
  -50.6621,
  -50.6528,
  -50.6426,
  -50.631,
  -50.6179,
  -50.6031,
  -50.5866,
  -50.5684,
  -50.5489,
  -50.5283,
  -50.507,
  -50.4852,
  -50.4632,
  -50.4415,
  -50.4205,
  -50.3993,
  -50.3798,
  -50.3606,
  -50.3415,
  -50.3222,
  -50.3027,
  -50.2834,
  -50.2642,
  -50.2454,
  -50.2268,
  -50.208,
  -50.1891,
  -50.1698,
  -50.15,
  -50.1294,
  -50.1078,
  -50.0852,
  -50.0617,
  -50.0378,
  -50.0139,
  -49.9908,
  -49.9685,
  -49.9472,
  -49.9265,
  -49.9059,
  -49.8854,
  -49.8648,
  -49.8445,
  -49.8242,
  -49.8038,
  -49.7828,
  -49.7608,
  -49.7381,
  -49.7148,
  -49.6912,
  -49.6674,
  -49.6435,
  -49.62,
  -49.5973,
  -49.575,
  -49.5557,
  -49.5383,
  -49.5229,
  -49.5089,
  -49.4956,
  -49.4825,
  -49.4692,
  -49.4554,
  -49.4413,
  -49.4271,
  -49.4131,
  -49.3996,
  -49.387,
  -49.3752,
  -49.3642,
  -49.3537,
  -49.3432,
  -49.3326,
  -49.3218,
  -49.3109,
  -49.3003,
  -49.2902,
  -49.2807,
  -49.2718,
  -49.2637,
  -48.6228,
  -48.6873,
  -48.7484,
  -48.8027,
  -48.8511,
  -48.892,
  -48.926,
  -48.9541,
  -48.9776,
  -48.9964,
  -49.0112,
  -49.0222,
  -49.0301,
  -49.0352,
  -49.038,
  -49.0389,
  -49.0385,
  -49.0375,
  -49.0355,
  -49.0352,
  -49.0364,
  -49.0394,
  -49.0442,
  -49.0503,
  -49.0568,
  -49.0635,
  -49.07,
  -49.0763,
  -49.0826,
  -49.0885,
  -49.0941,
  -49.0995,
  -49.1052,
  -49.1107,
  -49.1187,
  -49.1284,
  -49.1396,
  -49.1518,
  -49.1644,
  -49.1771,
  -49.1896,
  -49.2021,
  -49.214,
  -49.2252,
  -49.2356,
  -49.2453,
  -49.2546,
  -49.2638,
  -49.2734,
  -49.2823,
  -49.2926,
  -49.3031,
  -49.3139,
  -49.3252,
  -49.337,
  -49.3491,
  -49.3613,
  -49.3728,
  -49.3828,
  -49.3905,
  -49.3957,
  -49.3986,
  -49.3991,
  -49.3975,
  -49.3944,
  -49.3897,
  -49.3834,
  -49.3783,
  -49.3742,
  -49.3717,
  -49.371,
  -49.3723,
  -49.3758,
  -49.3812,
  -49.3881,
  -49.3958,
  -49.4036,
  -49.4109,
  -49.4172,
  -49.4219,
  -49.4247,
  -49.426,
  -49.4264,
  -49.4269,
  -49.4269,
  -49.4284,
  -49.43,
  -49.4312,
  -49.4318,
  -49.4316,
  -49.4311,
  -49.4307,
  -49.431,
  -49.4328,
  -49.4359,
  -49.4403,
  -49.4458,
  -49.452,
  -49.4588,
  -49.4659,
  -49.473,
  -49.48,
  -49.4868,
  -49.4923,
  -49.4984,
  -49.5042,
  -49.5094,
  -49.5142,
  -49.5187,
  -49.5229,
  -49.5272,
  -49.5318,
  -49.5367,
  -49.542,
  -49.5469,
  -49.5512,
  -49.5546,
  -49.557,
  -49.5585,
  -49.5598,
  -49.5618,
  -49.5651,
  -49.5704,
  -49.577,
  -49.5876,
  -49.6016,
  -49.619,
  -49.6399,
  -49.6636,
  -49.6895,
  -49.7165,
  -49.7437,
  -49.7703,
  -49.796,
  -49.8209,
  -49.8449,
  -49.8682,
  -49.891,
  -49.9133,
  -49.9352,
  -49.9564,
  -49.9765,
  -49.9953,
  -50.0125,
  -50.0274,
  -50.0426,
  -50.0575,
  -50.0729,
  -50.0896,
  -50.1074,
  -50.1273,
  -50.149,
  -50.1721,
  -50.1959,
  -50.2194,
  -50.242,
  -50.2632,
  -50.2824,
  -50.2998,
  -50.3154,
  -50.3296,
  -50.3426,
  -50.3552,
  -50.3678,
  -50.3812,
  -50.3959,
  -50.4124,
  -50.4305,
  -50.4492,
  -50.4698,
  -50.4915,
  -50.5135,
  -50.5353,
  -50.5571,
  -50.5787,
  -50.6002,
  -50.6212,
  -50.6412,
  -50.6596,
  -50.6762,
  -50.6912,
  -50.7052,
  -50.7185,
  -50.7316,
  -50.7451,
  -50.7594,
  -50.7749,
  -50.791,
  -50.8079,
  -50.8249,
  -50.8407,
  -50.8551,
  -50.8676,
  -50.8782,
  -50.8862,
  -50.8941,
  -50.9013,
  -50.9081,
  -50.9146,
  -50.9208,
  -50.9262,
  -50.93,
  -50.9316,
  -50.9309,
  -50.9284,
  -50.9241,
  -50.9183,
  -50.9108,
  -50.9013,
  -50.8901,
  -50.8779,
  -50.8651,
  -50.8521,
  -50.8393,
  -50.8269,
  -50.8148,
  -50.8029,
  -50.7914,
  -50.7805,
  -50.7702,
  -50.7604,
  -50.7507,
  -50.7406,
  -50.7296,
  -50.716,
  -50.702,
  -50.6865,
  -50.6695,
  -50.6508,
  -50.6308,
  -50.6096,
  -50.5877,
  -50.5651,
  -50.5423,
  -50.5196,
  -50.4975,
  -50.4761,
  -50.4554,
  -50.4352,
  -50.4147,
  -50.3938,
  -50.3728,
  -50.3518,
  -50.3313,
  -50.3112,
  -50.2914,
  -50.2715,
  -50.2512,
  -50.2305,
  -50.2092,
  -50.1872,
  -50.1644,
  -50.1408,
  -50.1165,
  -50.0919,
  -50.0679,
  -50.0449,
  -50.0229,
  -50.0019,
  -49.9814,
  -49.9601,
  -49.9397,
  -49.9196,
  -49.8995,
  -49.8793,
  -49.8589,
  -49.8379,
  -49.8158,
  -49.793,
  -49.7697,
  -49.746,
  -49.7221,
  -49.6979,
  -49.6738,
  -49.6505,
  -49.6287,
  -49.6089,
  -49.591,
  -49.5751,
  -49.5608,
  -49.5474,
  -49.5341,
  -49.5204,
  -49.5061,
  -49.4911,
  -49.476,
  -49.4609,
  -49.4464,
  -49.4328,
  -49.4199,
  -49.4076,
  -49.3956,
  -49.3836,
  -49.3714,
  -49.3591,
  -49.3469,
  -49.3351,
  -49.3238,
  -49.3133,
  -49.3038,
  -49.2953,
  -48.615,
  -48.681,
  -48.7438,
  -48.8012,
  -48.8521,
  -48.8959,
  -48.9329,
  -48.9638,
  -48.9894,
  -49.0101,
  -49.0262,
  -49.0381,
  -49.0453,
  -49.0506,
  -49.0535,
  -49.0546,
  -49.0544,
  -49.0534,
  -49.0524,
  -49.0522,
  -49.0537,
  -49.057,
  -49.0621,
  -49.0685,
  -49.0752,
  -49.0819,
  -49.0884,
  -49.0948,
  -49.1004,
  -49.1069,
  -49.1137,
  -49.1204,
  -49.1274,
  -49.1353,
  -49.1446,
  -49.1557,
  -49.1682,
  -49.1816,
  -49.1955,
  -49.2093,
  -49.2227,
  -49.2356,
  -49.2478,
  -49.2581,
  -49.2685,
  -49.2779,
  -49.287,
  -49.2959,
  -49.3049,
  -49.314,
  -49.3235,
  -49.3334,
  -49.344,
  -49.3555,
  -49.368,
  -49.3814,
  -49.3953,
  -49.4087,
  -49.4207,
  -49.4303,
  -49.4361,
  -49.44,
  -49.441,
  -49.4392,
  -49.4352,
  -49.4295,
  -49.423,
  -49.4168,
  -49.4118,
  -49.4087,
  -49.4077,
  -49.4091,
  -49.4129,
  -49.4187,
  -49.4264,
  -49.4352,
  -49.444,
  -49.4517,
  -49.4596,
  -49.4661,
  -49.4711,
  -49.4748,
  -49.4775,
  -49.4802,
  -49.4831,
  -49.4862,
  -49.4893,
  -49.4918,
  -49.4936,
  -49.4944,
  -49.4946,
  -49.4947,
  -49.4952,
  -49.4972,
  -49.5004,
  -49.5053,
  -49.5106,
  -49.5179,
  -49.5261,
  -49.5343,
  -49.5422,
  -49.5495,
  -49.5564,
  -49.5628,
  -49.5689,
  -49.5749,
  -49.5805,
  -49.5859,
  -49.5908,
  -49.5958,
  -49.601,
  -49.6067,
  -49.6131,
  -49.62,
  -49.6272,
  -49.633,
  -49.6388,
  -49.6435,
  -49.6473,
  -49.6507,
  -49.6546,
  -49.6595,
  -49.6661,
  -49.6747,
  -49.6858,
  -49.7,
  -49.7174,
  -49.7382,
  -49.7617,
  -49.7874,
  -49.8139,
  -49.8403,
  -49.8659,
  -49.8905,
  -49.9142,
  -49.9372,
  -49.9588,
  -49.9814,
  -50.0038,
  -50.026,
  -50.0476,
  -50.068,
  -50.0873,
  -50.1051,
  -50.1217,
  -50.1378,
  -50.1539,
  -50.1704,
  -50.1878,
  -50.2064,
  -50.2267,
  -50.2485,
  -50.2718,
  -50.2957,
  -50.3194,
  -50.342,
  -50.3632,
  -50.3825,
  -50.3999,
  -50.4147,
  -50.4291,
  -50.4423,
  -50.4552,
  -50.4682,
  -50.4822,
  -50.4976,
  -50.5147,
  -50.5336,
  -50.5542,
  -50.5759,
  -50.5985,
  -50.6213,
  -50.6438,
  -50.6661,
  -50.6879,
  -50.7089,
  -50.7292,
  -50.7483,
  -50.7659,
  -50.782,
  -50.7968,
  -50.8107,
  -50.8241,
  -50.8371,
  -50.8494,
  -50.8636,
  -50.8789,
  -50.8951,
  -50.9117,
  -50.9282,
  -50.9438,
  -50.9576,
  -50.9695,
  -50.9796,
  -50.9881,
  -50.9956,
  -51.0025,
  -51.0091,
  -51.0155,
  -51.0218,
  -51.0273,
  -51.0313,
  -51.0332,
  -51.0328,
  -51.0302,
  -51.026,
  -51.0201,
  -51.0122,
  -51.0023,
  -50.9907,
  -50.9781,
  -50.9648,
  -50.9504,
  -50.9373,
  -50.9245,
  -50.9121,
  -50.9001,
  -50.8883,
  -50.8767,
  -50.8655,
  -50.8548,
  -50.844,
  -50.8329,
  -50.8208,
  -50.8075,
  -50.793,
  -50.7768,
  -50.7592,
  -50.74,
  -50.7194,
  -50.6976,
  -50.6748,
  -50.6513,
  -50.6276,
  -50.6042,
  -50.5812,
  -50.559,
  -50.5374,
  -50.5159,
  -50.494,
  -50.4715,
  -50.4486,
  -50.4258,
  -50.4036,
  -50.3819,
  -50.3596,
  -50.3381,
  -50.3162,
  -50.2936,
  -50.2703,
  -50.2465,
  -50.2221,
  -50.1975,
  -50.1724,
  -50.1475,
  -50.1233,
  -50.1003,
  -50.0786,
  -50.0579,
  -50.0377,
  -50.0178,
  -49.9978,
  -49.978,
  -49.9583,
  -49.9385,
  -49.9181,
  -49.8969,
  -49.8747,
  -49.8517,
  -49.8282,
  -49.8045,
  -49.7805,
  -49.7562,
  -49.732,
  -49.7085,
  -49.6864,
  -49.6661,
  -49.6477,
  -49.6314,
  -49.6166,
  -49.6027,
  -49.5891,
  -49.5749,
  -49.5599,
  -49.5444,
  -49.5287,
  -49.5129,
  -49.4968,
  -49.4823,
  -49.4683,
  -49.4548,
  -49.4412,
  -49.4274,
  -49.4135,
  -49.3997,
  -49.3862,
  -49.3732,
  -49.3609,
  -49.3494,
  -49.339,
  -49.3298,
  -48.6132,
  -48.6794,
  -48.7424,
  -48.8007,
  -48.8532,
  -48.8994,
  -48.9391,
  -48.9717,
  -48.9997,
  -49.0225,
  -49.0402,
  -49.0534,
  -49.0624,
  -49.0683,
  -49.0713,
  -49.0724,
  -49.0721,
  -49.0711,
  -49.07,
  -49.0702,
  -49.072,
  -49.0758,
  -49.0803,
  -49.0869,
  -49.0938,
  -49.1004,
  -49.1069,
  -49.1133,
  -49.12,
  -49.127,
  -49.1347,
  -49.1425,
  -49.1509,
  -49.1601,
  -49.1708,
  -49.1832,
  -49.1971,
  -49.2119,
  -49.226,
  -49.241,
  -49.2554,
  -49.2691,
  -49.2816,
  -49.2931,
  -49.3036,
  -49.3132,
  -49.3224,
  -49.3312,
  -49.3397,
  -49.3483,
  -49.357,
  -49.366,
  -49.3761,
  -49.3875,
  -49.3994,
  -49.4137,
  -49.4289,
  -49.444,
  -49.4578,
  -49.4693,
  -49.4779,
  -49.4832,
  -49.4852,
  -49.4842,
  -49.4802,
  -49.4742,
  -49.4671,
  -49.4603,
  -49.4548,
  -49.4513,
  -49.4501,
  -49.4504,
  -49.4542,
  -49.4603,
  -49.4683,
  -49.4775,
  -49.4871,
  -49.4966,
  -49.5054,
  -49.5131,
  -49.5196,
  -49.5249,
  -49.5295,
  -49.534,
  -49.5386,
  -49.5434,
  -49.5481,
  -49.5523,
  -49.5556,
  -49.557,
  -49.5586,
  -49.56,
  -49.5618,
  -49.5646,
  -49.5684,
  -49.574,
  -49.5811,
  -49.5896,
  -49.5989,
  -49.608,
  -49.6165,
  -49.6239,
  -49.6305,
  -49.6365,
  -49.6423,
  -49.6478,
  -49.6531,
  -49.6583,
  -49.6622,
  -49.6677,
  -49.6737,
  -49.6806,
  -49.6887,
  -49.6978,
  -49.7074,
  -49.7169,
  -49.7257,
  -49.7335,
  -49.7404,
  -49.7465,
  -49.7529,
  -49.7601,
  -49.7682,
  -49.7779,
  -49.7899,
  -49.8043,
  -49.8218,
  -49.8424,
  -49.8647,
  -49.8897,
  -49.9155,
  -49.941,
  -49.9656,
  -49.9893,
  -50.0119,
  -50.034,
  -50.056,
  -50.0782,
  -50.1003,
  -50.1224,
  -50.1441,
  -50.1647,
  -50.1842,
  -50.2024,
  -50.2197,
  -50.2365,
  -50.2535,
  -50.271,
  -50.2893,
  -50.3088,
  -50.3286,
  -50.351,
  -50.3748,
  -50.399,
  -50.4229,
  -50.446,
  -50.4675,
  -50.4872,
  -50.505,
  -50.5211,
  -50.5357,
  -50.5494,
  -50.5627,
  -50.5765,
  -50.5912,
  -50.6075,
  -50.6254,
  -50.6451,
  -50.6663,
  -50.6888,
  -50.7119,
  -50.7352,
  -50.7582,
  -50.7806,
  -50.8011,
  -50.8216,
  -50.8412,
  -50.8594,
  -50.8765,
  -50.8923,
  -50.9071,
  -50.9211,
  -50.9343,
  -50.9473,
  -50.9605,
  -50.9744,
  -50.9895,
  -51.0053,
  -51.0214,
  -51.0373,
  -51.0521,
  -51.0653,
  -51.0766,
  -51.0861,
  -51.0941,
  -51.1011,
  -51.1076,
  -51.1139,
  -51.1203,
  -51.1266,
  -51.1323,
  -51.1358,
  -51.1383,
  -51.1385,
  -51.1362,
  -51.1321,
  -51.1259,
  -51.1177,
  -51.1074,
  -51.0954,
  -51.0823,
  -51.0687,
  -51.0549,
  -51.0414,
  -51.0284,
  -51.0157,
  -51.0033,
  -50.9912,
  -50.9791,
  -50.9672,
  -50.9554,
  -50.9436,
  -50.9314,
  -50.9185,
  -50.9044,
  -50.8891,
  -50.8723,
  -50.8539,
  -50.8339,
  -50.8126,
  -50.7899,
  -50.7662,
  -50.7409,
  -50.7164,
  -50.6922,
  -50.6686,
  -50.6458,
  -50.6232,
  -50.6007,
  -50.5776,
  -50.5536,
  -50.529,
  -50.5042,
  -50.48,
  -50.4564,
  -50.4331,
  -50.4097,
  -50.3858,
  -50.3611,
  -50.3359,
  -50.3102,
  -50.2843,
  -50.2583,
  -50.2325,
  -50.2071,
  -50.1829,
  -50.1601,
  -50.1386,
  -50.1181,
  -50.0981,
  -50.0785,
  -50.0588,
  -50.0395,
  -50.0199,
  -50.0003,
  -49.98,
  -49.9588,
  -49.9364,
  -49.9132,
  -49.8894,
  -49.8645,
  -49.8404,
  -49.816,
  -49.7919,
  -49.7684,
  -49.7462,
  -49.7256,
  -49.7069,
  -49.69,
  -49.6746,
  -49.6602,
  -49.646,
  -49.6313,
  -49.6159,
  -49.6002,
  -49.584,
  -49.5679,
  -49.5522,
  -49.537,
  -49.522,
  -49.5071,
  -49.4919,
  -49.4764,
  -49.4609,
  -49.4455,
  -49.4307,
  -49.4166,
  -49.4033,
  -49.3908,
  -49.3796,
  -49.3699,
  -48.6146,
  -48.68,
  -48.7415,
  -48.7999,
  -48.8531,
  -48.901,
  -48.943,
  -48.9793,
  -49.0101,
  -49.0349,
  -49.0545,
  -49.0691,
  -49.0795,
  -49.0862,
  -49.0898,
  -49.0913,
  -49.0898,
  -49.0885,
  -49.0876,
  -49.0879,
  -49.0901,
  -49.0944,
  -49.1004,
  -49.1073,
  -49.1142,
  -49.1207,
  -49.1271,
  -49.1335,
  -49.1403,
  -49.1479,
  -49.1563,
  -49.1652,
  -49.1739,
  -49.1846,
  -49.1967,
  -49.2105,
  -49.2257,
  -49.2418,
  -49.2582,
  -49.2743,
  -49.2896,
  -49.3039,
  -49.317,
  -49.3288,
  -49.3397,
  -49.3499,
  -49.3594,
  -49.3685,
  -49.376,
  -49.384,
  -49.392,
  -49.4002,
  -49.4097,
  -49.4208,
  -49.4339,
  -49.4487,
  -49.4648,
  -49.4811,
  -49.4965,
  -49.5098,
  -49.5203,
  -49.5276,
  -49.5314,
  -49.5316,
  -49.5286,
  -49.5221,
  -49.5153,
  -49.5086,
  -49.5031,
  -49.4995,
  -49.4981,
  -49.4992,
  -49.5028,
  -49.5088,
  -49.5167,
  -49.5259,
  -49.5356,
  -49.5453,
  -49.5544,
  -49.5625,
  -49.5696,
  -49.5759,
  -49.5808,
  -49.5868,
  -49.593,
  -49.5994,
  -49.6059,
  -49.6119,
  -49.6173,
  -49.622,
  -49.626,
  -49.6296,
  -49.633,
  -49.6374,
  -49.6424,
  -49.649,
  -49.6571,
  -49.6665,
  -49.6766,
  -49.6864,
  -49.6952,
  -49.7015,
  -49.7076,
  -49.7128,
  -49.7177,
  -49.7222,
  -49.7266,
  -49.731,
  -49.7357,
  -49.7411,
  -49.7479,
  -49.7561,
  -49.7661,
  -49.7776,
  -49.79,
  -49.8026,
  -49.8148,
  -49.8261,
  -49.8364,
  -49.8461,
  -49.8555,
  -49.8643,
  -49.8744,
  -49.8854,
  -49.8981,
  -49.9133,
  -49.9308,
  -49.9512,
  -49.974,
  -49.9983,
  -50.0232,
  -50.0479,
  -50.0717,
  -50.0944,
  -50.1163,
  -50.1378,
  -50.1593,
  -50.1808,
  -50.2027,
  -50.2245,
  -50.246,
  -50.2663,
  -50.2849,
  -50.3036,
  -50.3214,
  -50.339,
  -50.3567,
  -50.3749,
  -50.3939,
  -50.4142,
  -50.436,
  -50.459,
  -50.4834,
  -50.5083,
  -50.5328,
  -50.5565,
  -50.5786,
  -50.5988,
  -50.6172,
  -50.6338,
  -50.649,
  -50.6633,
  -50.6773,
  -50.6919,
  -50.7077,
  -50.7239,
  -50.7427,
  -50.7628,
  -50.7844,
  -50.8072,
  -50.8305,
  -50.8539,
  -50.8769,
  -50.8992,
  -50.9203,
  -50.9404,
  -50.9593,
  -50.9772,
  -50.994,
  -51.0098,
  -51.0247,
  -51.0389,
  -51.0522,
  -51.0648,
  -51.0776,
  -51.0911,
  -51.1056,
  -51.1207,
  -51.1361,
  -51.1512,
  -51.1654,
  -51.1769,
  -51.1876,
  -51.1965,
  -51.2039,
  -51.2103,
  -51.2164,
  -51.2223,
  -51.2285,
  -51.2348,
  -51.2409,
  -51.2461,
  -51.2494,
  -51.2504,
  -51.2487,
  -51.2446,
  -51.2382,
  -51.2293,
  -51.2184,
  -51.2059,
  -51.1923,
  -51.1783,
  -51.1643,
  -51.1505,
  -51.1373,
  -51.1243,
  -51.1117,
  -51.0995,
  -51.0871,
  -51.0746,
  -51.0608,
  -51.0479,
  -51.0347,
  -51.0207,
  -51.0057,
  -50.9896,
  -50.9719,
  -50.9526,
  -50.9316,
  -50.9091,
  -50.8853,
  -50.8605,
  -50.8352,
  -50.81,
  -50.7851,
  -50.761,
  -50.7376,
  -50.7144,
  -50.6907,
  -50.6665,
  -50.6411,
  -50.6151,
  -50.5882,
  -50.5619,
  -50.536,
  -50.5106,
  -50.485,
  -50.4589,
  -50.4321,
  -50.4049,
  -50.3776,
  -50.3503,
  -50.3232,
  -50.2966,
  -50.271,
  -50.2455,
  -50.2226,
  -50.2012,
  -50.1809,
  -50.1613,
  -50.1416,
  -50.122,
  -50.1027,
  -50.0835,
  -50.064,
  -50.0436,
  -50.0222,
  -49.9995,
  -49.9759,
  -49.9518,
  -49.9276,
  -49.9034,
  -49.8791,
  -49.8553,
  -49.832,
  -49.8099,
  -49.7893,
  -49.7703,
  -49.7528,
  -49.7366,
  -49.7214,
  -49.7065,
  -49.6914,
  -49.6758,
  -49.6598,
  -49.6436,
  -49.6273,
  -49.6113,
  -49.5953,
  -49.5793,
  -49.5631,
  -49.5464,
  -49.5293,
  -49.5122,
  -49.4955,
  -49.4795,
  -49.4643,
  -49.45,
  -49.4366,
  -49.4246,
  -49.4144,
  -48.6156,
  -48.6804,
  -48.7422,
  -48.8,
  -48.8536,
  -48.9028,
  -48.9469,
  -48.9858,
  -49.019,
  -49.0464,
  -49.068,
  -49.0835,
  -49.095,
  -49.1029,
  -49.1073,
  -49.1093,
  -49.109,
  -49.1079,
  -49.107,
  -49.1076,
  -49.1102,
  -49.115,
  -49.1215,
  -49.1286,
  -49.1356,
  -49.1423,
  -49.1476,
  -49.154,
  -49.1611,
  -49.1692,
  -49.1783,
  -49.1884,
  -49.1994,
  -49.2115,
  -49.225,
  -49.24,
  -49.2564,
  -49.2737,
  -49.2912,
  -49.3083,
  -49.3244,
  -49.3392,
  -49.3519,
  -49.3643,
  -49.3758,
  -49.3867,
  -49.3971,
  -49.4066,
  -49.4152,
  -49.4229,
  -49.4302,
  -49.4378,
  -49.4466,
  -49.4575,
  -49.4707,
  -49.4858,
  -49.5026,
  -49.5197,
  -49.5354,
  -49.5504,
  -49.563,
  -49.5726,
  -49.5786,
  -49.5808,
  -49.5795,
  -49.5753,
  -49.5697,
  -49.5638,
  -49.5589,
  -49.5555,
  -49.5542,
  -49.555,
  -49.5584,
  -49.5638,
  -49.5712,
  -49.5799,
  -49.5882,
  -49.5975,
  -49.6063,
  -49.6142,
  -49.6212,
  -49.6278,
  -49.6344,
  -49.6413,
  -49.6488,
  -49.6569,
  -49.6652,
  -49.6732,
  -49.681,
  -49.6883,
  -49.695,
  -49.7013,
  -49.7078,
  -49.7142,
  -49.72,
  -49.7279,
  -49.7373,
  -49.7475,
  -49.7583,
  -49.7684,
  -49.7773,
  -49.7845,
  -49.79,
  -49.7944,
  -49.7981,
  -49.8013,
  -49.8043,
  -49.8075,
  -49.8113,
  -49.8166,
  -49.8237,
  -49.8333,
  -49.8451,
  -49.8581,
  -49.8735,
  -49.8895,
  -49.9053,
  -49.9205,
  -49.9347,
  -49.9479,
  -49.9608,
  -49.9733,
  -49.9859,
  -49.9986,
  -50.0124,
  -50.0284,
  -50.0461,
  -50.0663,
  -50.0883,
  -50.1118,
  -50.1358,
  -50.1596,
  -50.1827,
  -50.2049,
  -50.2254,
  -50.2464,
  -50.2672,
  -50.2882,
  -50.3097,
  -50.3311,
  -50.3522,
  -50.3725,
  -50.3924,
  -50.4115,
  -50.4299,
  -50.4479,
  -50.4661,
  -50.4849,
  -50.5047,
  -50.5257,
  -50.5484,
  -50.5724,
  -50.5976,
  -50.6232,
  -50.6485,
  -50.6727,
  -50.6954,
  -50.7153,
  -50.7344,
  -50.7518,
  -50.7678,
  -50.783,
  -50.7981,
  -50.8139,
  -50.8309,
  -50.8491,
  -50.8687,
  -50.8891,
  -50.9108,
  -50.9332,
  -50.9561,
  -50.9792,
  -51.0019,
  -51.0237,
  -51.0445,
  -51.0643,
  -51.0831,
  -51.1009,
  -51.1179,
  -51.1338,
  -51.1492,
  -51.1623,
  -51.1753,
  -51.1877,
  -51.1999,
  -51.2128,
  -51.2264,
  -51.2408,
  -51.2556,
  -51.2701,
  -51.2835,
  -51.2955,
  -51.3056,
  -51.3138,
  -51.3205,
  -51.3263,
  -51.3317,
  -51.337,
  -51.3429,
  -51.3491,
  -51.3555,
  -51.3615,
  -51.3659,
  -51.3678,
  -51.3669,
  -51.3628,
  -51.3559,
  -51.3462,
  -51.3344,
  -51.3201,
  -51.306,
  -51.2916,
  -51.2773,
  -51.2633,
  -51.2498,
  -51.2366,
  -51.2242,
  -51.2117,
  -51.1991,
  -51.1859,
  -51.1726,
  -51.1587,
  -51.1443,
  -51.1293,
  -51.1133,
  -51.0961,
  -51.0774,
  -51.0569,
  -51.0345,
  -51.0106,
  -50.9854,
  -50.9594,
  -50.933,
  -50.9069,
  -50.8813,
  -50.8565,
  -50.8323,
  -50.8084,
  -50.784,
  -50.7589,
  -50.7324,
  -50.7048,
  -50.6753,
  -50.6467,
  -50.6184,
  -50.5905,
  -50.5625,
  -50.5343,
  -50.5057,
  -50.477,
  -50.4483,
  -50.4198,
  -50.392,
  -50.3648,
  -50.3387,
  -50.3139,
  -50.2908,
  -50.2693,
  -50.2487,
  -50.2287,
  -50.2089,
  -50.1893,
  -50.1699,
  -50.1506,
  -50.1309,
  -50.1102,
  -50.0884,
  -50.0654,
  -50.0414,
  -50.0169,
  -49.9924,
  -49.968,
  -49.944,
  -49.9205,
  -49.8976,
  -49.8759,
  -49.8553,
  -49.8361,
  -49.8182,
  -49.8014,
  -49.7856,
  -49.7701,
  -49.7536,
  -49.7378,
  -49.7217,
  -49.7056,
  -49.6892,
  -49.6726,
  -49.6558,
  -49.6387,
  -49.6212,
  -49.603,
  -49.5846,
  -49.5662,
  -49.5484,
  -49.5313,
  -49.5151,
  -49.4999,
  -49.4857,
  -49.4732,
  -49.4625,
  -48.6166,
  -48.6806,
  -48.7417,
  -48.7995,
  -48.8535,
  -48.9028,
  -48.9486,
  -48.9896,
  -49.025,
  -49.0547,
  -49.0786,
  -49.0969,
  -49.1104,
  -49.1197,
  -49.1254,
  -49.1281,
  -49.1286,
  -49.1281,
  -49.1279,
  -49.1289,
  -49.1311,
  -49.1361,
  -49.1427,
  -49.15,
  -49.1571,
  -49.1638,
  -49.1702,
  -49.177,
  -49.1846,
  -49.1933,
  -49.2032,
  -49.2143,
  -49.2266,
  -49.24,
  -49.2548,
  -49.2709,
  -49.2873,
  -49.3056,
  -49.3239,
  -49.3418,
  -49.3585,
  -49.3741,
  -49.3885,
  -49.4019,
  -49.4143,
  -49.426,
  -49.437,
  -49.4471,
  -49.4559,
  -49.4636,
  -49.4706,
  -49.4778,
  -49.4854,
  -49.4961,
  -49.5092,
  -49.5245,
  -49.5415,
  -49.5594,
  -49.5772,
  -49.5939,
  -49.6087,
  -49.6207,
  -49.6293,
  -49.6341,
  -49.635,
  -49.6329,
  -49.6289,
  -49.6244,
  -49.6204,
  -49.6166,
  -49.6155,
  -49.6163,
  -49.6191,
  -49.6239,
  -49.6305,
  -49.6384,
  -49.6469,
  -49.6554,
  -49.6634,
  -49.6706,
  -49.6772,
  -49.6835,
  -49.6903,
  -49.6978,
  -49.7062,
  -49.7155,
  -49.7255,
  -49.7347,
  -49.7448,
  -49.7547,
  -49.7643,
  -49.7738,
  -49.7831,
  -49.7923,
  -49.8017,
  -49.8116,
  -49.8223,
  -49.8336,
  -49.8449,
  -49.8554,
  -49.8642,
  -49.8711,
  -49.8762,
  -49.8798,
  -49.8824,
  -49.8845,
  -49.8853,
  -49.8874,
  -49.8905,
  -49.8954,
  -49.9028,
  -49.9133,
  -49.927,
  -49.9434,
  -49.9616,
  -49.9807,
  -50.0001,
  -50.0188,
  -50.0367,
  -50.0537,
  -50.0699,
  -50.0854,
  -50.1004,
  -50.1153,
  -50.1308,
  -50.1474,
  -50.1646,
  -50.1846,
  -50.2061,
  -50.2288,
  -50.2519,
  -50.2749,
  -50.2974,
  -50.3191,
  -50.3402,
  -50.3608,
  -50.3813,
  -50.4019,
  -50.4228,
  -50.4439,
  -50.4648,
  -50.4853,
  -50.5054,
  -50.525,
  -50.5442,
  -50.5629,
  -50.5817,
  -50.6011,
  -50.6206,
  -50.6426,
  -50.6662,
  -50.6912,
  -50.7172,
  -50.7435,
  -50.7693,
  -50.794,
  -50.8171,
  -50.8386,
  -50.8584,
  -50.8766,
  -50.8937,
  -50.9102,
  -50.9266,
  -50.9438,
  -50.9619,
  -50.9811,
  -51.0012,
  -51.0218,
  -51.0431,
  -51.0649,
  -51.0872,
  -51.1096,
  -51.1308,
  -51.1523,
  -51.173,
  -51.1929,
  -51.2118,
  -51.2299,
  -51.2472,
  -51.2635,
  -51.2788,
  -51.2928,
  -51.3055,
  -51.3173,
  -51.329,
  -51.3411,
  -51.3541,
  -51.368,
  -51.3821,
  -51.396,
  -51.4089,
  -51.4203,
  -51.4298,
  -51.4373,
  -51.4434,
  -51.4485,
  -51.4532,
  -51.458,
  -51.4624,
  -51.4686,
  -51.4753,
  -51.4818,
  -51.4869,
  -51.4895,
  -51.4889,
  -51.4849,
  -51.4775,
  -51.4671,
  -51.4543,
  -51.44,
  -51.425,
  -51.41,
  -51.3953,
  -51.381,
  -51.3674,
  -51.3543,
  -51.3418,
  -51.3293,
  -51.3166,
  -51.3032,
  -51.2892,
  -51.2747,
  -51.2595,
  -51.2435,
  -51.2265,
  -51.2082,
  -51.1881,
  -51.166,
  -51.1421,
  -51.1155,
  -51.0887,
  -51.0612,
  -51.0335,
  -51.0062,
  -50.9796,
  -50.9538,
  -50.9288,
  -50.904,
  -50.8789,
  -50.8529,
  -50.8254,
  -50.7965,
  -50.7664,
  -50.7358,
  -50.7051,
  -50.6747,
  -50.6445,
  -50.6143,
  -50.5841,
  -50.5541,
  -50.5244,
  -50.4952,
  -50.4666,
  -50.4388,
  -50.4121,
  -50.387,
  -50.3634,
  -50.3413,
  -50.3201,
  -50.2995,
  -50.2792,
  -50.2592,
  -50.2392,
  -50.2193,
  -50.199,
  -50.1778,
  -50.1546,
  -50.1313,
  -50.1071,
  -50.0825,
  -50.0579,
  -50.0336,
  -50.0098,
  -49.9865,
  -49.9639,
  -49.9423,
  -49.9218,
  -49.9025,
  -49.8844,
  -49.8676,
  -49.8515,
  -49.8359,
  -49.8203,
  -49.8045,
  -49.7884,
  -49.772,
  -49.7552,
  -49.738,
  -49.7203,
  -49.7021,
  -49.6834,
  -49.6641,
  -49.6445,
  -49.6251,
  -49.6061,
  -49.5879,
  -49.5706,
  -49.5545,
  -49.5397,
  -49.5267,
  -49.5158,
  -48.6131,
  -48.6772,
  -48.7383,
  -48.7965,
  -48.8514,
  -48.9029,
  -48.9505,
  -48.9935,
  -49.0313,
  -49.0634,
  -49.0894,
  -49.1098,
  -49.1252,
  -49.1362,
  -49.1433,
  -49.1463,
  -49.1482,
  -49.1487,
  -49.1493,
  -49.1509,
  -49.1544,
  -49.1597,
  -49.1665,
  -49.1738,
  -49.1811,
  -49.1882,
  -49.1951,
  -49.2025,
  -49.2108,
  -49.2202,
  -49.2297,
  -49.2419,
  -49.2552,
  -49.2698,
  -49.2856,
  -49.3027,
  -49.321,
  -49.34,
  -49.3591,
  -49.3776,
  -49.3951,
  -49.4114,
  -49.4267,
  -49.4412,
  -49.4548,
  -49.4673,
  -49.4778,
  -49.4884,
  -49.4974,
  -49.5052,
  -49.5125,
  -49.5196,
  -49.5282,
  -49.5389,
  -49.5521,
  -49.5675,
  -49.5847,
  -49.6031,
  -49.6219,
  -49.6401,
  -49.657,
  -49.6715,
  -49.6829,
  -49.6895,
  -49.6931,
  -49.6933,
  -49.6914,
  -49.6886,
  -49.686,
  -49.684,
  -49.6832,
  -49.6841,
  -49.6866,
  -49.6907,
  -49.6963,
  -49.7031,
  -49.7106,
  -49.7181,
  -49.7251,
  -49.7314,
  -49.7362,
  -49.742,
  -49.7485,
  -49.7561,
  -49.7651,
  -49.7754,
  -49.7868,
  -49.7988,
  -49.8111,
  -49.8235,
  -49.836,
  -49.8487,
  -49.8613,
  -49.8737,
  -49.886,
  -49.8982,
  -49.9105,
  -49.923,
  -49.935,
  -49.9448,
  -49.9538,
  -49.9609,
  -49.9657,
  -49.9692,
  -49.9711,
  -49.9721,
  -49.9728,
  -49.9742,
  -49.9765,
  -49.9807,
  -49.9882,
  -49.9994,
  -50.0148,
  -50.0334,
  -50.0544,
  -50.0767,
  -50.0991,
  -50.1212,
  -50.1425,
  -50.1618,
  -50.1811,
  -50.1994,
  -50.217,
  -50.234,
  -50.2513,
  -50.2693,
  -50.288,
  -50.3078,
  -50.3287,
  -50.3505,
  -50.3729,
  -50.3952,
  -50.4172,
  -50.4386,
  -50.4595,
  -50.48,
  -50.5003,
  -50.5207,
  -50.5414,
  -50.5622,
  -50.5819,
  -50.6025,
  -50.623,
  -50.6435,
  -50.6637,
  -50.6834,
  -50.7029,
  -50.7227,
  -50.7437,
  -50.7665,
  -50.7911,
  -50.8172,
  -50.8441,
  -50.871,
  -50.8975,
  -50.9224,
  -50.9457,
  -50.9676,
  -50.988,
  -51.0071,
  -51.0253,
  -51.0434,
  -51.0613,
  -51.079,
  -51.0985,
  -51.1187,
  -51.1393,
  -51.1599,
  -51.1806,
  -51.2014,
  -51.2225,
  -51.2442,
  -51.2658,
  -51.2871,
  -51.308,
  -51.3282,
  -51.3476,
  -51.3662,
  -51.3839,
  -51.4006,
  -51.4159,
  -51.4296,
  -51.4419,
  -51.4533,
  -51.4643,
  -51.4759,
  -51.4885,
  -51.502,
  -51.5148,
  -51.5287,
  -51.5409,
  -51.5519,
  -51.5607,
  -51.5676,
  -51.5728,
  -51.577,
  -51.581,
  -51.5851,
  -51.5899,
  -51.5957,
  -51.6025,
  -51.6092,
  -51.6147,
  -51.6178,
  -51.6174,
  -51.6133,
  -51.6055,
  -51.5942,
  -51.5801,
  -51.5646,
  -51.5486,
  -51.5328,
  -51.5177,
  -51.5033,
  -51.4896,
  -51.4767,
  -51.4643,
  -51.451,
  -51.4382,
  -51.4246,
  -51.4101,
  -51.3948,
  -51.3787,
  -51.3618,
  -51.3436,
  -51.324,
  -51.3025,
  -51.2789,
  -51.2532,
  -51.2258,
  -51.1972,
  -51.1681,
  -51.139,
  -51.1104,
  -51.0827,
  -51.0558,
  -51.0297,
  -51.0038,
  -50.9779,
  -50.9511,
  -50.9228,
  -50.8928,
  -50.8612,
  -50.8284,
  -50.7954,
  -50.7627,
  -50.7301,
  -50.6982,
  -50.6668,
  -50.6359,
  -50.6057,
  -50.575,
  -50.5458,
  -50.5175,
  -50.4901,
  -50.4644,
  -50.4399,
  -50.4167,
  -50.3944,
  -50.3728,
  -50.3516,
  -50.3307,
  -50.3099,
  -50.2891,
  -50.2678,
  -50.2458,
  -50.2229,
  -50.1992,
  -50.1749,
  -50.1503,
  -50.1258,
  -50.1016,
  -50.0779,
  -50.0548,
  -50.0323,
  -50.0108,
  -49.9903,
  -49.9711,
  -49.9533,
  -49.9367,
  -49.921,
  -49.9056,
  -49.8901,
  -49.8742,
  -49.8579,
  -49.8411,
  -49.8238,
  -49.8057,
  -49.787,
  -49.7678,
  -49.748,
  -49.7279,
  -49.7076,
  -49.6875,
  -49.6677,
  -49.6486,
  -49.6294,
  -49.6125,
  -49.5972,
  -49.5839,
  -49.573,
  -48.6062,
  -48.6709,
  -48.733,
  -48.7923,
  -48.8485,
  -48.9018,
  -48.9514,
  -48.9966,
  -49.0366,
  -49.0699,
  -49.0983,
  -49.121,
  -49.1385,
  -49.1514,
  -49.1605,
  -49.1665,
  -49.17,
  -49.1721,
  -49.1737,
  -49.1761,
  -49.1798,
  -49.185,
  -49.1916,
  -49.1989,
  -49.2053,
  -49.2128,
  -49.2205,
  -49.2286,
  -49.2377,
  -49.2481,
  -49.2597,
  -49.2727,
  -49.2872,
  -49.3029,
  -49.3198,
  -49.3379,
  -49.357,
  -49.3768,
  -49.3966,
  -49.4157,
  -49.4328,
  -49.45,
  -49.4663,
  -49.4817,
  -49.4963,
  -49.5095,
  -49.5218,
  -49.5328,
  -49.5424,
  -49.5507,
  -49.5584,
  -49.5663,
  -49.5752,
  -49.586,
  -49.5991,
  -49.6143,
  -49.6314,
  -49.6491,
  -49.6686,
  -49.6881,
  -49.7068,
  -49.7239,
  -49.7381,
  -49.7487,
  -49.7551,
  -49.758,
  -49.7584,
  -49.7575,
  -49.7563,
  -49.7553,
  -49.7551,
  -49.7559,
  -49.758,
  -49.7615,
  -49.7653,
  -49.771,
  -49.7774,
  -49.7839,
  -49.7899,
  -49.7952,
  -49.8002,
  -49.8053,
  -49.8113,
  -49.8186,
  -49.8277,
  -49.8385,
  -49.8509,
  -49.8645,
  -49.8787,
  -49.8934,
  -49.9086,
  -49.9243,
  -49.9391,
  -49.9547,
  -49.9699,
  -49.9847,
  -49.9992,
  -50.013,
  -50.0259,
  -50.0372,
  -50.0467,
  -50.0542,
  -50.0594,
  -50.0629,
  -50.0648,
  -50.0657,
  -50.0661,
  -50.067,
  -50.0689,
  -50.0732,
  -50.0809,
  -50.092,
  -50.1087,
  -50.1292,
  -50.1524,
  -50.1772,
  -50.2022,
  -50.227,
  -50.251,
  -50.274,
  -50.2959,
  -50.3166,
  -50.3364,
  -50.3554,
  -50.3742,
  -50.3934,
  -50.413,
  -50.4332,
  -50.4541,
  -50.4756,
  -50.4975,
  -50.5192,
  -50.5397,
  -50.5609,
  -50.5816,
  -50.6021,
  -50.6225,
  -50.643,
  -50.6637,
  -50.6844,
  -50.7052,
  -50.7259,
  -50.7469,
  -50.7682,
  -50.7896,
  -50.8105,
  -50.8309,
  -50.8515,
  -50.8731,
  -50.8967,
  -50.9221,
  -50.9492,
  -50.9769,
  -51.0045,
  -51.0301,
  -51.0554,
  -51.079,
  -51.1013,
  -51.1224,
  -51.1424,
  -51.1619,
  -51.1814,
  -51.2009,
  -51.2208,
  -51.2414,
  -51.2623,
  -51.283,
  -51.3032,
  -51.3232,
  -51.3431,
  -51.3634,
  -51.3845,
  -51.4059,
  -51.4274,
  -51.4487,
  -51.4694,
  -51.4892,
  -51.5082,
  -51.5263,
  -51.5422,
  -51.5575,
  -51.5712,
  -51.5832,
  -51.5942,
  -51.6049,
  -51.6161,
  -51.6283,
  -51.6416,
  -51.6553,
  -51.669,
  -51.6814,
  -51.6917,
  -51.6998,
  -51.7059,
  -51.7105,
  -51.7143,
  -51.7177,
  -51.7213,
  -51.7256,
  -51.731,
  -51.7374,
  -51.7438,
  -51.7491,
  -51.752,
  -51.7515,
  -51.747,
  -51.7374,
  -51.7252,
  -51.71,
  -51.6932,
  -51.6761,
  -51.6595,
  -51.6438,
  -51.6292,
  -51.6154,
  -51.6026,
  -51.5905,
  -51.5784,
  -51.5657,
  -51.5521,
  -51.5373,
  -51.5214,
  -51.5046,
  -51.4864,
  -51.4672,
  -51.446,
  -51.423,
  -51.3977,
  -51.3702,
  -51.341,
  -51.3106,
  -51.2797,
  -51.2491,
  -51.2192,
  -51.1902,
  -51.1621,
  -51.1348,
  -51.1079,
  -51.0799,
  -51.0521,
  -51.023,
  -50.9918,
  -50.9586,
  -50.9241,
  -50.889,
  -50.854,
  -50.8196,
  -50.786,
  -50.7533,
  -50.7215,
  -50.6905,
  -50.6602,
  -50.6306,
  -50.6018,
  -50.5741,
  -50.5475,
  -50.5221,
  -50.4976,
  -50.474,
  -50.4511,
  -50.429,
  -50.4067,
  -50.3847,
  -50.3626,
  -50.3401,
  -50.3169,
  -50.2932,
  -50.2689,
  -50.2443,
  -50.2196,
  -50.1951,
  -50.171,
  -50.1472,
  -50.124,
  -50.1014,
  -50.0797,
  -50.0592,
  -50.0391,
  -50.0216,
  -50.0054,
  -49.9903,
  -49.9754,
  -49.9602,
  -49.9441,
  -49.9278,
  -49.9108,
  -49.8929,
  -49.8743,
  -49.8549,
  -49.8349,
  -49.8145,
  -49.7938,
  -49.7732,
  -49.7527,
  -49.7326,
  -49.7129,
  -49.6942,
  -49.6768,
  -49.6614,
  -49.6481,
  -49.6374,
  -48.5943,
  -48.6606,
  -48.7243,
  -48.7855,
  -48.843,
  -48.8984,
  -48.9503,
  -48.9979,
  -49.0404,
  -49.0773,
  -49.108,
  -49.1331,
  -49.1528,
  -49.1681,
  -49.1795,
  -49.1878,
  -49.1934,
  -49.1972,
  -49.2002,
  -49.2023,
  -49.2061,
  -49.2112,
  -49.2174,
  -49.2245,
  -49.2322,
  -49.2402,
  -49.2487,
  -49.2578,
  -49.2679,
  -49.2792,
  -49.2918,
  -49.306,
  -49.3217,
  -49.3387,
  -49.3559,
  -49.3751,
  -49.3951,
  -49.4157,
  -49.4362,
  -49.4559,
  -49.4747,
  -49.4925,
  -49.5095,
  -49.5257,
  -49.5409,
  -49.5551,
  -49.568,
  -49.5797,
  -49.5901,
  -49.5995,
  -49.6072,
  -49.6159,
  -49.6255,
  -49.6365,
  -49.6494,
  -49.6642,
  -49.681,
  -49.6996,
  -49.7195,
  -49.74,
  -49.7605,
  -49.7797,
  -49.7966,
  -49.8101,
  -49.8195,
  -49.8251,
  -49.8279,
  -49.828,
  -49.8282,
  -49.8281,
  -49.8284,
  -49.8293,
  -49.8312,
  -49.8342,
  -49.8382,
  -49.843,
  -49.8485,
  -49.854,
  -49.8592,
  -49.8637,
  -49.8679,
  -49.8723,
  -49.8776,
  -49.8844,
  -49.8933,
  -49.9034,
  -49.9165,
  -49.9312,
  -49.9471,
  -49.9639,
  -49.9816,
  -49.9999,
  -50.0186,
  -50.0371,
  -50.0551,
  -50.0725,
  -50.0891,
  -50.1047,
  -50.1189,
  -50.1312,
  -50.1416,
  -50.1497,
  -50.1557,
  -50.1597,
  -50.1611,
  -50.1625,
  -50.1636,
  -50.1649,
  -50.1674,
  -50.1723,
  -50.1808,
  -50.1939,
  -50.2117,
  -50.2337,
  -50.2585,
  -50.285,
  -50.312,
  -50.3388,
  -50.3648,
  -50.3897,
  -50.4134,
  -50.4359,
  -50.4572,
  -50.4778,
  -50.4971,
  -50.5176,
  -50.5385,
  -50.5597,
  -50.581,
  -50.6026,
  -50.6242,
  -50.6456,
  -50.6667,
  -50.6876,
  -50.7082,
  -50.7289,
  -50.7497,
  -50.7705,
  -50.7915,
  -50.8124,
  -50.8334,
  -50.8545,
  -50.876,
  -50.8982,
  -50.9205,
  -50.9425,
  -50.963,
  -50.9845,
  -51.007,
  -51.0312,
  -51.0574,
  -51.085,
  -51.1132,
  -51.1411,
  -51.1682,
  -51.1939,
  -51.2182,
  -51.2413,
  -51.2635,
  -51.2848,
  -51.3057,
  -51.3264,
  -51.3473,
  -51.3683,
  -51.3896,
  -51.4106,
  -51.4311,
  -51.4509,
  -51.4702,
  -51.4886,
  -51.5084,
  -51.5291,
  -51.5505,
  -51.5723,
  -51.594,
  -51.6152,
  -51.6356,
  -51.6551,
  -51.6734,
  -51.6904,
  -51.7058,
  -51.7195,
  -51.7315,
  -51.7424,
  -51.7529,
  -51.7638,
  -51.7757,
  -51.7886,
  -51.8022,
  -51.8155,
  -51.8276,
  -51.8376,
  -51.8454,
  -51.8513,
  -51.8557,
  -51.8583,
  -51.8615,
  -51.8648,
  -51.8687,
  -51.8734,
  -51.879,
  -51.8847,
  -51.8893,
  -51.8915,
  -51.8902,
  -51.885,
  -51.8756,
  -51.8623,
  -51.8461,
  -51.8283,
  -51.8102,
  -51.7928,
  -51.7767,
  -51.7618,
  -51.748,
  -51.7353,
  -51.7233,
  -51.7114,
  -51.6989,
  -51.6852,
  -51.6702,
  -51.6537,
  -51.6358,
  -51.6165,
  -51.5957,
  -51.572,
  -51.5473,
  -51.5202,
  -51.491,
  -51.4599,
  -51.4278,
  -51.3954,
  -51.3633,
  -51.332,
  -51.3018,
  -51.2725,
  -51.2439,
  -51.2158,
  -51.1876,
  -51.1587,
  -51.1284,
  -51.096,
  -51.0615,
  -51.0254,
  -50.9886,
  -50.9517,
  -50.9155,
  -50.8802,
  -50.8461,
  -50.8132,
  -50.7813,
  -50.7503,
  -50.7202,
  -50.691,
  -50.6629,
  -50.6358,
  -50.6095,
  -50.5839,
  -50.559,
  -50.5346,
  -50.5108,
  -50.4872,
  -50.4627,
  -50.439,
  -50.4149,
  -50.3903,
  -50.3653,
  -50.3401,
  -50.3148,
  -50.2896,
  -50.2647,
  -50.2402,
  -50.2161,
  -50.1926,
  -50.1697,
  -50.1478,
  -50.1272,
  -50.1082,
  -50.091,
  -50.0753,
  -50.0606,
  -50.0462,
  -50.0314,
  -50.0158,
  -49.9993,
  -49.9819,
  -49.9637,
  -49.9447,
  -49.925,
  -49.9048,
  -49.8843,
  -49.8636,
  -49.843,
  -49.8227,
  -49.8026,
  -49.7832,
  -49.7646,
  -49.7475,
  -49.7322,
  -49.7193,
  -49.7087,
  -48.5771,
  -48.6456,
  -48.7118,
  -48.7756,
  -48.8368,
  -48.895,
  -48.9493,
  -48.9994,
  -49.0445,
  -49.0841,
  -49.1176,
  -49.1452,
  -49.1675,
  -49.1844,
  -49.1984,
  -49.2092,
  -49.2171,
  -49.223,
  -49.2273,
  -49.231,
  -49.235,
  -49.2398,
  -49.2456,
  -49.2527,
  -49.2608,
  -49.2694,
  -49.279,
  -49.2893,
  -49.3005,
  -49.312,
  -49.3259,
  -49.3413,
  -49.3583,
  -49.3767,
  -49.3963,
  -49.4166,
  -49.4375,
  -49.4588,
  -49.4799,
  -49.5004,
  -49.52,
  -49.5385,
  -49.5561,
  -49.5728,
  -49.5875,
  -49.6022,
  -49.6158,
  -49.6283,
  -49.6397,
  -49.6503,
  -49.6605,
  -49.6705,
  -49.6808,
  -49.6921,
  -49.7047,
  -49.7191,
  -49.7354,
  -49.7536,
  -49.7737,
  -49.795,
  -49.8169,
  -49.8371,
  -49.8564,
  -49.8725,
  -49.8846,
  -49.8928,
  -49.8979,
  -49.9009,
  -49.9026,
  -49.9036,
  -49.9045,
  -49.9056,
  -49.9074,
  -49.91,
  -49.9133,
  -49.9174,
  -49.9219,
  -49.9267,
  -49.9311,
  -49.934,
  -49.9376,
  -49.9413,
  -49.946,
  -49.9523,
  -49.961,
  -49.972,
  -49.9857,
  -50.0015,
  -50.0187,
  -50.0373,
  -50.0569,
  -50.0774,
  -50.0985,
  -50.1194,
  -50.1402,
  -50.1602,
  -50.1792,
  -50.1957,
  -50.2115,
  -50.2252,
  -50.2367,
  -50.2462,
  -50.2535,
  -50.2587,
  -50.2624,
  -50.2651,
  -50.2676,
  -50.2703,
  -50.2741,
  -50.2803,
  -50.2899,
  -50.304,
  -50.3229,
  -50.3457,
  -50.3715,
  -50.3991,
  -50.4274,
  -50.4543,
  -50.4816,
  -50.5079,
  -50.5327,
  -50.5563,
  -50.5787,
  -50.6003,
  -50.6219,
  -50.6441,
  -50.6664,
  -50.6888,
  -50.7111,
  -50.7331,
  -50.7547,
  -50.7759,
  -50.7966,
  -50.8172,
  -50.8378,
  -50.8589,
  -50.8803,
  -50.9019,
  -50.9225,
  -50.944,
  -50.9653,
  -50.9869,
  -51.0089,
  -51.0317,
  -51.055,
  -51.0782,
  -51.1007,
  -51.1232,
  -51.1467,
  -51.1715,
  -51.1983,
  -51.2263,
  -51.2547,
  -51.283,
  -51.3106,
  -51.337,
  -51.3623,
  -51.3865,
  -51.41,
  -51.4328,
  -51.4541,
  -51.4762,
  -51.4982,
  -51.52,
  -51.5416,
  -51.5625,
  -51.583,
  -51.6023,
  -51.6212,
  -51.6402,
  -51.6598,
  -51.6805,
  -51.7021,
  -51.7244,
  -51.7466,
  -51.7683,
  -51.7891,
  -51.8088,
  -51.8272,
  -51.8442,
  -51.8596,
  -51.873,
  -51.8852,
  -51.8962,
  -51.9068,
  -51.9167,
  -51.9284,
  -51.941,
  -51.9541,
  -51.967,
  -51.9787,
  -51.9884,
  -51.9962,
  -52.0023,
  -52.0067,
  -52.0106,
  -52.0139,
  -52.0172,
  -52.0207,
  -52.0248,
  -52.0295,
  -52.0339,
  -52.0371,
  -52.0381,
  -52.0356,
  -52.0295,
  -52.0193,
  -52.0052,
  -51.9882,
  -51.9695,
  -51.9507,
  -51.9327,
  -51.9163,
  -51.9011,
  -51.8863,
  -51.8737,
  -51.8617,
  -51.8498,
  -51.8372,
  -51.8232,
  -51.8076,
  -51.7902,
  -51.7712,
  -51.7504,
  -51.7279,
  -51.7034,
  -51.6769,
  -51.6481,
  -51.6172,
  -51.5846,
  -51.551,
  -51.5172,
  -51.4839,
  -51.4515,
  -51.42,
  -51.3894,
  -51.3595,
  -51.33,
  -51.3004,
  -51.2701,
  -51.2385,
  -51.2048,
  -51.169,
  -51.1316,
  -51.0933,
  -51.0549,
  -51.017,
  -50.9791,
  -50.9435,
  -50.9095,
  -50.8765,
  -50.8448,
  -50.8141,
  -50.7846,
  -50.7561,
  -50.7284,
  -50.7013,
  -50.6745,
  -50.6482,
  -50.6223,
  -50.5967,
  -50.5714,
  -50.5461,
  -50.5204,
  -50.4946,
  -50.4682,
  -50.4417,
  -50.4152,
  -50.389,
  -50.3629,
  -50.3372,
  -50.3119,
  -50.287,
  -50.2628,
  -50.2394,
  -50.2172,
  -50.1965,
  -50.1776,
  -50.1607,
  -50.1454,
  -50.1313,
  -50.1174,
  -50.1028,
  -50.0873,
  -50.0707,
  -50.0531,
  -50.0347,
  -50.0156,
  -49.996,
  -49.976,
  -49.9549,
  -49.9346,
  -49.9146,
  -49.8949,
  -49.8757,
  -49.8572,
  -49.8396,
  -49.8233,
  -49.8088,
  -49.7964,
  -49.7861,
  -48.5574,
  -48.6289,
  -48.6983,
  -48.7654,
  -48.8298,
  -48.8911,
  -48.9484,
  -49.001,
  -49.0476,
  -49.0898,
  -49.1258,
  -49.1561,
  -49.1812,
  -49.2019,
  -49.2186,
  -49.2321,
  -49.2425,
  -49.2502,
  -49.256,
  -49.2606,
  -49.2648,
  -49.2697,
  -49.2755,
  -49.2818,
  -49.2902,
  -49.2999,
  -49.3106,
  -49.3221,
  -49.3348,
  -49.3487,
  -49.364,
  -49.3809,
  -49.3994,
  -49.4192,
  -49.44,
  -49.4611,
  -49.483,
  -49.505,
  -49.5268,
  -49.547,
  -49.5673,
  -49.5865,
  -49.6045,
  -49.6215,
  -49.6376,
  -49.6528,
  -49.667,
  -49.6804,
  -49.693,
  -49.7051,
  -49.7168,
  -49.7283,
  -49.7396,
  -49.7512,
  -49.7638,
  -49.7767,
  -49.7925,
  -49.8103,
  -49.8303,
  -49.8521,
  -49.8749,
  -49.8976,
  -49.9188,
  -49.9372,
  -49.9517,
  -49.9624,
  -49.9698,
  -49.9747,
  -49.9779,
  -49.98,
  -49.9814,
  -49.9829,
  -49.9834,
  -49.9856,
  -49.9885,
  -49.9921,
  -49.996,
  -50.0001,
  -50.0039,
  -50.0073,
  -50.0106,
  -50.014,
  -50.0183,
  -50.0242,
  -50.0328,
  -50.0444,
  -50.0586,
  -50.0752,
  -50.0936,
  -50.1135,
  -50.1336,
  -50.1555,
  -50.1783,
  -50.2016,
  -50.2244,
  -50.2469,
  -50.268,
  -50.2878,
  -50.3055,
  -50.3209,
  -50.3342,
  -50.3453,
  -50.3544,
  -50.3615,
  -50.3672,
  -50.3719,
  -50.3766,
  -50.3816,
  -50.3876,
  -50.3947,
  -50.4059,
  -50.4215,
  -50.441,
  -50.4645,
  -50.4909,
  -50.5187,
  -50.5474,
  -50.5758,
  -50.6037,
  -50.6304,
  -50.6559,
  -50.68,
  -50.703,
  -50.7258,
  -50.7487,
  -50.7721,
  -50.7959,
  -50.8197,
  -50.8431,
  -50.8658,
  -50.8867,
  -50.9079,
  -50.9286,
  -50.9491,
  -50.9699,
  -50.9914,
  -51.0135,
  -51.0361,
  -51.0587,
  -51.0811,
  -51.1031,
  -51.1254,
  -51.148,
  -51.1715,
  -51.1952,
  -51.219,
  -51.2424,
  -51.266,
  -51.2902,
  -51.3158,
  -51.3429,
  -51.3711,
  -51.3988,
  -51.4274,
  -51.4556,
  -51.4831,
  -51.5097,
  -51.5355,
  -51.5605,
  -51.585,
  -51.609,
  -51.6324,
  -51.6554,
  -51.6777,
  -51.6997,
  -51.7206,
  -51.7405,
  -51.7597,
  -51.7784,
  -51.7974,
  -51.8172,
  -51.8382,
  -51.8601,
  -51.8828,
  -51.9054,
  -51.9273,
  -51.9474,
  -51.9672,
  -51.9856,
  -52.0025,
  -52.0177,
  -52.0313,
  -52.0433,
  -52.0546,
  -52.0654,
  -52.0764,
  -52.088,
  -52.1001,
  -52.1125,
  -52.125,
  -52.1363,
  -52.1459,
  -52.154,
  -52.1603,
  -52.1653,
  -52.1694,
  -52.1732,
  -52.1766,
  -52.1799,
  -52.1833,
  -52.1868,
  -52.1899,
  -52.1915,
  -52.1898,
  -52.186,
  -52.1786,
  -52.1674,
  -52.1528,
  -52.1353,
  -52.1163,
  -52.097,
  -52.0787,
  -52.0619,
  -52.0466,
  -52.0328,
  -52.0203,
  -52.0083,
  -51.9962,
  -51.983,
  -51.9683,
  -51.9518,
  -51.9333,
  -51.9126,
  -51.8901,
  -51.8656,
  -51.8393,
  -51.811,
  -51.7805,
  -51.7481,
  -51.7141,
  -51.6793,
  -51.6445,
  -51.6102,
  -51.5767,
  -51.543,
  -51.511,
  -51.4796,
  -51.4486,
  -51.4175,
  -51.3856,
  -51.3524,
  -51.3172,
  -51.2803,
  -51.2418,
  -51.2024,
  -51.1628,
  -51.1236,
  -51.0854,
  -51.0484,
  -51.0128,
  -50.9787,
  -50.9462,
  -50.9147,
  -50.8848,
  -50.8558,
  -50.8278,
  -50.8,
  -50.7723,
  -50.7447,
  -50.7172,
  -50.6897,
  -50.6624,
  -50.635,
  -50.6073,
  -50.5791,
  -50.5509,
  -50.5226,
  -50.4945,
  -50.4667,
  -50.4392,
  -50.4121,
  -50.3855,
  -50.3595,
  -50.3333,
  -50.3094,
  -50.2869,
  -50.2661,
  -50.2473,
  -50.2304,
  -50.2152,
  -50.2011,
  -50.1871,
  -50.1726,
  -50.1571,
  -50.1404,
  -50.1227,
  -50.1043,
  -50.0854,
  -50.0662,
  -50.0468,
  -50.0274,
  -50.0082,
  -49.9892,
  -49.9709,
  -49.9533,
  -49.9366,
  -49.9208,
  -49.9061,
  -49.8927,
  -49.8812,
  -49.8713,
  -48.5351,
  -48.6101,
  -48.6832,
  -48.7531,
  -48.821,
  -48.8854,
  -48.9458,
  -49.0012,
  -49.0514,
  -49.096,
  -49.1347,
  -49.1676,
  -49.1953,
  -49.2185,
  -49.2381,
  -49.2543,
  -49.2673,
  -49.2761,
  -49.2834,
  -49.289,
  -49.2941,
  -49.2994,
  -49.3057,
  -49.3135,
  -49.3228,
  -49.3336,
  -49.3456,
  -49.3588,
  -49.3731,
  -49.3884,
  -49.4055,
  -49.4239,
  -49.4438,
  -49.4637,
  -49.4852,
  -49.5074,
  -49.5299,
  -49.5525,
  -49.5751,
  -49.5972,
  -49.6183,
  -49.638,
  -49.6564,
  -49.6737,
  -49.69,
  -49.7055,
  -49.7202,
  -49.7346,
  -49.7486,
  -49.7613,
  -49.7746,
  -49.7875,
  -49.7999,
  -49.8122,
  -49.8248,
  -49.8385,
  -49.8538,
  -49.8712,
  -49.891,
  -49.913,
  -49.9364,
  -49.9601,
  -49.9828,
  -50.003,
  -50.0196,
  -50.0326,
  -50.0413,
  -50.0481,
  -50.0527,
  -50.0557,
  -50.0577,
  -50.0593,
  -50.0609,
  -50.0629,
  -50.0655,
  -50.0687,
  -50.0722,
  -50.0757,
  -50.079,
  -50.0823,
  -50.0855,
  -50.0888,
  -50.0935,
  -50.0987,
  -50.1075,
  -50.1194,
  -50.1342,
  -50.1517,
  -50.1712,
  -50.1921,
  -50.2143,
  -50.2375,
  -50.2615,
  -50.286,
  -50.3107,
  -50.335,
  -50.3583,
  -50.3803,
  -50.4001,
  -50.4175,
  -50.4327,
  -50.4457,
  -50.4561,
  -50.4657,
  -50.474,
  -50.4816,
  -50.4892,
  -50.4973,
  -50.5063,
  -50.5169,
  -50.5301,
  -50.5468,
  -50.5672,
  -50.5911,
  -50.6173,
  -50.645,
  -50.6732,
  -50.7014,
  -50.7293,
  -50.7561,
  -50.7815,
  -50.8061,
  -50.8289,
  -50.8524,
  -50.8762,
  -50.9007,
  -50.926,
  -50.9512,
  -50.9757,
  -50.9994,
  -51.022,
  -51.0437,
  -51.0646,
  -51.0854,
  -51.1067,
  -51.1287,
  -51.1516,
  -51.1752,
  -51.199,
  -51.2225,
  -51.2457,
  -51.2688,
  -51.2922,
  -51.3151,
  -51.3392,
  -51.3634,
  -51.3875,
  -51.4117,
  -51.4367,
  -51.4629,
  -51.4902,
  -51.5185,
  -51.5474,
  -51.5763,
  -51.6055,
  -51.6341,
  -51.6622,
  -51.6896,
  -51.7166,
  -51.7429,
  -51.7685,
  -51.7933,
  -51.8172,
  -51.8403,
  -51.8625,
  -51.8836,
  -51.9032,
  -51.9215,
  -51.9405,
  -51.9597,
  -51.9798,
  -52.0012,
  -52.0235,
  -52.0462,
  -52.0689,
  -52.091,
  -52.1121,
  -52.1318,
  -52.1502,
  -52.1669,
  -52.182,
  -52.1955,
  -52.2077,
  -52.2192,
  -52.2304,
  -52.2416,
  -52.2531,
  -52.2649,
  -52.2769,
  -52.2888,
  -52.2996,
  -52.3094,
  -52.3173,
  -52.3231,
  -52.3283,
  -52.3333,
  -52.3374,
  -52.3409,
  -52.3442,
  -52.347,
  -52.3495,
  -52.3511,
  -52.351,
  -52.3485,
  -52.3432,
  -52.3345,
  -52.3226,
  -52.3074,
  -52.2897,
  -52.2705,
  -52.2512,
  -52.2328,
  -52.2159,
  -52.2007,
  -52.187,
  -52.1745,
  -52.1623,
  -52.1496,
  -52.1355,
  -52.1196,
  -52.1017,
  -52.0815,
  -52.0582,
  -52.0336,
  -52.007,
  -51.9787,
  -51.9485,
  -51.9164,
  -51.8826,
  -51.8476,
  -51.812,
  -51.7764,
  -51.7413,
  -51.7067,
  -51.6728,
  -51.6393,
  -51.6063,
  -51.5736,
  -51.5407,
  -51.5072,
  -51.4724,
  -51.4358,
  -51.3977,
  -51.3583,
  -51.318,
  -51.2775,
  -51.2372,
  -51.1978,
  -51.1597,
  -51.1229,
  -51.0877,
  -51.054,
  -51.0219,
  -50.9914,
  -50.962,
  -50.9334,
  -50.9051,
  -50.8756,
  -50.8468,
  -50.8176,
  -50.7883,
  -50.7588,
  -50.7291,
  -50.699,
  -50.6686,
  -50.6381,
  -50.6078,
  -50.5777,
  -50.5479,
  -50.5185,
  -50.4896,
  -50.4613,
  -50.4339,
  -50.4077,
  -50.383,
  -50.3601,
  -50.3392,
  -50.3202,
  -50.303,
  -50.2872,
  -50.2725,
  -50.258,
  -50.2431,
  -50.2272,
  -50.2103,
  -50.1925,
  -50.1743,
  -50.1557,
  -50.1371,
  -50.1188,
  -50.1005,
  -50.0826,
  -50.0654,
  -50.0491,
  -50.0338,
  -50.0196,
  -50.0061,
  -49.9936,
  -49.982,
  -49.9715,
  -49.9619,
  -48.5096,
  -48.5891,
  -48.6661,
  -48.7408,
  -48.8123,
  -48.8801,
  -48.9432,
  -49.0013,
  -49.0541,
  -49.101,
  -49.1422,
  -49.1777,
  -49.2071,
  -49.233,
  -49.2553,
  -49.274,
  -49.2894,
  -49.3015,
  -49.3106,
  -49.3177,
  -49.3241,
  -49.3305,
  -49.338,
  -49.347,
  -49.3576,
  -49.3698,
  -49.3834,
  -49.3973,
  -49.4134,
  -49.4306,
  -49.4491,
  -49.4687,
  -49.4895,
  -49.5112,
  -49.5335,
  -49.5563,
  -49.5793,
  -49.6028,
  -49.6262,
  -49.6492,
  -49.6711,
  -49.6916,
  -49.7105,
  -49.7268,
  -49.7433,
  -49.7592,
  -49.7744,
  -49.7897,
  -49.8049,
  -49.8201,
  -49.835,
  -49.8494,
  -49.863,
  -49.876,
  -49.889,
  -49.9027,
  -49.9178,
  -49.935,
  -49.9547,
  -49.9756,
  -49.9992,
  -50.0235,
  -50.0471,
  -50.0687,
  -50.0873,
  -50.1023,
  -50.1141,
  -50.1228,
  -50.1288,
  -50.1327,
  -50.1352,
  -50.137,
  -50.1387,
  -50.1408,
  -50.1433,
  -50.1463,
  -50.1495,
  -50.1517,
  -50.1548,
  -50.158,
  -50.1615,
  -50.1655,
  -50.1705,
  -50.1773,
  -50.1868,
  -50.1994,
  -50.215,
  -50.2334,
  -50.2538,
  -50.2757,
  -50.2988,
  -50.3227,
  -50.3475,
  -50.3729,
  -50.3988,
  -50.4235,
  -50.4488,
  -50.4727,
  -50.4946,
  -50.5143,
  -50.5318,
  -50.5471,
  -50.5606,
  -50.5732,
  -50.5846,
  -50.5956,
  -50.6067,
  -50.6183,
  -50.6307,
  -50.6442,
  -50.6598,
  -50.6781,
  -50.6989,
  -50.7226,
  -50.7474,
  -50.7744,
  -50.802,
  -50.8297,
  -50.8571,
  -50.8836,
  -50.9091,
  -50.9337,
  -50.9578,
  -50.9819,
  -51.0066,
  -51.032,
  -51.0584,
  -51.0849,
  -51.1107,
  -51.1355,
  -51.1593,
  -51.182,
  -51.2039,
  -51.2255,
  -51.2475,
  -51.2694,
  -51.2932,
  -51.3177,
  -51.3427,
  -51.3674,
  -51.3918,
  -51.416,
  -51.4401,
  -51.4643,
  -51.4887,
  -51.5133,
  -51.5378,
  -51.5626,
  -51.5884,
  -51.615,
  -51.6425,
  -51.6709,
  -51.7,
  -51.7297,
  -51.7595,
  -51.7893,
  -51.8189,
  -51.8479,
  -51.8755,
  -51.9036,
  -51.931,
  -51.9575,
  -51.9827,
  -52.0067,
  -52.0294,
  -52.0509,
  -52.0711,
  -52.0905,
  -52.1098,
  -52.1296,
  -52.1503,
  -52.172,
  -52.1944,
  -52.217,
  -52.2394,
  -52.2612,
  -52.282,
  -52.3016,
  -52.3198,
  -52.3364,
  -52.3515,
  -52.365,
  -52.3774,
  -52.3882,
  -52.3996,
  -52.4111,
  -52.4226,
  -52.4343,
  -52.4461,
  -52.4577,
  -52.4685,
  -52.4781,
  -52.4862,
  -52.4928,
  -52.4986,
  -52.5034,
  -52.5079,
  -52.5114,
  -52.5146,
  -52.5171,
  -52.5187,
  -52.519,
  -52.5173,
  -52.5133,
  -52.5064,
  -52.4966,
  -52.4837,
  -52.4681,
  -52.4504,
  -52.4313,
  -52.4122,
  -52.3929,
  -52.376,
  -52.3609,
  -52.3472,
  -52.3347,
  -52.3223,
  -52.3087,
  -52.2935,
  -52.276,
  -52.2562,
  -52.2341,
  -52.2097,
  -52.183,
  -52.1542,
  -52.1238,
  -52.0918,
  -52.0583,
  -52.0235,
  -51.9876,
  -51.9513,
  -51.9151,
  -51.8792,
  -51.8437,
  -51.8084,
  -51.7735,
  -51.7387,
  -51.7042,
  -51.6695,
  -51.6342,
  -51.5977,
  -51.5598,
  -51.5206,
  -51.4802,
  -51.4382,
  -51.397,
  -51.3559,
  -51.3157,
  -51.2765,
  -51.2388,
  -51.2026,
  -51.1682,
  -51.1353,
  -51.104,
  -51.0739,
  -51.0448,
  -51.0158,
  -50.9867,
  -50.9568,
  -50.926,
  -50.8947,
  -50.8629,
  -50.8307,
  -50.798,
  -50.7652,
  -50.7324,
  -50.6999,
  -50.6676,
  -50.6355,
  -50.6039,
  -50.5729,
  -50.5427,
  -50.5139,
  -50.4866,
  -50.4611,
  -50.4377,
  -50.4162,
  -50.3966,
  -50.3786,
  -50.3618,
  -50.3458,
  -50.3298,
  -50.3137,
  -50.2973,
  -50.2799,
  -50.2611,
  -50.2429,
  -50.2249,
  -50.2069,
  -50.1895,
  -50.1727,
  -50.1566,
  -50.1416,
  -50.1278,
  -50.1153,
  -50.1039,
  -50.0933,
  -50.0832,
  -50.0735,
  -50.0643,
  -50.0553,
  -48.4835,
  -48.5675,
  -48.6492,
  -48.7279,
  -48.8029,
  -48.8737,
  -48.9385,
  -48.9991,
  -49.054,
  -49.1031,
  -49.1464,
  -49.1844,
  -49.2176,
  -49.2463,
  -49.2715,
  -49.2929,
  -49.3107,
  -49.3249,
  -49.3359,
  -49.345,
  -49.3532,
  -49.3605,
  -49.3699,
  -49.3807,
  -49.3932,
  -49.4072,
  -49.4228,
  -49.4395,
  -49.4575,
  -49.4763,
  -49.4961,
  -49.5167,
  -49.5382,
  -49.5604,
  -49.5831,
  -49.6063,
  -49.6301,
  -49.6534,
  -49.6778,
  -49.7018,
  -49.7245,
  -49.7458,
  -49.7651,
  -49.783,
  -49.7997,
  -49.8156,
  -49.8313,
  -49.8473,
  -49.8636,
  -49.88,
  -49.8963,
  -49.9121,
  -49.9271,
  -49.9401,
  -49.9538,
  -49.9678,
  -49.9831,
  -50.0003,
  -50.0198,
  -50.0416,
  -50.0652,
  -50.0897,
  -50.1137,
  -50.1364,
  -50.1566,
  -50.1737,
  -50.1875,
  -50.1979,
  -50.2052,
  -50.21,
  -50.2121,
  -50.2145,
  -50.2165,
  -50.2189,
  -50.2217,
  -50.2247,
  -50.2277,
  -50.2306,
  -50.2337,
  -50.2371,
  -50.2409,
  -50.2455,
  -50.2513,
  -50.2592,
  -50.2697,
  -50.2833,
  -50.3,
  -50.3193,
  -50.3397,
  -50.3625,
  -50.3863,
  -50.4109,
  -50.4361,
  -50.4621,
  -50.4887,
  -50.5156,
  -50.5422,
  -50.5678,
  -50.5917,
  -50.6135,
  -50.6333,
  -50.6512,
  -50.6677,
  -50.683,
  -50.6979,
  -50.7125,
  -50.7274,
  -50.7417,
  -50.7575,
  -50.7741,
  -50.792,
  -50.8114,
  -50.8327,
  -50.856,
  -50.8812,
  -50.9075,
  -50.9345,
  -50.9614,
  -50.9882,
  -51.0141,
  -51.0394,
  -51.064,
  -51.0884,
  -51.1133,
  -51.1389,
  -51.1651,
  -51.1923,
  -51.2198,
  -51.2459,
  -51.2718,
  -51.2972,
  -51.3216,
  -51.3451,
  -51.3685,
  -51.3918,
  -51.4155,
  -51.4402,
  -51.4656,
  -51.4916,
  -51.5176,
  -51.5432,
  -51.5684,
  -51.5934,
  -51.6182,
  -51.6429,
  -51.6678,
  -51.6928,
  -51.7183,
  -51.7447,
  -51.7707,
  -51.7985,
  -51.8271,
  -51.8565,
  -51.8866,
  -51.9172,
  -51.948,
  -51.9785,
  -52.0089,
  -52.039,
  -52.069,
  -52.0984,
  -52.1268,
  -52.1537,
  -52.179,
  -52.2027,
  -52.2249,
  -52.2458,
  -52.266,
  -52.286,
  -52.3065,
  -52.3277,
  -52.3496,
  -52.3718,
  -52.3932,
  -52.4152,
  -52.4363,
  -52.4566,
  -52.4758,
  -52.4936,
  -52.51,
  -52.525,
  -52.5387,
  -52.5513,
  -52.5636,
  -52.5752,
  -52.5867,
  -52.5982,
  -52.6099,
  -52.6218,
  -52.6334,
  -52.6444,
  -52.654,
  -52.6622,
  -52.669,
  -52.6745,
  -52.6793,
  -52.6835,
  -52.687,
  -52.6901,
  -52.6923,
  -52.6923,
  -52.6917,
  -52.6888,
  -52.6834,
  -52.6752,
  -52.6642,
  -52.6504,
  -52.6343,
  -52.6164,
  -52.5976,
  -52.5787,
  -52.5606,
  -52.5439,
  -52.5288,
  -52.5151,
  -52.5023,
  -52.4892,
  -52.4747,
  -52.458,
  -52.4387,
  -52.4169,
  -52.3927,
  -52.366,
  -52.3372,
  -52.3065,
  -52.2742,
  -52.2405,
  -52.2058,
  -52.17,
  -52.1335,
  -52.0967,
  -52.0588,
  -52.0221,
  -51.9856,
  -51.9491,
  -51.9126,
  -51.876,
  -51.8396,
  -51.803,
  -51.7658,
  -51.7277,
  -51.6884,
  -51.648,
  -51.6068,
  -51.5651,
  -51.5235,
  -51.482,
  -51.4411,
  -51.4014,
  -51.363,
  -51.3262,
  -51.2911,
  -51.2575,
  -51.2254,
  -51.1945,
  -51.1645,
  -51.1346,
  -51.1044,
  -51.0733,
  -51.0408,
  -51.0077,
  -50.9736,
  -50.9388,
  -50.9036,
  -50.8684,
  -50.8334,
  -50.7985,
  -50.7638,
  -50.7283,
  -50.6943,
  -50.6612,
  -50.6293,
  -50.5989,
  -50.5705,
  -50.544,
  -50.5197,
  -50.4973,
  -50.4766,
  -50.4573,
  -50.4387,
  -50.4208,
  -50.4033,
  -50.3854,
  -50.3674,
  -50.3494,
  -50.3312,
  -50.313,
  -50.2952,
  -50.278,
  -50.2617,
  -50.2464,
  -50.2324,
  -50.2197,
  -50.2086,
  -50.1989,
  -50.1904,
  -50.1828,
  -50.1752,
  -50.1675,
  -50.1596,
  -50.1517,
  -48.4557,
  -48.5439,
  -48.6302,
  -48.7129,
  -48.7913,
  -48.8648,
  -48.9329,
  -48.9956,
  -49.0525,
  -49.1037,
  -49.1492,
  -49.1894,
  -49.2252,
  -49.2569,
  -49.285,
  -49.3092,
  -49.3286,
  -49.3451,
  -49.3585,
  -49.3697,
  -49.38,
  -49.3906,
  -49.4024,
  -49.4157,
  -49.4308,
  -49.4472,
  -49.4651,
  -49.4841,
  -49.5039,
  -49.5244,
  -49.5453,
  -49.5658,
  -49.5876,
  -49.6098,
  -49.6327,
  -49.6564,
  -49.681,
  -49.7063,
  -49.7316,
  -49.7566,
  -49.7805,
  -49.8027,
  -49.8227,
  -49.8412,
  -49.8582,
  -49.8743,
  -49.8902,
  -49.9056,
  -49.9225,
  -49.9398,
  -49.9574,
  -49.9745,
  -49.9908,
  -50.0062,
  -50.021,
  -50.0359,
  -50.0517,
  -50.0691,
  -50.0887,
  -50.1103,
  -50.1337,
  -50.158,
  -50.1822,
  -50.2055,
  -50.226,
  -50.2449,
  -50.2606,
  -50.2728,
  -50.2816,
  -50.2877,
  -50.2917,
  -50.2949,
  -50.2978,
  -50.3007,
  -50.3038,
  -50.3068,
  -50.3097,
  -50.3125,
  -50.3156,
  -50.3191,
  -50.3234,
  -50.3286,
  -50.3344,
  -50.3434,
  -50.3552,
  -50.37,
  -50.3879,
  -50.4084,
  -50.4309,
  -50.4546,
  -50.4791,
  -50.5042,
  -50.5299,
  -50.5563,
  -50.5835,
  -50.6111,
  -50.6387,
  -50.6655,
  -50.6911,
  -50.7149,
  -50.736,
  -50.7565,
  -50.7759,
  -50.7947,
  -50.813,
  -50.8312,
  -50.8496,
  -50.8682,
  -50.887,
  -50.9061,
  -50.9257,
  -50.9462,
  -50.968,
  -50.9914,
  -51.0164,
  -51.0424,
  -51.069,
  -51.0956,
  -51.122,
  -51.1477,
  -51.1717,
  -51.1965,
  -51.2212,
  -51.2463,
  -51.2723,
  -51.2994,
  -51.3273,
  -51.3554,
  -51.3835,
  -51.411,
  -51.438,
  -51.4644,
  -51.4901,
  -51.5154,
  -51.5405,
  -51.5659,
  -51.5917,
  -51.6182,
  -51.6451,
  -51.6722,
  -51.6992,
  -51.7247,
  -51.7506,
  -51.7761,
  -51.8014,
  -51.8269,
  -51.8523,
  -51.8783,
  -51.905,
  -51.9325,
  -51.9606,
  -51.9894,
  -52.0191,
  -52.0497,
  -52.0807,
  -52.112,
  -52.1434,
  -52.1748,
  -52.2064,
  -52.2381,
  -52.2697,
  -52.3002,
  -52.3292,
  -52.356,
  -52.3801,
  -52.4034,
  -52.4254,
  -52.4467,
  -52.4678,
  -52.4891,
  -52.5109,
  -52.5329,
  -52.555,
  -52.577,
  -52.5983,
  -52.619,
  -52.6382,
  -52.6566,
  -52.6738,
  -52.6898,
  -52.7046,
  -52.7184,
  -52.7314,
  -52.7438,
  -52.7556,
  -52.7673,
  -52.7789,
  -52.7907,
  -52.8028,
  -52.8149,
  -52.8253,
  -52.8354,
  -52.8438,
  -52.8508,
  -52.8563,
  -52.8606,
  -52.8643,
  -52.8674,
  -52.8702,
  -52.8722,
  -52.8727,
  -52.8712,
  -52.8673,
  -52.8609,
  -52.8517,
  -52.8396,
  -52.825,
  -52.8083,
  -52.7902,
  -52.7715,
  -52.7526,
  -52.7347,
  -52.7181,
  -52.703,
  -52.6889,
  -52.6754,
  -52.6612,
  -52.6453,
  -52.6271,
  -52.605,
  -52.5813,
  -52.555,
  -52.5263,
  -52.4956,
  -52.4631,
  -52.4291,
  -52.3941,
  -52.3582,
  -52.3217,
  -52.2845,
  -52.247,
  -52.2094,
  -52.1718,
  -52.1342,
  -52.0965,
  -52.0585,
  -52.0202,
  -51.9819,
  -51.9433,
  -51.9042,
  -51.8644,
  -51.8238,
  -51.7823,
  -51.7403,
  -51.6983,
  -51.6563,
  -51.6147,
  -51.5738,
  -51.5339,
  -51.4953,
  -51.4581,
  -51.4224,
  -51.388,
  -51.3549,
  -51.3218,
  -51.2904,
  -51.259,
  -51.2272,
  -51.1944,
  -51.1603,
  -51.1249,
  -51.0888,
  -51.0518,
  -51.0146,
  -50.9774,
  -50.9401,
  -50.903,
  -50.8659,
  -50.8291,
  -50.7929,
  -50.7578,
  -50.7241,
  -50.6922,
  -50.6624,
  -50.6347,
  -50.6091,
  -50.5854,
  -50.5633,
  -50.5421,
  -50.5218,
  -50.5019,
  -50.4821,
  -50.4621,
  -50.4421,
  -50.4225,
  -50.4034,
  -50.3847,
  -50.3669,
  -50.3502,
  -50.335,
  -50.3213,
  -50.3093,
  -50.2991,
  -50.2906,
  -50.2837,
  -50.2778,
  -50.2726,
  -50.2674,
  -50.2615,
  -50.2541,
  -50.2476,
  -48.4258,
  -48.5201,
  -48.6111,
  -48.6978,
  -48.7795,
  -48.8555,
  -48.9259,
  -48.9904,
  -49.0489,
  -49.1019,
  -49.1485,
  -49.191,
  -49.2292,
  -49.2638,
  -49.2945,
  -49.3215,
  -49.3446,
  -49.3637,
  -49.3796,
  -49.3933,
  -49.4062,
  -49.4194,
  -49.4341,
  -49.4504,
  -49.4684,
  -49.4878,
  -49.5075,
  -49.5291,
  -49.5512,
  -49.5735,
  -49.5956,
  -49.6176,
  -49.6396,
  -49.6619,
  -49.685,
  -49.7092,
  -49.7345,
  -49.7607,
  -49.7872,
  -49.8133,
  -49.8381,
  -49.8602,
  -49.8812,
  -49.9002,
  -49.9177,
  -49.9341,
  -49.9501,
  -49.9665,
  -49.9838,
  -50.0019,
  -50.0204,
  -50.0388,
  -50.0565,
  -50.0734,
  -50.0896,
  -50.1057,
  -50.1225,
  -50.1404,
  -50.159,
  -50.1806,
  -50.2037,
  -50.2277,
  -50.2521,
  -50.2759,
  -50.2985,
  -50.3189,
  -50.3364,
  -50.3504,
  -50.3609,
  -50.3685,
  -50.3741,
  -50.3785,
  -50.3824,
  -50.3862,
  -50.3896,
  -50.3917,
  -50.3945,
  -50.397,
  -50.4002,
  -50.4038,
  -50.4082,
  -50.4141,
  -50.4218,
  -50.4321,
  -50.4452,
  -50.4615,
  -50.4808,
  -50.5026,
  -50.5262,
  -50.5509,
  -50.5761,
  -50.6017,
  -50.6278,
  -50.6535,
  -50.6811,
  -50.7092,
  -50.7374,
  -50.7651,
  -50.792,
  -50.8176,
  -50.8418,
  -50.865,
  -50.8874,
  -50.9094,
  -50.9311,
  -50.9526,
  -50.974,
  -50.9955,
  -51.0168,
  -51.0379,
  -51.059,
  -51.0805,
  -51.103,
  -51.1259,
  -51.1512,
  -51.1776,
  -51.2044,
  -51.2311,
  -51.2576,
  -51.2834,
  -51.3086,
  -51.3335,
  -51.3584,
  -51.384,
  -51.4104,
  -51.4379,
  -51.4662,
  -51.4951,
  -51.5239,
  -51.5527,
  -51.5813,
  -51.6097,
  -51.6377,
  -51.6643,
  -51.6915,
  -51.7187,
  -51.7463,
  -51.7742,
  -51.8025,
  -51.8309,
  -51.859,
  -51.8867,
  -51.9138,
  -51.9403,
  -51.9664,
  -51.9924,
  -52.0184,
  -52.0449,
  -52.0718,
  -52.0993,
  -52.1276,
  -52.1568,
  -52.1868,
  -52.2175,
  -52.2488,
  -52.2803,
  -52.3112,
  -52.3435,
  -52.3766,
  -52.4103,
  -52.4439,
  -52.4766,
  -52.5076,
  -52.5364,
  -52.5628,
  -52.5877,
  -52.6112,
  -52.634,
  -52.6566,
  -52.679,
  -52.7015,
  -52.7238,
  -52.7458,
  -52.7672,
  -52.7878,
  -52.8074,
  -52.8259,
  -52.8433,
  -52.8597,
  -52.875,
  -52.8886,
  -52.9022,
  -52.9153,
  -52.9279,
  -52.94,
  -52.9517,
  -52.9635,
  -52.9756,
  -52.9882,
  -53.0009,
  -53.013,
  -53.0238,
  -53.0329,
  -53.0402,
  -53.0456,
  -53.0496,
  -53.0528,
  -53.0555,
  -53.0578,
  -53.0593,
  -53.0593,
  -53.057,
  -53.0524,
  -53.045,
  -53.0351,
  -53.0221,
  -53.0066,
  -52.9893,
  -52.97,
  -52.9511,
  -52.9324,
  -52.9146,
  -52.8979,
  -52.8822,
  -52.8674,
  -52.8526,
  -52.837,
  -52.8196,
  -52.7995,
  -52.7768,
  -52.7513,
  -52.7233,
  -52.6929,
  -52.6605,
  -52.6265,
  -52.5911,
  -52.555,
  -52.5182,
  -52.4808,
  -52.4429,
  -52.4045,
  -52.3659,
  -52.3271,
  -52.2884,
  -52.2494,
  -52.21,
  -52.1702,
  -52.13,
  -52.0894,
  -52.0486,
  -52.0061,
  -51.9642,
  -51.9218,
  -51.8793,
  -51.837,
  -51.7951,
  -51.7536,
  -51.7128,
  -51.6731,
  -51.6347,
  -51.5973,
  -51.561,
  -51.5255,
  -51.4913,
  -51.4576,
  -51.4242,
  -51.3907,
  -51.3568,
  -51.3219,
  -51.2858,
  -51.2485,
  -51.2106,
  -51.1718,
  -51.1329,
  -51.0938,
  -51.0546,
  -51.0154,
  -50.9762,
  -50.9373,
  -50.8992,
  -50.8621,
  -50.8267,
  -50.7932,
  -50.7617,
  -50.7325,
  -50.7055,
  -50.6802,
  -50.656,
  -50.6332,
  -50.6109,
  -50.5878,
  -50.5654,
  -50.5429,
  -50.5206,
  -50.4989,
  -50.4782,
  -50.4586,
  -50.4405,
  -50.424,
  -50.4096,
  -50.3973,
  -50.3872,
  -50.3793,
  -50.3732,
  -50.3685,
  -50.3647,
  -50.3617,
  -50.3581,
  -50.3539,
  -50.3492,
  -50.3444,
  -48.3956,
  -48.4954,
  -48.5912,
  -48.6817,
  -48.7667,
  -48.8444,
  -48.9169,
  -48.9829,
  -49.043,
  -49.0974,
  -49.1468,
  -49.1914,
  -49.2319,
  -49.2687,
  -49.3019,
  -49.3314,
  -49.3569,
  -49.3788,
  -49.3973,
  -49.4141,
  -49.4292,
  -49.4458,
  -49.4638,
  -49.4835,
  -49.5048,
  -49.5277,
  -49.5515,
  -49.5761,
  -49.6009,
  -49.6252,
  -49.6487,
  -49.6715,
  -49.694,
  -49.7166,
  -49.7399,
  -49.7634,
  -49.7893,
  -49.8162,
  -49.8436,
  -49.8707,
  -49.8966,
  -49.9207,
  -49.9426,
  -49.9625,
  -49.9804,
  -49.997,
  -50.0132,
  -50.0298,
  -50.0473,
  -50.0659,
  -50.0853,
  -50.1048,
  -50.1229,
  -50.1412,
  -50.1589,
  -50.1764,
  -50.1941,
  -50.2127,
  -50.2326,
  -50.2542,
  -50.2771,
  -50.3011,
  -50.3256,
  -50.35,
  -50.3735,
  -50.3954,
  -50.4146,
  -50.4306,
  -50.4432,
  -50.4519,
  -50.4593,
  -50.4653,
  -50.4706,
  -50.4752,
  -50.4791,
  -50.4823,
  -50.4849,
  -50.4873,
  -50.4901,
  -50.4936,
  -50.4984,
  -50.5047,
  -50.5132,
  -50.5246,
  -50.5391,
  -50.5569,
  -50.5768,
  -50.5999,
  -50.6247,
  -50.6503,
  -50.6762,
  -50.7024,
  -50.7289,
  -50.756,
  -50.7837,
  -50.812,
  -50.8405,
  -50.8689,
  -50.8968,
  -50.924,
  -50.9502,
  -50.9759,
  -51.0012,
  -51.0262,
  -51.0509,
  -51.0743,
  -51.0983,
  -51.122,
  -51.1454,
  -51.1682,
  -51.1907,
  -51.2134,
  -51.2369,
  -51.2617,
  -51.2879,
  -51.315,
  -51.3426,
  -51.3701,
  -51.3972,
  -51.4236,
  -51.4493,
  -51.4747,
  -51.5002,
  -51.5261,
  -51.5529,
  -51.5796,
  -51.6081,
  -51.6373,
  -51.6668,
  -51.6966,
  -51.7267,
  -51.7569,
  -51.787,
  -51.8169,
  -51.8465,
  -51.876,
  -51.9055,
  -51.9352,
  -51.9651,
  -51.995,
  -52.0247,
  -52.0538,
  -52.0821,
  -52.1097,
  -52.1367,
  -52.1634,
  -52.19,
  -52.2157,
  -52.2428,
  -52.2704,
  -52.2987,
  -52.328,
  -52.3581,
  -52.389,
  -52.4204,
  -52.4523,
  -52.4847,
  -52.518,
  -52.5524,
  -52.5877,
  -52.6231,
  -52.6577,
  -52.6905,
  -52.7211,
  -52.7495,
  -52.7761,
  -52.8015,
  -52.8262,
  -52.8505,
  -52.8745,
  -52.8981,
  -52.92,
  -52.9421,
  -52.9632,
  -52.9832,
  -53.0019,
  -53.0194,
  -53.0358,
  -53.0511,
  -53.0656,
  -53.0795,
  -53.0929,
  -53.106,
  -53.1187,
  -53.1309,
  -53.1427,
  -53.1547,
  -53.1672,
  -53.1803,
  -53.1936,
  -53.2063,
  -53.2179,
  -53.2277,
  -53.2355,
  -53.2412,
  -53.2452,
  -53.2482,
  -53.2496,
  -53.2514,
  -53.2524,
  -53.2516,
  -53.2487,
  -53.2433,
  -53.2352,
  -53.2243,
  -53.2105,
  -53.1944,
  -53.1767,
  -53.1581,
  -53.1392,
  -53.1205,
  -53.1025,
  -53.0853,
  -53.0689,
  -53.0528,
  -53.0365,
  -53.0191,
  -52.9997,
  -52.978,
  -52.9537,
  -52.9266,
  -52.8971,
  -52.8654,
  -52.8317,
  -52.7965,
  -52.7602,
  -52.723,
  -52.6853,
  -52.646,
  -52.6071,
  -52.5675,
  -52.5276,
  -52.4875,
  -52.4472,
  -52.4067,
  -52.3658,
  -52.3243,
  -52.2824,
  -52.2402,
  -52.1977,
  -52.1549,
  -52.1118,
  -52.0688,
  -52.026,
  -51.9837,
  -51.942,
  -51.901,
  -51.8606,
  -51.8212,
  -51.7827,
  -51.745,
  -51.708,
  -51.6715,
  -51.6355,
  -51.5998,
  -51.5641,
  -51.5282,
  -51.4918,
  -51.4547,
  -51.4166,
  -51.3776,
  -51.3379,
  -51.2977,
  -51.2573,
  -51.2156,
  -51.1747,
  -51.1337,
  -51.0927,
  -51.0521,
  -51.0122,
  -50.9735,
  -50.9364,
  -50.9011,
  -50.8679,
  -50.8368,
  -50.8078,
  -50.7805,
  -50.7547,
  -50.7299,
  -50.7054,
  -50.6808,
  -50.6558,
  -50.6306,
  -50.6057,
  -50.5818,
  -50.5592,
  -50.5385,
  -50.5197,
  -50.5032,
  -50.4893,
  -50.4781,
  -50.4694,
  -50.463,
  -50.4585,
  -50.4555,
  -50.4534,
  -50.4516,
  -50.4494,
  -50.4466,
  -50.4437,
  -50.441,
  -48.3615,
  -48.4676,
  -48.5686,
  -48.6637,
  -48.7521,
  -48.8336,
  -48.9082,
  -48.976,
  -49.0375,
  -49.0932,
  -49.1438,
  -49.1899,
  -49.2321,
  -49.2706,
  -49.3046,
  -49.3361,
  -49.3639,
  -49.3883,
  -49.41,
  -49.4303,
  -49.4503,
  -49.471,
  -49.4933,
  -49.5169,
  -49.5423,
  -49.5687,
  -49.5961,
  -49.6239,
  -49.6514,
  -49.6781,
  -49.7023,
  -49.7264,
  -49.7497,
  -49.773,
  -49.7968,
  -49.8218,
  -49.8483,
  -49.8759,
  -49.9041,
  -49.9319,
  -49.9588,
  -49.9837,
  -50.0066,
  -50.0272,
  -50.0456,
  -50.0625,
  -50.0778,
  -50.0945,
  -50.1124,
  -50.1316,
  -50.1517,
  -50.1723,
  -50.1926,
  -50.2123,
  -50.2315,
  -50.2503,
  -50.2691,
  -50.2884,
  -50.3086,
  -50.3302,
  -50.3532,
  -50.3773,
  -50.4011,
  -50.426,
  -50.4505,
  -50.4736,
  -50.4945,
  -50.5126,
  -50.5275,
  -50.5395,
  -50.5492,
  -50.5573,
  -50.5642,
  -50.57,
  -50.5747,
  -50.5783,
  -50.5808,
  -50.5834,
  -50.5858,
  -50.5892,
  -50.5929,
  -50.5994,
  -50.6085,
  -50.6207,
  -50.6364,
  -50.6557,
  -50.6779,
  -50.7024,
  -50.7281,
  -50.7545,
  -50.7812,
  -50.808,
  -50.8351,
  -50.8626,
  -50.8905,
  -50.9189,
  -50.9474,
  -50.9762,
  -51.0038,
  -51.0323,
  -51.0603,
  -51.0883,
  -51.1161,
  -51.1439,
  -51.1714,
  -51.1983,
  -51.2245,
  -51.2499,
  -51.2747,
  -51.2992,
  -51.3232,
  -51.3473,
  -51.3722,
  -51.3985,
  -51.4261,
  -51.4548,
  -51.4837,
  -51.5124,
  -51.5397,
  -51.5672,
  -51.594,
  -51.6206,
  -51.6468,
  -51.6731,
  -51.7001,
  -51.7277,
  -51.7562,
  -51.7853,
  -51.8151,
  -51.8456,
  -51.8768,
  -51.9086,
  -51.9407,
  -51.9727,
  -52.0046,
  -52.0363,
  -52.0679,
  -52.0997,
  -52.1314,
  -52.1621,
  -52.1935,
  -52.2242,
  -52.254,
  -52.2831,
  -52.3112,
  -52.3386,
  -52.3658,
  -52.3927,
  -52.4198,
  -52.4473,
  -52.4757,
  -52.5049,
  -52.5352,
  -52.5661,
  -52.5976,
  -52.6296,
  -52.6626,
  -52.6969,
  -52.7329,
  -52.7698,
  -52.8068,
  -52.843,
  -52.8765,
  -52.9088,
  -52.939,
  -52.9675,
  -52.9951,
  -53.022,
  -53.0484,
  -53.0742,
  -53.099,
  -53.1227,
  -53.145,
  -53.1659,
  -53.1855,
  -53.2036,
  -53.2203,
  -53.2357,
  -53.2501,
  -53.2639,
  -53.2773,
  -53.2905,
  -53.3034,
  -53.3158,
  -53.3279,
  -53.3399,
  -53.3522,
  -53.3641,
  -53.3776,
  -53.3915,
  -53.4049,
  -53.4173,
  -53.4279,
  -53.4366,
  -53.4428,
  -53.4473,
  -53.4503,
  -53.4524,
  -53.4537,
  -53.4539,
  -53.4524,
  -53.4488,
  -53.4427,
  -53.4339,
  -53.4221,
  -53.4077,
  -53.3908,
  -53.3726,
  -53.3536,
  -53.3345,
  -53.3157,
  -53.2974,
  -53.2795,
  -53.2619,
  -53.2444,
  -53.2262,
  -53.2058,
  -53.1846,
  -53.1611,
  -53.1354,
  -53.1071,
  -53.0765,
  -53.0437,
  -53.009,
  -52.973,
  -52.9358,
  -52.8978,
  -52.859,
  -52.8195,
  -52.7791,
  -52.738,
  -52.6963,
  -52.6545,
  -52.6124,
  -52.5702,
  -52.5278,
  -52.4849,
  -52.4416,
  -52.3979,
  -52.3541,
  -52.3103,
  -52.2665,
  -52.2229,
  -52.1801,
  -52.138,
  -52.0968,
  -52.0563,
  -52.0164,
  -51.9772,
  -51.9387,
  -51.8995,
  -51.8615,
  -51.8237,
  -51.7856,
  -51.7475,
  -51.7092,
  -51.6706,
  -51.6316,
  -51.5921,
  -51.552,
  -51.5114,
  -51.4702,
  -51.4287,
  -51.387,
  -51.3449,
  -51.3025,
  -51.2599,
  -51.2173,
  -51.1751,
  -51.1339,
  -51.0937,
  -51.055,
  -51.0179,
  -50.9827,
  -50.9496,
  -50.9184,
  -50.889,
  -50.8611,
  -50.8341,
  -50.8074,
  -50.7804,
  -50.7529,
  -50.7251,
  -50.6977,
  -50.6715,
  -50.6471,
  -50.6251,
  -50.6056,
  -50.5888,
  -50.5751,
  -50.5644,
  -50.5564,
  -50.5509,
  -50.5462,
  -50.5439,
  -50.5424,
  -50.541,
  -50.5394,
  -50.5379,
  -50.5366,
  -50.5362,
  -48.3257,
  -48.4388,
  -48.546,
  -48.646,
  -48.7383,
  -48.8227,
  -48.8996,
  -48.9691,
  -49.0317,
  -49.0873,
  -49.1384,
  -49.1851,
  -49.2279,
  -49.2671,
  -49.303,
  -49.3358,
  -49.3658,
  -49.3931,
  -49.4184,
  -49.4428,
  -49.4674,
  -49.4932,
  -49.5204,
  -49.549,
  -49.5779,
  -49.6086,
  -49.6398,
  -49.6711,
  -49.7017,
  -49.7309,
  -49.7585,
  -49.7843,
  -49.8092,
  -49.8335,
  -49.8581,
  -49.8838,
  -49.9107,
  -49.9388,
  -49.9674,
  -49.996,
  -50.0227,
  -50.0487,
  -50.0726,
  -50.0939,
  -50.1129,
  -50.1303,
  -50.1469,
  -50.1638,
  -50.182,
  -50.2016,
  -50.2223,
  -50.2436,
  -50.2649,
  -50.2858,
  -50.3062,
  -50.326,
  -50.3448,
  -50.3649,
  -50.3858,
  -50.4078,
  -50.4312,
  -50.4556,
  -50.4809,
  -50.5066,
  -50.5318,
  -50.5561,
  -50.5787,
  -50.5986,
  -50.6158,
  -50.6304,
  -50.6427,
  -50.653,
  -50.6619,
  -50.6682,
  -50.674,
  -50.6783,
  -50.6814,
  -50.6838,
  -50.6861,
  -50.6893,
  -50.6939,
  -50.7004,
  -50.7099,
  -50.7228,
  -50.7396,
  -50.7601,
  -50.7835,
  -50.8089,
  -50.8355,
  -50.8626,
  -50.8899,
  -50.9162,
  -50.9436,
  -50.9713,
  -50.9996,
  -51.0283,
  -51.0571,
  -51.0863,
  -51.1157,
  -51.1453,
  -51.1749,
  -51.2049,
  -51.2351,
  -51.2653,
  -51.2951,
  -51.3241,
  -51.352,
  -51.3789,
  -51.4054,
  -51.4313,
  -51.4569,
  -51.4817,
  -51.5085,
  -51.5367,
  -51.5662,
  -51.5966,
  -51.6272,
  -51.6576,
  -51.6872,
  -51.7162,
  -51.7445,
  -51.7721,
  -51.7994,
  -51.826,
  -51.8531,
  -51.8807,
  -51.9091,
  -51.9378,
  -51.9678,
  -51.9986,
  -52.0307,
  -52.0628,
  -52.0965,
  -52.1304,
  -52.1644,
  -52.1983,
  -52.2321,
  -52.2661,
  -52.2999,
  -52.3338,
  -52.367,
  -52.3996,
  -52.4311,
  -52.4617,
  -52.4908,
  -52.5192,
  -52.5469,
  -52.5742,
  -52.6015,
  -52.6291,
  -52.6575,
  -52.6868,
  -52.7171,
  -52.7472,
  -52.7789,
  -52.8115,
  -52.8451,
  -52.8806,
  -52.9179,
  -52.9563,
  -52.9942,
  -53.0315,
  -53.0673,
  -53.1011,
  -53.1332,
  -53.1638,
  -53.1936,
  -53.2228,
  -53.2515,
  -53.2793,
  -53.3058,
  -53.3307,
  -53.3537,
  -53.3749,
  -53.3944,
  -53.4122,
  -53.4284,
  -53.4431,
  -53.4559,
  -53.4691,
  -53.4822,
  -53.495,
  -53.5076,
  -53.5199,
  -53.532,
  -53.544,
  -53.5564,
  -53.5694,
  -53.5831,
  -53.5971,
  -53.6109,
  -53.6238,
  -53.6352,
  -53.6446,
  -53.6517,
  -53.6568,
  -53.6601,
  -53.6623,
  -53.6632,
  -53.6629,
  -53.6606,
  -53.6562,
  -53.6492,
  -53.6397,
  -53.6273,
  -53.6112,
  -53.5939,
  -53.5752,
  -53.5559,
  -53.5367,
  -53.5176,
  -53.4986,
  -53.4798,
  -53.4608,
  -53.4416,
  -53.4215,
  -53.4001,
  -53.3769,
  -53.3517,
  -53.3247,
  -53.2951,
  -53.2636,
  -53.2297,
  -53.1942,
  -53.1576,
  -53.1197,
  -53.0808,
  -53.041,
  -53.0002,
  -52.9584,
  -52.9155,
  -52.8719,
  -52.8279,
  -52.7838,
  -52.7399,
  -52.696,
  -52.6516,
  -52.6058,
  -52.561,
  -52.5163,
  -52.4717,
  -52.4272,
  -52.3832,
  -52.3404,
  -52.2988,
  -52.258,
  -52.2179,
  -52.1782,
  -52.139,
  -52.1002,
  -52.0613,
  -52.022,
  -51.9823,
  -51.9421,
  -51.9015,
  -51.8607,
  -51.8193,
  -51.778,
  -51.7363,
  -51.6942,
  -51.652,
  -51.6094,
  -51.5666,
  -51.5235,
  -51.4802,
  -51.4365,
  -51.3925,
  -51.3486,
  -51.3053,
  -51.2629,
  -51.2215,
  -51.1813,
  -51.1427,
  -51.1057,
  -51.0706,
  -51.0373,
  -51.0046,
  -50.9742,
  -50.9446,
  -50.9153,
  -50.8857,
  -50.8556,
  -50.8254,
  -50.7957,
  -50.7676,
  -50.7418,
  -50.7187,
  -50.6985,
  -50.6813,
  -50.6673,
  -50.6564,
  -50.6482,
  -50.6425,
  -50.6386,
  -50.6358,
  -50.6339,
  -50.6325,
  -50.6312,
  -50.6306,
  -50.631,
  -50.6328,
  -48.287,
  -48.4079,
  -48.5218,
  -48.6275,
  -48.7234,
  -48.8113,
  -48.8904,
  -48.9614,
  -49.0248,
  -49.0816,
  -49.1323,
  -49.1781,
  -49.22,
  -49.2586,
  -49.2945,
  -49.328,
  -49.3598,
  -49.3901,
  -49.4197,
  -49.4483,
  -49.4787,
  -49.5106,
  -49.5439,
  -49.5784,
  -49.6134,
  -49.6489,
  -49.6845,
  -49.7195,
  -49.7534,
  -49.7856,
  -49.8158,
  -49.8441,
  -49.8709,
  -49.8968,
  -49.9218,
  -49.9483,
  -49.9756,
  -50.0042,
  -50.0333,
  -50.0628,
  -50.0914,
  -50.1184,
  -50.1433,
  -50.1656,
  -50.1851,
  -50.203,
  -50.2202,
  -50.2375,
  -50.256,
  -50.2758,
  -50.2958,
  -50.3176,
  -50.3395,
  -50.3613,
  -50.3826,
  -50.4035,
  -50.4242,
  -50.4452,
  -50.4669,
  -50.4896,
  -50.5136,
  -50.5386,
  -50.5644,
  -50.5907,
  -50.6168,
  -50.6421,
  -50.666,
  -50.6866,
  -50.706,
  -50.7231,
  -50.738,
  -50.7509,
  -50.762,
  -50.7712,
  -50.7787,
  -50.7843,
  -50.7883,
  -50.7913,
  -50.7939,
  -50.7969,
  -50.8013,
  -50.8077,
  -50.8174,
  -50.8308,
  -50.8484,
  -50.8686,
  -50.8927,
  -50.9187,
  -50.9457,
  -50.9733,
  -51.0009,
  -51.0287,
  -51.0565,
  -51.0846,
  -51.1133,
  -51.1423,
  -51.1718,
  -51.2015,
  -51.2317,
  -51.2625,
  -51.2937,
  -51.3255,
  -51.3578,
  -51.389,
  -51.4208,
  -51.4516,
  -51.481,
  -51.5094,
  -51.5372,
  -51.5648,
  -51.5922,
  -51.6202,
  -51.6493,
  -51.6797,
  -51.7116,
  -51.7441,
  -51.7766,
  -51.8088,
  -51.8403,
  -51.8712,
  -51.9011,
  -51.9301,
  -51.9583,
  -51.9847,
  -52.0122,
  -52.0391,
  -52.0667,
  -52.0951,
  -52.1249,
  -52.1559,
  -52.1887,
  -52.2225,
  -52.2575,
  -52.2929,
  -52.3286,
  -52.3645,
  -52.4005,
  -52.4366,
  -52.4728,
  -52.5087,
  -52.5441,
  -52.5787,
  -52.6119,
  -52.6439,
  -52.6746,
  -52.7031,
  -52.7314,
  -52.7593,
  -52.7869,
  -52.8146,
  -52.8431,
  -52.8726,
  -52.9031,
  -52.9344,
  -52.9665,
  -52.9998,
  -53.0345,
  -53.0712,
  -53.1095,
  -53.1487,
  -53.1878,
  -53.2258,
  -53.2625,
  -53.2976,
  -53.3314,
  -53.364,
  -53.396,
  -53.4276,
  -53.4576,
  -53.4875,
  -53.516,
  -53.5424,
  -53.5667,
  -53.5886,
  -53.6085,
  -53.6263,
  -53.6424,
  -53.6569,
  -53.6703,
  -53.6833,
  -53.6961,
  -53.709,
  -53.7214,
  -53.7334,
  -53.7454,
  -53.7574,
  -53.7698,
  -53.7828,
  -53.7964,
  -53.8104,
  -53.8242,
  -53.8374,
  -53.8494,
  -53.8596,
  -53.8677,
  -53.8726,
  -53.8765,
  -53.8787,
  -53.8794,
  -53.8783,
  -53.8752,
  -53.8698,
  -53.8621,
  -53.8517,
  -53.8389,
  -53.8235,
  -53.806,
  -53.787,
  -53.7676,
  -53.7481,
  -53.7284,
  -53.7086,
  -53.6886,
  -53.668,
  -53.6468,
  -53.6247,
  -53.6012,
  -53.5763,
  -53.5496,
  -53.5212,
  -53.4906,
  -53.4579,
  -53.4232,
  -53.3869,
  -53.3485,
  -53.3099,
  -53.2703,
  -53.2294,
  -53.1872,
  -53.1438,
  -53.099,
  -53.0533,
  -53.0073,
  -52.9612,
  -52.9154,
  -52.8695,
  -52.8238,
  -52.7779,
  -52.7322,
  -52.6866,
  -52.6413,
  -52.5963,
  -52.5524,
  -52.5095,
  -52.468,
  -52.4276,
  -52.3879,
  -52.3483,
  -52.3088,
  -52.2693,
  -52.2291,
  -52.1881,
  -52.1462,
  -52.1036,
  -52.0606,
  -52.0172,
  -51.9735,
  -51.9299,
  -51.8861,
  -51.8426,
  -51.7978,
  -51.7538,
  -51.7096,
  -51.6651,
  -51.6207,
  -51.5758,
  -51.5305,
  -51.4855,
  -51.4411,
  -51.3977,
  -51.3554,
  -51.3141,
  -51.2742,
  -51.2356,
  -51.1987,
  -51.1632,
  -51.1291,
  -51.0962,
  -51.0638,
  -51.0317,
  -50.9996,
  -50.967,
  -50.9348,
  -50.9032,
  -50.8736,
  -50.8465,
  -50.8225,
  -50.8017,
  -50.784,
  -50.7694,
  -50.7577,
  -50.7486,
  -50.7416,
  -50.7364,
  -50.7324,
  -50.7293,
  -50.727,
  -50.7256,
  -50.7254,
  -50.7272,
  -50.7311,
  -48.2443,
  -48.3744,
  -48.4957,
  -48.6076,
  -48.7093,
  -48.8008,
  -48.8824,
  -48.9546,
  -49.0179,
  -49.0737,
  -49.1225,
  -49.1661,
  -49.2055,
  -49.2412,
  -49.2759,
  -49.3095,
  -49.3428,
  -49.3765,
  -49.4112,
  -49.4472,
  -49.4849,
  -49.5242,
  -49.5651,
  -49.6063,
  -49.6477,
  -49.6888,
  -49.7289,
  -49.7679,
  -49.8043,
  -49.8398,
  -49.8731,
  -49.9042,
  -49.9335,
  -49.9617,
  -49.9893,
  -50.0171,
  -50.0453,
  -50.0746,
  -50.1043,
  -50.1345,
  -50.164,
  -50.192,
  -50.218,
  -50.2411,
  -50.2607,
  -50.2792,
  -50.2968,
  -50.315,
  -50.3338,
  -50.3538,
  -50.3749,
  -50.3968,
  -50.4192,
  -50.4415,
  -50.4635,
  -50.4855,
  -50.5072,
  -50.5292,
  -50.5518,
  -50.5754,
  -50.6,
  -50.6247,
  -50.6511,
  -50.6778,
  -50.7043,
  -50.7304,
  -50.7552,
  -50.7782,
  -50.7994,
  -50.8189,
  -50.8365,
  -50.8521,
  -50.8658,
  -50.8773,
  -50.8869,
  -50.8944,
  -50.9002,
  -50.9044,
  -50.9068,
  -50.91,
  -50.9144,
  -50.9209,
  -50.9306,
  -50.9444,
  -50.9622,
  -50.9837,
  -51.008,
  -51.034,
  -51.061,
  -51.0884,
  -51.1161,
  -51.1441,
  -51.1723,
  -51.201,
  -51.2302,
  -51.2599,
  -51.2892,
  -51.3199,
  -51.3514,
  -51.3834,
  -51.4161,
  -51.4498,
  -51.484,
  -51.5182,
  -51.5516,
  -51.5839,
  -51.615,
  -51.6451,
  -51.6745,
  -51.7037,
  -51.7331,
  -51.7634,
  -51.795,
  -51.8281,
  -51.8623,
  -51.8972,
  -51.9309,
  -51.9652,
  -51.9987,
  -52.0315,
  -52.0632,
  -52.0937,
  -52.1231,
  -52.1511,
  -52.1779,
  -52.205,
  -52.2319,
  -52.2597,
  -52.2888,
  -52.3199,
  -52.3529,
  -52.3876,
  -52.4235,
  -52.4601,
  -52.4972,
  -52.5347,
  -52.5727,
  -52.6099,
  -52.6483,
  -52.6864,
  -52.7238,
  -52.7604,
  -52.7954,
  -52.8289,
  -52.8608,
  -52.8913,
  -52.9208,
  -52.9494,
  -52.9776,
  -53.0058,
  -53.0346,
  -53.0642,
  -53.095,
  -53.1268,
  -53.1596,
  -53.1937,
  -53.2296,
  -53.2674,
  -53.3069,
  -53.3468,
  -53.3853,
  -53.4238,
  -53.4612,
  -53.4975,
  -53.5329,
  -53.5675,
  -53.6016,
  -53.6353,
  -53.6686,
  -53.7007,
  -53.7312,
  -53.7597,
  -53.7856,
  -53.8086,
  -53.8288,
  -53.8474,
  -53.8635,
  -53.878,
  -53.8914,
  -53.9046,
  -53.9178,
  -53.9308,
  -53.9434,
  -53.9556,
  -53.9676,
  -53.9788,
  -53.9911,
  -54.004,
  -54.0174,
  -54.0309,
  -54.0446,
  -54.0579,
  -54.0703,
  -54.0812,
  -54.0902,
  -54.097,
  -54.1015,
  -54.1038,
  -54.1038,
  -54.1017,
  -54.0974,
  -54.0912,
  -54.0826,
  -54.0718,
  -54.0587,
  -54.0433,
  -54.026,
  -54.0073,
  -53.9877,
  -53.9677,
  -53.9474,
  -53.9266,
  -53.9051,
  -53.8818,
  -53.8586,
  -53.8343,
  -53.8089,
  -53.7822,
  -53.7541,
  -53.7244,
  -53.6928,
  -53.6591,
  -53.6233,
  -53.5858,
  -53.5474,
  -53.508,
  -53.4676,
  -53.4259,
  -53.3825,
  -53.3374,
  -53.2909,
  -53.2432,
  -53.1952,
  -53.1471,
  -53.0992,
  -53.0516,
  -53.0044,
  -52.9575,
  -52.9108,
  -52.8646,
  -52.8189,
  -52.7737,
  -52.7294,
  -52.6865,
  -52.645,
  -52.6049,
  -52.5643,
  -52.5244,
  -52.4843,
  -52.4435,
  -52.4017,
  -52.3585,
  -52.3142,
  -52.2691,
  -52.2235,
  -52.1778,
  -52.1322,
  -52.087,
  -52.0416,
  -51.9966,
  -51.9513,
  -51.9059,
  -51.8602,
  -51.8144,
  -51.7685,
  -51.7223,
  -51.676,
  -51.6299,
  -51.5845,
  -51.5402,
  -51.4972,
  -51.4553,
  -51.4144,
  -51.3746,
  -51.336,
  -51.2986,
  -51.2622,
  -51.2264,
  -51.1912,
  -51.1562,
  -51.1212,
  -51.0863,
  -51.0523,
  -51.0193,
  -50.9887,
  -50.9608,
  -50.936,
  -50.9146,
  -50.8953,
  -50.8798,
  -50.8669,
  -50.8563,
  -50.8477,
  -50.8405,
  -50.8345,
  -50.8296,
  -50.8258,
  -50.8236,
  -50.8237,
  -50.8265,
  -50.8318,
  -48.2011,
  -48.3407,
  -48.47,
  -48.5886,
  -48.6954,
  -48.7904,
  -48.8742,
  -48.947,
  -49.0083,
  -49.0617,
  -49.107,
  -49.1462,
  -49.1814,
  -49.2143,
  -49.2466,
  -49.2797,
  -49.3146,
  -49.3523,
  -49.3932,
  -49.4373,
  -49.4842,
  -49.5331,
  -49.5827,
  -49.6317,
  -49.6802,
  -49.7273,
  -49.7725,
  -49.8157,
  -49.8567,
  -49.8955,
  -49.9319,
  -49.9662,
  -49.9986,
  -50.0295,
  -50.0594,
  -50.0892,
  -50.119,
  -50.1491,
  -50.1786,
  -50.2093,
  -50.2395,
  -50.2683,
  -50.2949,
  -50.3192,
  -50.3412,
  -50.3608,
  -50.3796,
  -50.3985,
  -50.4179,
  -50.4382,
  -50.4594,
  -50.4815,
  -50.5039,
  -50.5267,
  -50.5494,
  -50.5711,
  -50.5939,
  -50.617,
  -50.6406,
  -50.6649,
  -50.69,
  -50.716,
  -50.7425,
  -50.7694,
  -50.7961,
  -50.8224,
  -50.8478,
  -50.8721,
  -50.8952,
  -50.9169,
  -50.9371,
  -50.9556,
  -50.9712,
  -50.9854,
  -50.9976,
  -51.0075,
  -51.0153,
  -51.0212,
  -51.0259,
  -51.0301,
  -51.035,
  -51.0421,
  -51.0522,
  -51.0661,
  -51.0839,
  -51.105,
  -51.1288,
  -51.1542,
  -51.1804,
  -51.2071,
  -51.2334,
  -51.2612,
  -51.2896,
  -51.3188,
  -51.3488,
  -51.3797,
  -51.4114,
  -51.4437,
  -51.4766,
  -51.5102,
  -51.5447,
  -51.5802,
  -51.6163,
  -51.6523,
  -51.6875,
  -51.7216,
  -51.7546,
  -51.7866,
  -51.8178,
  -51.8478,
  -51.8791,
  -51.9116,
  -51.9456,
  -51.9812,
  -52.018,
  -52.0553,
  -52.0924,
  -52.1291,
  -52.1648,
  -52.1994,
  -52.2326,
  -52.2643,
  -52.2943,
  -52.3227,
  -52.3497,
  -52.3762,
  -52.4027,
  -52.4299,
  -52.4588,
  -52.4889,
  -52.5223,
  -52.5577,
  -52.5945,
  -52.6322,
  -52.6705,
  -52.7094,
  -52.7488,
  -52.7886,
  -52.8287,
  -52.8683,
  -52.9074,
  -52.9456,
  -52.9823,
  -53.0172,
  -53.0507,
  -53.0828,
  -53.1136,
  -53.1434,
  -53.1726,
  -53.2016,
  -53.2308,
  -53.26,
  -53.2912,
  -53.3236,
  -53.3573,
  -53.3922,
  -53.429,
  -53.4677,
  -53.508,
  -53.5486,
  -53.5887,
  -53.6278,
  -53.6663,
  -53.7038,
  -53.7407,
  -53.777,
  -53.8129,
  -53.8484,
  -53.8836,
  -53.9177,
  -53.9501,
  -53.9802,
  -54.0077,
  -54.0318,
  -54.0534,
  -54.0711,
  -54.088,
  -54.103,
  -54.1172,
  -54.1311,
  -54.145,
  -54.1588,
  -54.1722,
  -54.185,
  -54.1975,
  -54.2098,
  -54.2223,
  -54.2351,
  -54.2482,
  -54.2614,
  -54.2749,
  -54.2883,
  -54.3012,
  -54.3128,
  -54.3224,
  -54.3297,
  -54.3345,
  -54.3364,
  -54.3357,
  -54.3325,
  -54.3269,
  -54.3194,
  -54.3089,
  -54.2976,
  -54.2846,
  -54.2693,
  -54.2523,
  -54.2339,
  -54.2145,
  -54.1942,
  -54.1732,
  -54.1514,
  -54.1286,
  -54.1046,
  -54.0793,
  -54.0528,
  -54.0251,
  -53.9965,
  -53.9667,
  -53.9355,
  -53.9026,
  -53.8679,
  -53.8313,
  -53.793,
  -53.7536,
  -53.7133,
  -53.6721,
  -53.6295,
  -53.585,
  -53.5385,
  -53.4903,
  -53.4409,
  -53.391,
  -53.3399,
  -53.29,
  -53.2408,
  -53.1922,
  -53.1442,
  -53.097,
  -53.0504,
  -53.0045,
  -52.9593,
  -52.915,
  -52.872,
  -52.8301,
  -52.7896,
  -52.7494,
  -52.7089,
  -52.6677,
  -52.6252,
  -52.5813,
  -52.5361,
  -52.4897,
  -52.4424,
  -52.3945,
  -52.3467,
  -52.2995,
  -52.2527,
  -52.206,
  -52.1592,
  -52.1123,
  -52.0653,
  -52.0181,
  -51.9708,
  -51.9234,
  -51.8761,
  -51.8287,
  -51.7817,
  -51.7356,
  -51.6906,
  -51.6468,
  -51.6032,
  -51.5615,
  -51.5206,
  -51.4803,
  -51.4407,
  -51.4019,
  -51.3633,
  -51.3249,
  -51.287,
  -51.2495,
  -51.2127,
  -51.1771,
  -51.1433,
  -51.1119,
  -51.0835,
  -51.0584,
  -51.0365,
  -51.0176,
  -51.0011,
  -50.9869,
  -50.9747,
  -50.964,
  -50.9544,
  -50.946,
  -50.9388,
  -50.9333,
  -50.93,
  -50.9296,
  -50.9326,
  -50.9386,
  -48.1598,
  -48.3086,
  -48.4447,
  -48.569,
  -48.6803,
  -48.7781,
  -48.8629,
  -48.9351,
  -48.9952,
  -49.0445,
  -49.0846,
  -49.1177,
  -49.1468,
  -49.1745,
  -49.2033,
  -49.2354,
  -49.2724,
  -49.314,
  -49.3627,
  -49.4168,
  -49.475,
  -49.5354,
  -49.5962,
  -49.6559,
  -49.7129,
  -49.7667,
  -49.8173,
  -49.8647,
  -49.9094,
  -49.9515,
  -49.9911,
  -50.0287,
  -50.0635,
  -50.0978,
  -50.1309,
  -50.1631,
  -50.1948,
  -50.2264,
  -50.2579,
  -50.2891,
  -50.3197,
  -50.3492,
  -50.3768,
  -50.4023,
  -50.4255,
  -50.4469,
  -50.4672,
  -50.4874,
  -50.5066,
  -50.5272,
  -50.5485,
  -50.5706,
  -50.5933,
  -50.6165,
  -50.6398,
  -50.6633,
  -50.6869,
  -50.711,
  -50.7354,
  -50.7603,
  -50.7857,
  -50.8117,
  -50.838,
  -50.8646,
  -50.8912,
  -50.9166,
  -50.9426,
  -50.9679,
  -50.9927,
  -51.0166,
  -51.0393,
  -51.0606,
  -51.0801,
  -51.0974,
  -51.1123,
  -51.1248,
  -51.1351,
  -51.1433,
  -51.1499,
  -51.1558,
  -51.1621,
  -51.1701,
  -51.1809,
  -51.194,
  -51.2115,
  -51.2319,
  -51.2545,
  -51.2785,
  -51.3034,
  -51.329,
  -51.3553,
  -51.3826,
  -51.4111,
  -51.4408,
  -51.4719,
  -51.5042,
  -51.5376,
  -51.5718,
  -51.6068,
  -51.6423,
  -51.6786,
  -51.716,
  -51.753,
  -51.791,
  -51.8281,
  -51.8642,
  -51.8992,
  -51.9332,
  -51.9665,
  -51.9994,
  -52.0328,
  -52.0674,
  -52.1039,
  -52.1421,
  -52.1814,
  -52.2213,
  -52.261,
  -52.3001,
  -52.3381,
  -52.3744,
  -52.409,
  -52.4405,
  -52.4709,
  -52.4992,
  -52.5263,
  -52.5527,
  -52.579,
  -52.6062,
  -52.6351,
  -52.6664,
  -52.7002,
  -52.7362,
  -52.7738,
  -52.8123,
  -52.8515,
  -52.8913,
  -52.9317,
  -52.9725,
  -53.0135,
  -53.0543,
  -53.0946,
  -53.134,
  -53.1722,
  -53.2078,
  -53.243,
  -53.2768,
  -53.3093,
  -53.3407,
  -53.3712,
  -53.4013,
  -53.4314,
  -53.4622,
  -53.4942,
  -53.5275,
  -53.5621,
  -53.5981,
  -53.6359,
  -53.6752,
  -53.7159,
  -53.7569,
  -53.7975,
  -53.8373,
  -53.8766,
  -53.9153,
  -53.9535,
  -53.9912,
  -54.0276,
  -54.0648,
  -54.1015,
  -54.1373,
  -54.1713,
  -54.203,
  -54.2318,
  -54.2575,
  -54.28,
  -54.2999,
  -54.3178,
  -54.334,
  -54.3495,
  -54.3646,
  -54.3797,
  -54.3947,
  -54.4094,
  -54.4234,
  -54.4368,
  -54.4499,
  -54.4627,
  -54.4756,
  -54.4884,
  -54.5015,
  -54.515,
  -54.5284,
  -54.5405,
  -54.5526,
  -54.5627,
  -54.57,
  -54.5744,
  -54.5756,
  -54.5736,
  -54.5687,
  -54.5618,
  -54.5531,
  -54.5428,
  -54.5314,
  -54.5183,
  -54.5034,
  -54.4869,
  -54.469,
  -54.4498,
  -54.4293,
  -54.4077,
  -54.3849,
  -54.3608,
  -54.3354,
  -54.3083,
  -54.2797,
  -54.2499,
  -54.2192,
  -54.1876,
  -54.1549,
  -54.1207,
  -54.0839,
  -54.0462,
  -54.007,
  -53.9664,
  -53.9251,
  -53.883,
  -53.8395,
  -53.7941,
  -53.7463,
  -53.6967,
  -53.6457,
  -53.594,
  -53.5421,
  -53.4907,
  -53.4397,
  -53.3897,
  -53.3407,
  -53.2928,
  -53.246,
  -53.2001,
  -53.155,
  -53.1107,
  -53.0674,
  -53.0251,
  -52.9835,
  -52.9422,
  -52.9004,
  -52.8574,
  -52.813,
  -52.7669,
  -52.7193,
  -52.6709,
  -52.6217,
  -52.5724,
  -52.5233,
  -52.4735,
  -52.4252,
  -52.3771,
  -52.3287,
  -52.2801,
  -52.2313,
  -52.1823,
  -52.1334,
  -52.0846,
  -52.036,
  -51.9877,
  -51.94,
  -51.8933,
  -51.8478,
  -51.8034,
  -51.7603,
  -51.7178,
  -51.6759,
  -51.6343,
  -51.5925,
  -51.5509,
  -51.5097,
  -51.4683,
  -51.4276,
  -51.3877,
  -51.3491,
  -51.3123,
  -51.2778,
  -51.246,
  -51.2174,
  -51.192,
  -51.1696,
  -51.1497,
  -51.1324,
  -51.1168,
  -51.1028,
  -51.0899,
  -51.078,
  -51.067,
  -51.0574,
  -51.0499,
  -51.0453,
  -51.0442,
  -51.0467,
  -51.0527,
  -48.1242,
  -48.2801,
  -48.4233,
  -48.5522,
  -48.6661,
  -48.765,
  -48.8491,
  -48.9188,
  -48.9748,
  -49.0184,
  -49.0516,
  -49.0771,
  -49.0976,
  -49.1188,
  -49.1434,
  -49.1745,
  -49.2143,
  -49.2634,
  -49.3218,
  -49.3881,
  -49.4597,
  -49.5338,
  -49.6074,
  -49.6782,
  -49.7447,
  -49.8061,
  -49.8623,
  -49.9132,
  -49.9614,
  -50.0065,
  -50.0493,
  -50.0903,
  -50.1299,
  -50.168,
  -50.2047,
  -50.2402,
  -50.2744,
  -50.3078,
  -50.3405,
  -50.3725,
  -50.4035,
  -50.4335,
  -50.462,
  -50.4879,
  -50.5129,
  -50.5362,
  -50.5584,
  -50.58,
  -50.6013,
  -50.6227,
  -50.6444,
  -50.6667,
  -50.6898,
  -50.7134,
  -50.7372,
  -50.7614,
  -50.7858,
  -50.8104,
  -50.8355,
  -50.8598,
  -50.8852,
  -50.9109,
  -50.9369,
  -50.9631,
  -50.9893,
  -51.0159,
  -51.0423,
  -51.0687,
  -51.0949,
  -51.1207,
  -51.1457,
  -51.1696,
  -51.1919,
  -51.212,
  -51.2299,
  -51.2453,
  -51.2571,
  -51.268,
  -51.2771,
  -51.2853,
  -51.2937,
  -51.3034,
  -51.3152,
  -51.3297,
  -51.3468,
  -51.3661,
  -51.3871,
  -51.4093,
  -51.4325,
  -51.4567,
  -51.4819,
  -51.5086,
  -51.5368,
  -51.5671,
  -51.5992,
  -51.6319,
  -51.6671,
  -51.7034,
  -51.7405,
  -51.7783,
  -51.8169,
  -51.8563,
  -51.8963,
  -51.9362,
  -51.9755,
  -52.0139,
  -52.0512,
  -52.0874,
  -52.1228,
  -52.1579,
  -52.1934,
  -52.2303,
  -52.2693,
  -52.3101,
  -52.3512,
  -52.3936,
  -52.4359,
  -52.4774,
  -52.5174,
  -52.5554,
  -52.5908,
  -52.6239,
  -52.6545,
  -52.6832,
  -52.7104,
  -52.7369,
  -52.7632,
  -52.7909,
  -52.8203,
  -52.8522,
  -52.8866,
  -52.9231,
  -52.9611,
  -53.0001,
  -53.0398,
  -53.079,
  -53.1197,
  -53.1608,
  -53.2022,
  -53.2436,
  -53.2845,
  -53.3251,
  -53.3647,
  -53.4029,
  -53.4399,
  -53.4756,
  -53.5101,
  -53.5433,
  -53.5754,
  -53.6068,
  -53.6382,
  -53.6702,
  -53.7033,
  -53.7379,
  -53.7736,
  -53.8107,
  -53.8493,
  -53.8882,
  -53.929,
  -53.9702,
  -54.0111,
  -54.0516,
  -54.0917,
  -54.1314,
  -54.1707,
  -54.2096,
  -54.2482,
  -54.2865,
  -54.3243,
  -54.3612,
  -54.3965,
  -54.4295,
  -54.4595,
  -54.4865,
  -54.5105,
  -54.532,
  -54.5513,
  -54.5693,
  -54.5866,
  -54.6035,
  -54.6203,
  -54.637,
  -54.6523,
  -54.668,
  -54.683,
  -54.6972,
  -54.711,
  -54.7245,
  -54.7371,
  -54.7503,
  -54.7641,
  -54.7774,
  -54.7905,
  -54.8024,
  -54.8124,
  -54.8196,
  -54.8232,
  -54.8231,
  -54.8196,
  -54.8132,
  -54.8046,
  -54.7944,
  -54.7835,
  -54.7716,
  -54.7585,
  -54.7442,
  -54.7283,
  -54.7108,
  -54.6919,
  -54.6714,
  -54.6483,
  -54.6248,
  -54.5998,
  -54.5731,
  -54.5446,
  -54.5144,
  -54.4828,
  -54.45,
  -54.4165,
  -54.3821,
  -54.3463,
  -54.3093,
  -54.2706,
  -54.2304,
  -54.189,
  -54.1467,
  -54.1033,
  -54.0584,
  -54.0119,
  -53.963,
  -53.9121,
  -53.8599,
  -53.8068,
  -53.7535,
  -53.7006,
  -53.6482,
  -53.5967,
  -53.5467,
  -53.4982,
  -53.4511,
  -53.4051,
  -53.3601,
  -53.3158,
  -53.271,
  -53.2277,
  -53.1848,
  -53.1417,
  -53.0979,
  -53.0527,
  -53.0059,
  -52.9575,
  -52.9079,
  -52.8576,
  -52.8069,
  -52.7563,
  -52.706,
  -52.6561,
  -52.6065,
  -52.5569,
  -52.507,
  -52.4567,
  -52.4061,
  -52.3554,
  -52.3049,
  -52.2546,
  -52.2048,
  -52.1557,
  -52.1075,
  -52.0604,
  -52.0145,
  -51.9697,
  -51.9259,
  -51.8826,
  -51.8396,
  -51.7964,
  -51.7526,
  -51.7086,
  -51.6645,
  -51.6206,
  -51.5773,
  -51.5353,
  -51.4951,
  -51.4573,
  -51.4213,
  -51.3893,
  -51.3604,
  -51.3346,
  -51.3115,
  -51.2912,
  -51.2726,
  -51.2557,
  -51.2397,
  -51.2247,
  -51.2104,
  -51.1969,
  -51.185,
  -51.1757,
  -51.1697,
  -51.1676,
  -51.1694,
  -51.1747,
  -48.1009,
  -48.2606,
  -48.4067,
  -48.5373,
  -48.6514,
  -48.749,
  -48.8293,
  -48.8944,
  -48.9442,
  -48.9801,
  -49.0047,
  -49.0212,
  -49.034,
  -49.0485,
  -49.0688,
  -49.0995,
  -49.143,
  -49.2005,
  -49.2706,
  -49.3511,
  -49.4385,
  -49.5272,
  -49.6151,
  -49.6984,
  -49.7751,
  -49.8445,
  -49.9069,
  -49.9632,
  -50.0148,
  -50.063,
  -50.1089,
  -50.1532,
  -50.1966,
  -50.2388,
  -50.2796,
  -50.3188,
  -50.3562,
  -50.3909,
  -50.4251,
  -50.4577,
  -50.4893,
  -50.5199,
  -50.5494,
  -50.5777,
  -50.6048,
  -50.6304,
  -50.6549,
  -50.6783,
  -50.7011,
  -50.7234,
  -50.746,
  -50.7688,
  -50.7924,
  -50.8154,
  -50.8398,
  -50.8644,
  -50.8894,
  -50.9146,
  -50.9398,
  -50.9652,
  -50.9905,
  -51.016,
  -51.0417,
  -51.0674,
  -51.0936,
  -51.1202,
  -51.1472,
  -51.1745,
  -51.2019,
  -51.2291,
  -51.255,
  -51.2811,
  -51.3057,
  -51.3285,
  -51.3492,
  -51.3674,
  -51.3831,
  -51.3967,
  -51.4088,
  -51.4198,
  -51.4309,
  -51.4429,
  -51.4562,
  -51.4715,
  -51.4884,
  -51.5067,
  -51.526,
  -51.5463,
  -51.5667,
  -51.5893,
  -51.6134,
  -51.6393,
  -51.6673,
  -51.6979,
  -51.7306,
  -51.7657,
  -51.8026,
  -51.8409,
  -51.8801,
  -51.9202,
  -51.9611,
  -52.0025,
  -52.0446,
  -52.0866,
  -52.1283,
  -52.1693,
  -52.2092,
  -52.247,
  -52.2848,
  -52.3222,
  -52.3601,
  -52.3995,
  -52.441,
  -52.4844,
  -52.5291,
  -52.5743,
  -52.619,
  -52.6626,
  -52.7043,
  -52.7436,
  -52.78,
  -52.8136,
  -52.8441,
  -52.8729,
  -52.9006,
  -52.9277,
  -52.9553,
  -52.9825,
  -53.0128,
  -53.0456,
  -53.0806,
  -53.1175,
  -53.1557,
  -53.1949,
  -53.2347,
  -53.2748,
  -53.3153,
  -53.3562,
  -53.3975,
  -53.4389,
  -53.4804,
  -53.5216,
  -53.5625,
  -53.6023,
  -53.6411,
  -53.6788,
  -53.7152,
  -53.7502,
  -53.784,
  -53.8161,
  -53.849,
  -53.8826,
  -53.9172,
  -53.9532,
  -53.9905,
  -54.0289,
  -54.0683,
  -54.1086,
  -54.1494,
  -54.1906,
  -54.232,
  -54.273,
  -54.3138,
  -54.3544,
  -54.3946,
  -54.4343,
  -54.4737,
  -54.5127,
  -54.5511,
  -54.5887,
  -54.6248,
  -54.6586,
  -54.6898,
  -54.7173,
  -54.743,
  -54.7665,
  -54.788,
  -54.8082,
  -54.8276,
  -54.8467,
  -54.8655,
  -54.8842,
  -54.9024,
  -54.92,
  -54.9368,
  -54.9527,
  -54.9678,
  -54.9818,
  -54.9953,
  -55.009,
  -55.0229,
  -55.0363,
  -55.0491,
  -55.0609,
  -55.0703,
  -55.0766,
  -55.079,
  -55.0774,
  -55.0723,
  -55.0632,
  -55.0532,
  -55.0421,
  -55.0302,
  -55.0178,
  -55.0048,
  -54.9909,
  -54.9757,
  -54.9587,
  -54.9399,
  -54.9194,
  -54.8969,
  -54.8727,
  -54.847,
  -54.8195,
  -54.7901,
  -54.7588,
  -54.7258,
  -54.6914,
  -54.6559,
  -54.6196,
  -54.5821,
  -54.5438,
  -54.5039,
  -54.4629,
  -54.4207,
  -54.3773,
  -54.3325,
  -54.2862,
  -54.2383,
  -54.1882,
  -54.1353,
  -54.0822,
  -54.0281,
  -53.9736,
  -53.9194,
  -53.8657,
  -53.8131,
  -53.7619,
  -53.7125,
  -53.6648,
  -53.6186,
  -53.5732,
  -53.5286,
  -53.4842,
  -53.4396,
  -53.3949,
  -53.3495,
  -53.3032,
  -53.2555,
  -53.2064,
  -53.1558,
  -53.1042,
  -53.0524,
  -53.0003,
  -52.9486,
  -52.8975,
  -52.8465,
  -52.7956,
  -52.7445,
  -52.693,
  -52.6411,
  -52.5891,
  -52.5367,
  -52.4845,
  -52.4329,
  -52.3821,
  -52.3323,
  -52.2827,
  -52.2352,
  -52.189,
  -52.1437,
  -52.0991,
  -52.0548,
  -52.0105,
  -51.9656,
  -51.9199,
  -51.8736,
  -51.8271,
  -51.781,
  -51.7357,
  -51.692,
  -51.6505,
  -51.6117,
  -51.576,
  -51.5435,
  -51.5142,
  -51.488,
  -51.4645,
  -51.4431,
  -51.4235,
  -51.4051,
  -51.3874,
  -51.3701,
  -51.3534,
  -51.3376,
  -51.3238,
  -51.3129,
  -51.3057,
  -51.3025,
  -51.3033,
  -51.3074,
  -48.0924,
  -48.2503,
  -48.3948,
  -48.5233,
  -48.6344,
  -48.7275,
  -48.803,
  -48.8613,
  -48.9027,
  -48.9293,
  -48.9437,
  -48.9503,
  -48.9547,
  -48.9625,
  -48.9798,
  -49.0116,
  -49.0599,
  -49.1274,
  -49.2113,
  -49.3083,
  -49.4129,
  -49.5193,
  -49.6227,
  -49.7191,
  -49.8065,
  -49.8842,
  -49.9528,
  -50.0139,
  -50.0689,
  -50.1201,
  -50.169,
  -50.2159,
  -50.263,
  -50.3095,
  -50.3546,
  -50.3977,
  -50.4385,
  -50.4769,
  -50.5128,
  -50.5469,
  -50.5793,
  -50.6107,
  -50.6413,
  -50.6712,
  -50.7003,
  -50.7283,
  -50.7552,
  -50.7798,
  -50.8044,
  -50.8283,
  -50.852,
  -50.876,
  -50.9001,
  -50.9245,
  -50.9493,
  -50.9744,
  -50.9995,
  -51.0249,
  -51.0502,
  -51.0756,
  -51.101,
  -51.1265,
  -51.152,
  -51.1777,
  -51.2029,
  -51.2296,
  -51.257,
  -51.2848,
  -51.313,
  -51.3412,
  -51.3694,
  -51.3971,
  -51.4236,
  -51.4487,
  -51.4717,
  -51.4928,
  -51.5115,
  -51.5281,
  -51.5434,
  -51.5578,
  -51.5719,
  -51.5856,
  -51.6009,
  -51.6172,
  -51.6342,
  -51.6519,
  -51.6701,
  -51.6889,
  -51.7087,
  -51.73,
  -51.7532,
  -51.7785,
  -51.8064,
  -51.8369,
  -51.8702,
  -51.9061,
  -51.9441,
  -51.9838,
  -52.0246,
  -52.0665,
  -52.1084,
  -52.1521,
  -52.1964,
  -52.2408,
  -52.2851,
  -52.3291,
  -52.3721,
  -52.4138,
  -52.4544,
  -52.4945,
  -52.5351,
  -52.5772,
  -52.6212,
  -52.667,
  -52.7141,
  -52.7617,
  -52.8087,
  -52.8543,
  -52.8975,
  -52.9369,
  -52.9742,
  -53.0083,
  -53.0397,
  -53.0693,
  -53.0976,
  -53.1255,
  -53.154,
  -53.1835,
  -53.2148,
  -53.2483,
  -53.2839,
  -53.3212,
  -53.3597,
  -53.3988,
  -53.4383,
  -53.4781,
  -53.5183,
  -53.5588,
  -53.5998,
  -53.6411,
  -53.6826,
  -53.7237,
  -53.7653,
  -53.8066,
  -53.8471,
  -53.8864,
  -53.9244,
  -53.9611,
  -53.9965,
  -54.0312,
  -54.0658,
  -54.101,
  -54.1373,
  -54.175,
  -54.2138,
  -54.2534,
  -54.2939,
  -54.3348,
  -54.376,
  -54.4175,
  -54.4592,
  -54.5008,
  -54.5423,
  -54.5836,
  -54.6233,
  -54.6636,
  -54.7035,
  -54.743,
  -54.7817,
  -54.8196,
  -54.8563,
  -54.891,
  -54.9233,
  -54.9531,
  -54.9807,
  -55.0062,
  -55.0303,
  -55.053,
  -55.0749,
  -55.0963,
  -55.1174,
  -55.1381,
  -55.1584,
  -55.1779,
  -55.1965,
  -55.2143,
  -55.2309,
  -55.2463,
  -55.2608,
  -55.274,
  -55.2879,
  -55.3013,
  -55.314,
  -55.3251,
  -55.3338,
  -55.339,
  -55.3403,
  -55.3374,
  -55.3308,
  -55.3215,
  -55.3104,
  -55.2984,
  -55.286,
  -55.2733,
  -55.2604,
  -55.2469,
  -55.2322,
  -55.2158,
  -55.1972,
  -55.1766,
  -55.1538,
  -55.1292,
  -55.103,
  -55.0747,
  -55.0444,
  -55.0123,
  -54.9783,
  -54.9426,
  -54.9044,
  -54.8662,
  -54.8273,
  -54.7874,
  -54.7468,
  -54.705,
  -54.6619,
  -54.6174,
  -54.5714,
  -54.5236,
  -54.4739,
  -54.4225,
  -54.3695,
  -54.3156,
  -54.2606,
  -54.2051,
  -54.1496,
  -54.0947,
  -54.041,
  -53.9886,
  -53.938,
  -53.8892,
  -53.842,
  -53.7959,
  -53.7503,
  -53.7046,
  -53.6582,
  -53.6115,
  -53.5638,
  -53.515,
  -53.4647,
  -53.4132,
  -53.3607,
  -53.3075,
  -53.253,
  -53.1997,
  -53.1468,
  -53.0947,
  -53.0426,
  -52.9904,
  -52.9381,
  -52.8853,
  -52.8321,
  -52.7786,
  -52.7248,
  -52.6713,
  -52.6185,
  -52.5666,
  -52.5162,
  -52.4674,
  -52.4194,
  -52.3727,
  -52.3268,
  -52.2813,
  -52.2359,
  -52.1901,
  -52.1435,
  -52.0961,
  -52.0479,
  -51.9996,
  -51.9517,
  -51.9049,
  -51.86,
  -51.8174,
  -51.7775,
  -51.741,
  -51.7077,
  -51.6777,
  -51.6507,
  -51.6264,
  -51.6041,
  -51.5833,
  -51.5633,
  -51.5437,
  -51.5243,
  -51.5055,
  -51.4879,
  -51.4725,
  -51.4602,
  -51.4507,
  -51.4464,
  -51.4459,
  -51.4486,
  -48.0991,
  -48.252,
  -48.3902,
  -48.5118,
  -48.6159,
  -48.7015,
  -48.7686,
  -48.8172,
  -48.8483,
  -48.864,
  -48.8669,
  -48.8639,
  -48.8603,
  -48.8632,
  -48.8792,
  -48.9141,
  -48.9711,
  -49.0507,
  -49.1503,
  -49.2649,
  -49.3876,
  -49.5116,
  -49.6307,
  -49.7405,
  -49.8387,
  -49.9238,
  -49.9986,
  -50.0643,
  -50.123,
  -50.1773,
  -50.2295,
  -50.2808,
  -50.3319,
  -50.3825,
  -50.4318,
  -50.479,
  -50.5234,
  -50.5648,
  -50.6031,
  -50.6389,
  -50.6726,
  -50.7042,
  -50.7361,
  -50.7676,
  -50.7987,
  -50.829,
  -50.8583,
  -50.8863,
  -50.9131,
  -50.9389,
  -50.9642,
  -50.9893,
  -51.0142,
  -51.0394,
  -51.0645,
  -51.0898,
  -51.1152,
  -51.1396,
  -51.165,
  -51.1904,
  -51.216,
  -51.2416,
  -51.2672,
  -51.2932,
  -51.3196,
  -51.3466,
  -51.374,
  -51.4021,
  -51.4307,
  -51.4594,
  -51.4882,
  -51.5168,
  -51.5447,
  -51.5715,
  -51.5968,
  -51.6192,
  -51.6408,
  -51.6607,
  -51.6793,
  -51.6973,
  -51.7149,
  -51.7327,
  -51.7507,
  -51.7685,
  -51.7863,
  -51.8039,
  -51.8216,
  -51.8397,
  -51.8586,
  -51.8791,
  -51.9016,
  -51.9265,
  -51.9541,
  -51.9835,
  -52.0166,
  -52.0525,
  -52.0908,
  -52.1312,
  -52.1731,
  -52.2162,
  -52.261,
  -52.3068,
  -52.3536,
  -52.4008,
  -52.4482,
  -52.4953,
  -52.5415,
  -52.5866,
  -52.6304,
  -52.6735,
  -52.717,
  -52.7618,
  -52.8074,
  -52.8556,
  -52.9049,
  -52.9544,
  -53.0032,
  -53.0505,
  -53.0951,
  -53.1367,
  -53.1749,
  -53.2099,
  -53.2424,
  -53.2728,
  -53.3022,
  -53.3315,
  -53.3612,
  -53.3921,
  -53.4246,
  -53.4589,
  -53.4951,
  -53.5328,
  -53.5714,
  -53.6095,
  -53.6488,
  -53.6882,
  -53.7278,
  -53.7679,
  -53.8085,
  -53.8498,
  -53.8916,
  -53.9337,
  -53.9762,
  -54.0184,
  -54.0599,
  -54.1005,
  -54.1398,
  -54.1777,
  -54.2144,
  -54.2505,
  -54.2869,
  -54.324,
  -54.362,
  -54.4014,
  -54.4418,
  -54.482,
  -54.5234,
  -54.5653,
  -54.6071,
  -54.6493,
  -54.6916,
  -54.7341,
  -54.7762,
  -54.818,
  -54.8593,
  -54.9,
  -54.9401,
  -54.9797,
  -55.0186,
  -55.0567,
  -55.0936,
  -55.1288,
  -55.1622,
  -55.1935,
  -55.223,
  -55.251,
  -55.2777,
  -55.3032,
  -55.3278,
  -55.3517,
  -55.374,
  -55.3966,
  -55.4189,
  -55.4404,
  -55.461,
  -55.4808,
  -55.4991,
  -55.516,
  -55.5316,
  -55.5462,
  -55.5602,
  -55.5738,
  -55.5863,
  -55.5968,
  -55.6046,
  -55.6087,
  -55.6088,
  -55.6048,
  -55.5972,
  -55.5869,
  -55.575,
  -55.5626,
  -55.5499,
  -55.5373,
  -55.5246,
  -55.5115,
  -55.4974,
  -55.4805,
  -55.4621,
  -55.4412,
  -55.418,
  -55.3928,
  -55.3659,
  -55.3368,
  -55.306,
  -55.2734,
  -55.2388,
  -55.2023,
  -55.164,
  -55.1242,
  -55.0838,
  -55.0428,
  -55.0013,
  -54.9588,
  -54.9151,
  -54.8696,
  -54.8225,
  -54.7732,
  -54.7219,
  -54.669,
  -54.6149,
  -54.5599,
  -54.5042,
  -54.4477,
  -54.3912,
  -54.335,
  -54.28,
  -54.2262,
  -54.1742,
  -54.1229,
  -54.074,
  -54.026,
  -53.9785,
  -53.9309,
  -53.8827,
  -53.8335,
  -53.7834,
  -53.732,
  -53.6794,
  -53.6256,
  -53.5712,
  -53.5165,
  -53.4618,
  -53.4073,
  -53.3534,
  -53.2999,
  -53.2468,
  -53.1936,
  -53.14,
  -53.086,
  -53.0315,
  -52.9767,
  -52.9219,
  -52.8672,
  -52.8132,
  -52.7606,
  -52.7097,
  -52.6605,
  -52.6122,
  -52.5647,
  -52.518,
  -52.4715,
  -52.4247,
  -52.3773,
  -52.3291,
  -52.2797,
  -52.23,
  -52.1804,
  -52.1314,
  -52.0825,
  -52.0365,
  -51.9926,
  -51.9518,
  -51.914,
  -51.8797,
  -51.8487,
  -51.8206,
  -51.7954,
  -51.772,
  -51.7498,
  -51.7282,
  -51.7068,
  -51.6856,
  -51.6651,
  -51.646,
  -51.6293,
  -51.6158,
  -51.6062,
  -51.6007,
  -51.5989,
  -51.6001,
  -48.1213,
  -48.2631,
  -48.3898,
  -48.5002,
  -48.5933,
  -48.667,
  -48.723,
  -48.7599,
  -48.7796,
  -48.7838,
  -48.7774,
  -48.7659,
  -48.7563,
  -48.7566,
  -48.7743,
  -48.8151,
  -48.8823,
  -48.9758,
  -49.0922,
  -49.2248,
  -49.3648,
  -49.5056,
  -49.6399,
  -49.7626,
  -49.8711,
  -49.9653,
  -50.0463,
  -50.1167,
  -50.1794,
  -50.2372,
  -50.2928,
  -50.3477,
  -50.4027,
  -50.4574,
  -50.5109,
  -50.5612,
  -50.6094,
  -50.6539,
  -50.695,
  -50.733,
  -50.7687,
  -50.8027,
  -50.8361,
  -50.8693,
  -50.9023,
  -50.9349,
  -50.9665,
  -50.9969,
  -51.0261,
  -51.054,
  -51.0811,
  -51.1064,
  -51.1327,
  -51.1586,
  -51.1843,
  -51.2099,
  -51.2353,
  -51.2608,
  -51.2863,
  -51.3119,
  -51.3378,
  -51.3638,
  -51.3899,
  -51.4163,
  -51.4429,
  -51.47,
  -51.4976,
  -51.5257,
  -51.5532,
  -51.582,
  -51.6109,
  -51.6399,
  -51.6686,
  -51.6966,
  -51.7235,
  -51.7489,
  -51.7732,
  -51.7963,
  -51.8186,
  -51.8403,
  -51.8617,
  -51.8831,
  -51.904,
  -51.9243,
  -51.9436,
  -51.9621,
  -51.9792,
  -51.9974,
  -52.0163,
  -52.0367,
  -52.0588,
  -52.0834,
  -52.1105,
  -52.1404,
  -52.1731,
  -52.2083,
  -52.2462,
  -52.2863,
  -52.3283,
  -52.3722,
  -52.4181,
  -52.466,
  -52.5154,
  -52.5658,
  -52.6164,
  -52.6658,
  -52.7155,
  -52.7641,
  -52.8114,
  -52.858,
  -52.9045,
  -52.9522,
  -53.0013,
  -53.0517,
  -53.1028,
  -53.1538,
  -53.204,
  -53.2526,
  -53.2984,
  -53.3411,
  -53.3804,
  -53.4166,
  -53.4504,
  -53.4823,
  -53.5132,
  -53.5428,
  -53.5741,
  -53.6065,
  -53.6402,
  -53.6755,
  -53.7121,
  -53.7504,
  -53.7893,
  -53.8286,
  -53.8678,
  -53.9069,
  -53.9462,
  -53.986,
  -54.0264,
  -54.0676,
  -54.1094,
  -54.1518,
  -54.1946,
  -54.2373,
  -54.2795,
  -54.3207,
  -54.3606,
  -54.3982,
  -54.4361,
  -54.4737,
  -54.5116,
  -54.5504,
  -54.5902,
  -54.6311,
  -54.6731,
  -54.7159,
  -54.7589,
  -54.8018,
  -54.8447,
  -54.8878,
  -54.9311,
  -54.9744,
  -55.0177,
  -55.06,
  -55.1017,
  -55.1427,
  -55.1828,
  -55.2225,
  -55.2614,
  -55.2996,
  -55.3357,
  -55.3715,
  -55.4059,
  -55.4388,
  -55.4703,
  -55.5006,
  -55.5299,
  -55.5582,
  -55.5857,
  -55.6121,
  -55.6376,
  -55.6624,
  -55.6865,
  -55.7099,
  -55.7323,
  -55.7539,
  -55.7739,
  -55.7923,
  -55.8089,
  -55.8243,
  -55.8385,
  -55.852,
  -55.864,
  -55.874,
  -55.8811,
  -55.8844,
  -55.8836,
  -55.8778,
  -55.8695,
  -55.8588,
  -55.8467,
  -55.834,
  -55.8215,
  -55.8093,
  -55.7971,
  -55.7844,
  -55.7707,
  -55.755,
  -55.7367,
  -55.7154,
  -55.6914,
  -55.6655,
  -55.6379,
  -55.6085,
  -55.5773,
  -55.5442,
  -55.5094,
  -55.4725,
  -55.4335,
  -55.3928,
  -55.3512,
  -55.3091,
  -55.2669,
  -55.2239,
  -55.1795,
  -55.1332,
  -55.0851,
  -55.0333,
  -54.9807,
  -54.9267,
  -54.8713,
  -54.8152,
  -54.7582,
  -54.7006,
  -54.6427,
  -54.5851,
  -54.5286,
  -54.4732,
  -54.4195,
  -54.3669,
  -54.3156,
  -54.2654,
  -54.2154,
  -54.1653,
  -54.1146,
  -54.0629,
  -54.0103,
  -53.9564,
  -53.9014,
  -53.8456,
  -53.7894,
  -53.7333,
  -53.6773,
  -53.6218,
  -53.5669,
  -53.5123,
  -53.458,
  -53.4037,
  -53.3491,
  -53.294,
  -53.2383,
  -53.1823,
  -53.1263,
  -53.0695,
  -53.0146,
  -52.9613,
  -52.9099,
  -52.8601,
  -52.8115,
  -52.7634,
  -52.7156,
  -52.6678,
  -52.6195,
  -52.5705,
  -52.5206,
  -52.4697,
  -52.4184,
  -52.3678,
  -52.318,
  -52.2695,
  -52.2226,
  -52.1778,
  -52.1357,
  -52.0968,
  -52.0612,
  -52.0289,
  -51.9996,
  -51.973,
  -51.9482,
  -51.9244,
  -51.9011,
  -51.878,
  -51.8553,
  -51.8335,
  -51.8133,
  -51.7956,
  -51.7811,
  -51.7703,
  -51.7635,
  -51.7604,
  -51.7599,
  -48.152,
  -48.2778,
  -48.3888,
  -48.4837,
  -48.5622,
  -48.623,
  -48.6654,
  -48.6896,
  -48.6971,
  -48.6903,
  -48.6752,
  -48.6578,
  -48.6455,
  -48.6469,
  -48.6689,
  -48.7192,
  -48.7993,
  -48.9085,
  -49.0422,
  -49.1925,
  -49.3503,
  -49.5068,
  -49.6545,
  -49.7886,
  -49.9065,
  -50.0083,
  -50.0952,
  -50.1704,
  -50.2373,
  -50.299,
  -50.3574,
  -50.4163,
  -50.4754,
  -50.5342,
  -50.5918,
  -50.647,
  -50.6989,
  -50.7469,
  -50.7911,
  -50.8319,
  -50.8698,
  -50.9058,
  -50.9409,
  -50.976,
  -51.0109,
  -51.0445,
  -51.0783,
  -51.1111,
  -51.1425,
  -51.1726,
  -51.2015,
  -51.2295,
  -51.257,
  -51.2838,
  -51.3104,
  -51.3365,
  -51.3623,
  -51.388,
  -51.4138,
  -51.4398,
  -51.4661,
  -51.4927,
  -51.5184,
  -51.5452,
  -51.5721,
  -51.5993,
  -51.6268,
  -51.6547,
  -51.6829,
  -51.7115,
  -51.7403,
  -51.7693,
  -51.7982,
  -51.8269,
  -51.8548,
  -51.8821,
  -51.9086,
  -51.9347,
  -51.9605,
  -51.9861,
  -52.0107,
  -52.036,
  -52.0605,
  -52.0837,
  -52.1055,
  -52.1259,
  -52.1455,
  -52.1648,
  -52.1844,
  -52.2052,
  -52.2276,
  -52.2518,
  -52.2784,
  -52.3074,
  -52.3391,
  -52.3733,
  -52.4099,
  -52.4487,
  -52.4889,
  -52.5329,
  -52.5796,
  -52.6294,
  -52.6814,
  -52.7348,
  -52.7888,
  -52.8428,
  -52.8958,
  -52.9482,
  -52.9992,
  -53.0493,
  -53.0994,
  -53.1503,
  -53.2019,
  -53.2541,
  -53.3065,
  -53.3589,
  -53.4101,
  -53.4597,
  -53.5053,
  -53.549,
  -53.5897,
  -53.6275,
  -53.6629,
  -53.6964,
  -53.7289,
  -53.7613,
  -53.7941,
  -53.8279,
  -53.8629,
  -53.899,
  -53.9367,
  -53.9756,
  -54.0149,
  -54.0544,
  -54.0937,
  -54.133,
  -54.1723,
  -54.212,
  -54.2525,
  -54.2928,
  -54.3348,
  -54.3773,
  -54.4202,
  -54.463,
  -54.5052,
  -54.5464,
  -54.5864,
  -54.6253,
  -54.6638,
  -54.7025,
  -54.7419,
  -54.7823,
  -54.8238,
  -54.8666,
  -54.9104,
  -54.9546,
  -54.9991,
  -55.0434,
  -55.0877,
  -55.1321,
  -55.1766,
  -55.2202,
  -55.2643,
  -55.3075,
  -55.3496,
  -55.3907,
  -55.4309,
  -55.4706,
  -55.5095,
  -55.5479,
  -55.5853,
  -55.6217,
  -55.6571,
  -55.6914,
  -55.7248,
  -55.7575,
  -55.7893,
  -55.8205,
  -55.8506,
  -55.8797,
  -55.9076,
  -55.9342,
  -55.9599,
  -55.9848,
  -56.009,
  -56.0325,
  -56.0541,
  -56.0725,
  -56.0902,
  -56.1062,
  -56.1211,
  -56.1344,
  -56.1464,
  -56.156,
  -56.1626,
  -56.1653,
  -56.1638,
  -56.1585,
  -56.1501,
  -56.1395,
  -56.1276,
  -56.1154,
  -56.1032,
  -56.0916,
  -56.0799,
  -56.0677,
  -56.0542,
  -56.0383,
  -56.0194,
  -55.9975,
  -55.9729,
  -55.9463,
  -55.9179,
  -55.8881,
  -55.8568,
  -55.8229,
  -55.7879,
  -55.7509,
  -55.7116,
  -55.6706,
  -55.6285,
  -55.5858,
  -55.5428,
  -55.4989,
  -55.4538,
  -55.4069,
  -55.3575,
  -55.3058,
  -55.2519,
  -55.1967,
  -55.1404,
  -55.0828,
  -55.0243,
  -54.9652,
  -54.9057,
  -54.8466,
  -54.7882,
  -54.7309,
  -54.6749,
  -54.62,
  -54.5661,
  -54.5128,
  -54.4599,
  -54.4069,
  -54.3535,
  -54.2993,
  -54.244,
  -54.1876,
  -54.1303,
  -54.0715,
  -54.0136,
  -53.9559,
  -53.8987,
  -53.842,
  -53.786,
  -53.7305,
  -53.6752,
  -53.6199,
  -53.5642,
  -53.5081,
  -53.4515,
  -53.3944,
  -53.3371,
  -53.2802,
  -53.2245,
  -53.1706,
  -53.1186,
  -53.0683,
  -53.019,
  -52.9701,
  -52.9212,
  -52.8717,
  -52.8217,
  -52.7708,
  -52.7191,
  -52.6668,
  -52.6146,
  -52.5631,
  -52.5128,
  -52.4637,
  -52.4163,
  -52.3707,
  -52.3276,
  -52.2874,
  -52.2505,
  -52.2168,
  -52.1861,
  -52.1579,
  -52.1313,
  -52.1057,
  -52.0806,
  -52.0559,
  -52.031,
  -52.0082,
  -51.9873,
  -51.9689,
  -51.9535,
  -51.9416,
  -51.9334,
  -51.9288,
  -51.9266,
  -48.186,
  -48.2927,
  -48.3845,
  -48.4606,
  -48.5209,
  -48.5649,
  -48.5919,
  -48.6026,
  -48.5979,
  -48.5812,
  -48.56,
  -48.5403,
  -48.5303,
  -48.5378,
  -48.571,
  -48.6345,
  -48.7302,
  -48.8561,
  -49.0064,
  -49.1726,
  -49.3452,
  -49.5147,
  -49.674,
  -49.8178,
  -49.943,
  -50.0515,
  -50.1443,
  -50.2244,
  -50.2959,
  -50.3622,
  -50.426,
  -50.4892,
  -50.5524,
  -50.6151,
  -50.6768,
  -50.7359,
  -50.7915,
  -50.843,
  -50.8904,
  -50.9342,
  -50.9738,
  -51.0124,
  -51.0501,
  -51.0871,
  -51.124,
  -51.1608,
  -51.1967,
  -51.2315,
  -51.2649,
  -51.2969,
  -51.3274,
  -51.357,
  -51.3856,
  -51.4138,
  -51.4413,
  -51.4684,
  -51.4941,
  -51.5207,
  -51.5471,
  -51.5739,
  -51.601,
  -51.6282,
  -51.6555,
  -51.6826,
  -51.7097,
  -51.7369,
  -51.7644,
  -51.7921,
  -51.82,
  -51.8481,
  -51.8765,
  -51.9051,
  -51.9338,
  -51.9614,
  -51.99,
  -52.0185,
  -52.047,
  -52.0758,
  -52.1051,
  -52.1349,
  -52.1647,
  -52.1941,
  -52.2225,
  -52.2494,
  -52.2744,
  -52.2977,
  -52.3195,
  -52.3407,
  -52.3618,
  -52.3836,
  -52.4064,
  -52.4296,
  -52.4556,
  -52.4837,
  -52.5141,
  -52.5467,
  -52.5815,
  -52.6185,
  -52.6584,
  -52.7018,
  -52.7489,
  -52.7996,
  -52.8534,
  -52.9093,
  -52.9665,
  -53.024,
  -53.0806,
  -53.1366,
  -53.1914,
  -53.2456,
  -53.2987,
  -53.3526,
  -53.4068,
  -53.4611,
  -53.5153,
  -53.5689,
  -53.6211,
  -53.6713,
  -53.7191,
  -53.7639,
  -53.8056,
  -53.8448,
  -53.8817,
  -53.9169,
  -53.9513,
  -53.9855,
  -54.0202,
  -54.0556,
  -54.092,
  -54.1295,
  -54.1681,
  -54.2064,
  -54.246,
  -54.2857,
  -54.3253,
  -54.3647,
  -54.4042,
  -54.4445,
  -54.4851,
  -54.5266,
  -54.569,
  -54.6116,
  -54.6542,
  -54.697,
  -54.7391,
  -54.7798,
  -54.8196,
  -54.8585,
  -54.8977,
  -54.937,
  -54.9776,
  -55.0193,
  -55.0625,
  -55.1059,
  -55.1513,
  -55.1973,
  -55.2435,
  -55.2896,
  -55.3355,
  -55.3813,
  -55.427,
  -55.4726,
  -55.5174,
  -55.5612,
  -55.6037,
  -55.645,
  -55.6854,
  -55.7253,
  -55.7646,
  -55.8033,
  -55.8413,
  -55.8784,
  -55.9148,
  -55.9506,
  -55.9859,
  -56.0207,
  -56.055,
  -56.0877,
  -56.1207,
  -56.1523,
  -56.1825,
  -56.211,
  -56.2385,
  -56.2649,
  -56.2907,
  -56.3154,
  -56.3384,
  -56.3591,
  -56.3782,
  -56.3952,
  -56.4104,
  -56.4241,
  -56.436,
  -56.4452,
  -56.4513,
  -56.4535,
  -56.4516,
  -56.4462,
  -56.438,
  -56.4279,
  -56.4168,
  -56.4054,
  -56.3941,
  -56.3831,
  -56.371,
  -56.359,
  -56.3451,
  -56.3287,
  -56.3092,
  -56.2866,
  -56.2612,
  -56.2338,
  -56.2048,
  -56.1747,
  -56.1434,
  -56.1107,
  -56.076,
  -56.0391,
  -56.0001,
  -55.9591,
  -55.9168,
  -55.8736,
  -55.8296,
  -55.7846,
  -55.7386,
  -55.6906,
  -55.6402,
  -55.5875,
  -55.5327,
  -55.4763,
  -55.4187,
  -55.3598,
  -55.2998,
  -55.239,
  -55.178,
  -55.1171,
  -55.0556,
  -54.9962,
  -54.9376,
  -54.8801,
  -54.8234,
  -54.7672,
  -54.7113,
  -54.6553,
  -54.5991,
  -54.5424,
  -54.4845,
  -54.4257,
  -54.3661,
  -54.3062,
  -54.2465,
  -54.187,
  -54.1283,
  -54.0703,
  -54.0133,
  -53.9569,
  -53.9007,
  -53.8446,
  -53.7881,
  -53.7311,
  -53.6732,
  -53.6147,
  -53.5563,
  -53.4985,
  -53.4419,
  -53.3871,
  -53.3342,
  -53.283,
  -53.2327,
  -53.1826,
  -53.1323,
  -53.0812,
  -53.0294,
  -52.9769,
  -52.9238,
  -52.8694,
  -52.8164,
  -52.7643,
  -52.7134,
  -52.6638,
  -52.6158,
  -52.5695,
  -52.5255,
  -52.4842,
  -52.4461,
  -52.4111,
  -52.3786,
  -52.3484,
  -52.3196,
  -52.2919,
  -52.2649,
  -52.2388,
  -52.2138,
  -52.1904,
  -52.1691,
  -52.1502,
  -52.1343,
  -52.1217,
  -52.1125,
  -52.1064,
  -52.1026,
  -48.2152,
  -48.3004,
  -48.3707,
  -48.4257,
  -48.4649,
  -48.4902,
  -48.5007,
  -48.4971,
  -48.4819,
  -48.4592,
  -48.4354,
  -48.4179,
  -48.4148,
  -48.4341,
  -48.4821,
  -48.5627,
  -48.6768,
  -48.821,
  -48.9863,
  -49.1669,
  -49.3518,
  -49.5317,
  -49.6991,
  -49.8501,
  -49.9827,
  -50.0971,
  -50.1953,
  -50.2807,
  -50.3573,
  -50.4287,
  -50.4976,
  -50.5656,
  -50.6332,
  -50.7004,
  -50.7649,
  -50.8277,
  -50.8867,
  -50.9416,
  -50.9925,
  -51.0396,
  -51.0836,
  -51.1251,
  -51.1654,
  -51.2048,
  -51.244,
  -51.2827,
  -51.3206,
  -51.3571,
  -51.3922,
  -51.426,
  -51.4571,
  -51.4881,
  -51.5183,
  -51.5479,
  -51.5768,
  -51.6052,
  -51.6333,
  -51.661,
  -51.6886,
  -51.7163,
  -51.7443,
  -51.7724,
  -51.8002,
  -51.8278,
  -51.855,
  -51.8824,
  -51.9098,
  -51.9363,
  -51.9638,
  -51.9916,
  -52.0195,
  -52.0475,
  -52.0757,
  -52.1039,
  -52.1326,
  -52.1619,
  -52.1922,
  -52.2235,
  -52.2561,
  -52.2898,
  -52.324,
  -52.3578,
  -52.3905,
  -52.4212,
  -52.4491,
  -52.4758,
  -52.5007,
  -52.5244,
  -52.5475,
  -52.5708,
  -52.5942,
  -52.6185,
  -52.6439,
  -52.6708,
  -52.6997,
  -52.7304,
  -52.7632,
  -52.7982,
  -52.8363,
  -52.8785,
  -52.9253,
  -52.9766,
  -53.0316,
  -53.0883,
  -53.148,
  -53.2085,
  -53.2688,
  -53.3283,
  -53.3871,
  -53.4454,
  -53.5033,
  -53.5609,
  -53.618,
  -53.6745,
  -53.7306,
  -53.7856,
  -53.839,
  -53.8903,
  -53.9389,
  -53.9847,
  -54.0277,
  -54.0683,
  -54.1068,
  -54.1427,
  -54.179,
  -54.2151,
  -54.2518,
  -54.289,
  -54.3269,
  -54.3657,
  -54.405,
  -54.4448,
  -54.4847,
  -54.5244,
  -54.5641,
  -54.6038,
  -54.6439,
  -54.6846,
  -54.726,
  -54.7679,
  -54.8104,
  -54.8533,
  -54.8959,
  -54.9381,
  -54.9796,
  -55.0191,
  -55.0586,
  -55.0976,
  -55.1369,
  -55.1772,
  -55.2182,
  -55.261,
  -55.3054,
  -55.3514,
  -55.3984,
  -55.4461,
  -55.494,
  -55.542,
  -55.5897,
  -55.6372,
  -55.6843,
  -55.7309,
  -55.7766,
  -55.8209,
  -55.8637,
  -55.9052,
  -55.9459,
  -55.9861,
  -56.0249,
  -56.0641,
  -56.1027,
  -56.1407,
  -56.1782,
  -56.2154,
  -56.2524,
  -56.2892,
  -56.3258,
  -56.3621,
  -56.3976,
  -56.4317,
  -56.4641,
  -56.4946,
  -56.5235,
  -56.5511,
  -56.578,
  -56.6039,
  -56.6281,
  -56.6504,
  -56.6706,
  -56.6888,
  -56.7049,
  -56.7191,
  -56.7311,
  -56.7401,
  -56.745,
  -56.747,
  -56.7453,
  -56.7402,
  -56.7326,
  -56.7235,
  -56.7135,
  -56.7032,
  -56.6931,
  -56.6827,
  -56.672,
  -56.6599,
  -56.6455,
  -56.6283,
  -56.6078,
  -56.5844,
  -56.5583,
  -56.5302,
  -56.5007,
  -56.4701,
  -56.4388,
  -56.4062,
  -56.3719,
  -56.3355,
  -56.2966,
  -56.2559,
  -56.2135,
  -56.1699,
  -56.1251,
  -56.079,
  -56.0306,
  -55.9816,
  -55.93,
  -55.8762,
  -55.8201,
  -55.7625,
  -55.7034,
  -55.6432,
  -55.5818,
  -55.5194,
  -55.4566,
  -55.3938,
  -55.3315,
  -55.2698,
  -55.2087,
  -55.1486,
  -55.0892,
  -55.0303,
  -54.9715,
  -54.9127,
  -54.8538,
  -54.7945,
  -54.7343,
  -54.6732,
  -54.6113,
  -54.5494,
  -54.4876,
  -54.4263,
  -54.3658,
  -54.3061,
  -54.248,
  -54.1908,
  -54.1339,
  -54.077,
  -54.0196,
  -53.9605,
  -53.9014,
  -53.8417,
  -53.7819,
  -53.7228,
  -53.6652,
  -53.6094,
  -53.5555,
  -53.5031,
  -53.4513,
  -53.3996,
  -53.3475,
  -53.2946,
  -53.241,
  -53.1869,
  -53.1326,
  -53.0783,
  -53.0246,
  -52.9719,
  -52.9203,
  -52.8701,
  -52.8215,
  -52.7746,
  -52.7299,
  -52.6879,
  -52.6487,
  -52.6123,
  -52.5783,
  -52.5458,
  -52.5146,
  -52.4847,
  -52.4559,
  -52.4284,
  -52.4025,
  -52.3786,
  -52.3571,
  -52.3381,
  -52.3219,
  -52.3087,
  -52.2985,
  -52.2911,
  -52.2856,
  -48.2329,
  -48.2951,
  -48.3427,
  -48.3758,
  -48.3945,
  -48.3999,
  -48.3934,
  -48.3763,
  -48.3519,
  -48.325,
  -48.3024,
  -48.2918,
  -48.3004,
  -48.3352,
  -48.4029,
  -48.5042,
  -48.6384,
  -48.8007,
  -48.9831,
  -49.1765,
  -49.3711,
  -49.5584,
  -49.7321,
  -49.8882,
  -50.0254,
  -50.1445,
  -50.2478,
  -50.3387,
  -50.4199,
  -50.4968,
  -50.5712,
  -50.6444,
  -50.7169,
  -50.7883,
  -50.8578,
  -50.9242,
  -50.9866,
  -51.0449,
  -51.0993,
  -51.1499,
  -51.1974,
  -51.2424,
  -51.2858,
  -51.328,
  -51.3685,
  -51.4092,
  -51.4489,
  -51.4871,
  -51.5239,
  -51.5592,
  -51.593,
  -51.6255,
  -51.6572,
  -51.6883,
  -51.7188,
  -51.7489,
  -51.7787,
  -51.8081,
  -51.8373,
  -51.8663,
  -51.8954,
  -51.9233,
  -51.952,
  -51.98,
  -52.0078,
  -52.0352,
  -52.0626,
  -52.0902,
  -52.1176,
  -52.1451,
  -52.1725,
  -52.1999,
  -52.2274,
  -52.2551,
  -52.2836,
  -52.3134,
  -52.3449,
  -52.3786,
  -52.4134,
  -52.4509,
  -52.4891,
  -52.5272,
  -52.5642,
  -52.5993,
  -52.6322,
  -52.6627,
  -52.691,
  -52.7179,
  -52.7435,
  -52.7683,
  -52.7927,
  -52.817,
  -52.8418,
  -52.8675,
  -52.8946,
  -52.9233,
  -52.9528,
  -52.9859,
  -53.0224,
  -53.0632,
  -53.1093,
  -53.1601,
  -53.2155,
  -53.2745,
  -53.3361,
  -53.399,
  -53.4622,
  -53.5253,
  -53.5881,
  -53.6505,
  -53.7124,
  -53.7736,
  -53.834,
  -53.8934,
  -53.9517,
  -54.0085,
  -54.0624,
  -54.1151,
  -54.1649,
  -54.2119,
  -54.2562,
  -54.2982,
  -54.3382,
  -54.3768,
  -54.4149,
  -54.4531,
  -54.4918,
  -54.531,
  -54.5707,
  -54.6106,
  -54.6506,
  -54.6906,
  -54.7303,
  -54.7699,
  -54.8096,
  -54.8495,
  -54.8901,
  -54.9304,
  -54.9725,
  -55.0149,
  -55.058,
  -55.1008,
  -55.1435,
  -55.1854,
  -55.2266,
  -55.2666,
  -55.306,
  -55.3451,
  -55.3847,
  -55.425,
  -55.4668,
  -55.5103,
  -55.5556,
  -55.6026,
  -55.651,
  -55.7002,
  -55.7499,
  -55.7996,
  -55.8492,
  -55.8975,
  -55.9462,
  -55.9939,
  -56.0404,
  -56.0852,
  -56.1284,
  -56.1704,
  -56.2116,
  -56.2524,
  -56.2929,
  -56.3328,
  -56.3721,
  -56.4109,
  -56.4495,
  -56.488,
  -56.5265,
  -56.5651,
  -56.6037,
  -56.6423,
  -56.6803,
  -56.7169,
  -56.7513,
  -56.7835,
  -56.814,
  -56.8432,
  -56.8701,
  -56.897,
  -56.9222,
  -56.9457,
  -56.9671,
  -56.9864,
  -57.0035,
  -57.0182,
  -57.0303,
  -57.0395,
  -57.0453,
  -57.0475,
  -57.0463,
  -57.0421,
  -57.0357,
  -57.028,
  -57.0194,
  -57.0103,
  -57.0012,
  -56.9919,
  -56.9815,
  -56.9691,
  -56.9539,
  -56.9358,
  -56.9145,
  -56.8903,
  -56.8634,
  -56.8346,
  -56.8036,
  -56.7727,
  -56.7411,
  -56.7085,
  -56.6742,
  -56.638,
  -56.5995,
  -56.559,
  -56.5167,
  -56.4726,
  -56.4271,
  -56.3796,
  -56.3309,
  -56.2801,
  -56.2271,
  -56.1718,
  -56.1143,
  -56.0552,
  -55.9949,
  -55.9331,
  -55.8703,
  -55.8065,
  -55.7424,
  -55.6777,
  -55.6134,
  -55.5498,
  -55.4867,
  -55.4243,
  -55.3623,
  -55.3007,
  -55.2394,
  -55.1782,
  -55.1169,
  -55.0543,
  -54.9919,
  -54.9287,
  -54.8648,
  -54.8008,
  -54.7368,
  -54.6733,
  -54.6108,
  -54.5496,
  -54.49,
  -54.4315,
  -54.3738,
  -54.3161,
  -54.2577,
  -54.1983,
  -54.1377,
  -54.0764,
  -54.0152,
  -53.9548,
  -53.8961,
  -53.8392,
  -53.7838,
  -53.7297,
  -53.6761,
  -53.6225,
  -53.5683,
  -53.5136,
  -53.4584,
  -53.4028,
  -53.3474,
  -53.2922,
  -53.2376,
  -53.1839,
  -53.1317,
  -53.0806,
  -53.0312,
  -52.9838,
  -52.9386,
  -52.8961,
  -52.8561,
  -52.8184,
  -52.7824,
  -52.747,
  -52.7137,
  -52.6818,
  -52.6513,
  -52.6224,
  -52.5957,
  -52.5713,
  -52.5495,
  -52.5305,
  -52.5141,
  -52.5006,
  -52.4897,
  -52.481,
  -52.4739,
  -48.2372,
  -48.2767,
  -48.3012,
  -48.3114,
  -48.3085,
  -48.294,
  -48.2703,
  -48.2407,
  -48.208,
  -48.1801,
  -48.1629,
  -48.1636,
  -48.1891,
  -48.2456,
  -48.3358,
  -48.46,
  -48.6152,
  -48.7956,
  -48.9929,
  -49.1971,
  -49.3994,
  -49.5923,
  -49.7702,
  -49.929,
  -50.0699,
  -50.1931,
  -50.3012,
  -50.3975,
  -50.4855,
  -50.5684,
  -50.6486,
  -50.7271,
  -50.8043,
  -50.8801,
  -50.9534,
  -51.0236,
  -51.0896,
  -51.1515,
  -51.2086,
  -51.263,
  -51.3141,
  -51.3628,
  -51.4097,
  -51.455,
  -51.4991,
  -51.5419,
  -51.5834,
  -51.6232,
  -51.6615,
  -51.6982,
  -51.7334,
  -51.7676,
  -51.8009,
  -51.8339,
  -51.8655,
  -51.8977,
  -51.9294,
  -51.9606,
  -51.9914,
  -52.022,
  -52.0524,
  -52.0825,
  -52.1121,
  -52.1412,
  -52.1696,
  -52.1977,
  -52.2255,
  -52.2533,
  -52.2808,
  -52.3082,
  -52.3353,
  -52.3611,
  -52.3881,
  -52.4154,
  -52.4437,
  -52.4739,
  -52.5067,
  -52.5425,
  -52.581,
  -52.6217,
  -52.6636,
  -52.7058,
  -52.7469,
  -52.7862,
  -52.8229,
  -52.8573,
  -52.8893,
  -52.9193,
  -52.9476,
  -52.9732,
  -52.9988,
  -53.0235,
  -53.0478,
  -53.0722,
  -53.0974,
  -53.124,
  -53.1525,
  -53.1836,
  -53.2183,
  -53.2575,
  -53.3024,
  -53.3525,
  -53.4076,
  -53.4671,
  -53.5298,
  -53.5948,
  -53.6607,
  -53.7272,
  -53.7925,
  -53.8586,
  -53.9245,
  -53.9897,
  -54.0538,
  -54.1166,
  -54.1775,
  -54.2368,
  -54.2937,
  -54.348,
  -54.3994,
  -54.4476,
  -54.4932,
  -54.5365,
  -54.5782,
  -54.6187,
  -54.6588,
  -54.6992,
  -54.7401,
  -54.7814,
  -54.8226,
  -54.8624,
  -54.9029,
  -54.9427,
  -54.9822,
  -55.0214,
  -55.0609,
  -55.1009,
  -55.1418,
  -55.1836,
  -55.2261,
  -55.2691,
  -55.3123,
  -55.3554,
  -55.398,
  -55.4397,
  -55.4806,
  -55.5205,
  -55.5598,
  -55.5988,
  -55.6382,
  -55.6787,
  -55.7209,
  -55.764,
  -55.8101,
  -55.8584,
  -55.9079,
  -55.9586,
  -56.01,
  -56.0614,
  -56.1129,
  -56.164,
  -56.2143,
  -56.2636,
  -56.3111,
  -56.3569,
  -56.4009,
  -56.4436,
  -56.4854,
  -56.5271,
  -56.5683,
  -56.6089,
  -56.649,
  -56.6887,
  -56.7282,
  -56.7678,
  -56.8076,
  -56.8467,
  -56.8871,
  -56.9278,
  -56.9679,
  -57.0067,
  -57.0432,
  -57.0774,
  -57.1097,
  -57.1402,
  -57.1694,
  -57.1973,
  -57.2235,
  -57.2479,
  -57.2704,
  -57.2904,
  -57.308,
  -57.3231,
  -57.3354,
  -57.3446,
  -57.3506,
  -57.3533,
  -57.3528,
  -57.3498,
  -57.3449,
  -57.3387,
  -57.3317,
  -57.3243,
  -57.3156,
  -57.3071,
  -57.2968,
  -57.2842,
  -57.2685,
  -57.2497,
  -57.2275,
  -57.2024,
  -57.175,
  -57.1459,
  -57.1152,
  -57.0839,
  -57.052,
  -57.0191,
  -56.9848,
  -56.9486,
  -56.9102,
  -56.8695,
  -56.8268,
  -56.782,
  -56.7353,
  -56.6866,
  -56.6358,
  -56.5829,
  -56.5281,
  -56.4712,
  -56.4122,
  -56.3517,
  -56.2899,
  -56.2271,
  -56.1632,
  -56.0972,
  -56.0317,
  -55.9658,
  -55.9004,
  -55.8353,
  -55.7704,
  -55.706,
  -55.6419,
  -55.5781,
  -55.5145,
  -55.451,
  -55.3875,
  -55.3237,
  -55.2593,
  -55.1941,
  -55.1283,
  -55.0622,
  -54.9961,
  -54.9304,
  -54.8659,
  -54.8027,
  -54.7412,
  -54.6813,
  -54.6222,
  -54.5633,
  -54.5035,
  -54.4425,
  -54.3804,
  -54.3175,
  -54.2548,
  -54.193,
  -54.1328,
  -54.0744,
  -54.0173,
  -53.9613,
  -53.9056,
  -53.8497,
  -53.7934,
  -53.7359,
  -53.679,
  -53.622,
  -53.5653,
  -53.5089,
  -53.4533,
  -53.3988,
  -53.3455,
  -53.2936,
  -53.2435,
  -53.1957,
  -53.1501,
  -53.107,
  -53.0661,
  -53.0272,
  -52.9897,
  -52.9535,
  -52.9184,
  -52.8846,
  -52.8526,
  -52.8225,
  -52.7948,
  -52.7699,
  -52.7478,
  -52.7285,
  -52.7119,
  -52.6979,
  -52.6863,
  -52.6766,
  -52.6683,
  -48.2263,
  -48.2435,
  -48.2441,
  -48.2318,
  -48.2072,
  -48.1732,
  -48.133,
  -48.0921,
  -48.0556,
  -48.0296,
  -48.0213,
  -48.0378,
  -48.084,
  -48.1643,
  -48.2799,
  -48.4283,
  -48.6052,
  -48.802,
  -49.0124,
  -49.2259,
  -49.4342,
  -49.6307,
  -49.8111,
  -49.9733,
  -50.1173,
  -50.2446,
  -50.3578,
  -50.4598,
  -50.5541,
  -50.6431,
  -50.729,
  -50.8129,
  -50.894,
  -50.9739,
  -51.0509,
  -51.1244,
  -51.1941,
  -51.2599,
  -51.3218,
  -51.3803,
  -51.4357,
  -51.4883,
  -51.5388,
  -51.5874,
  -51.6343,
  -51.6792,
  -51.7225,
  -51.7639,
  -51.8026,
  -51.8409,
  -51.8778,
  -51.9137,
  -51.9488,
  -51.9836,
  -52.0184,
  -52.0529,
  -52.0869,
  -52.1203,
  -52.153,
  -52.1853,
  -52.2171,
  -52.2486,
  -52.2796,
  -52.31,
  -52.3398,
  -52.3679,
  -52.3967,
  -52.425,
  -52.4529,
  -52.4804,
  -52.5075,
  -52.5342,
  -52.5608,
  -52.588,
  -52.6166,
  -52.6473,
  -52.6813,
  -52.7186,
  -52.7594,
  -52.803,
  -52.8482,
  -52.8938,
  -52.9386,
  -52.9805,
  -53.0211,
  -53.0591,
  -53.0946,
  -53.1277,
  -53.1585,
  -53.1873,
  -53.2142,
  -53.2393,
  -53.2632,
  -53.2866,
  -53.3104,
  -53.3351,
  -53.3618,
  -53.3911,
  -53.4242,
  -53.4621,
  -53.5052,
  -53.5531,
  -53.6073,
  -53.6665,
  -53.7299,
  -53.7962,
  -53.8643,
  -53.9333,
  -54.0028,
  -54.0727,
  -54.1423,
  -54.2115,
  -54.2795,
  -54.3459,
  -54.4104,
  -54.4725,
  -54.5318,
  -54.588,
  -54.641,
  -54.691,
  -54.7381,
  -54.7821,
  -54.8253,
  -54.8677,
  -54.9101,
  -54.9528,
  -54.9959,
  -55.039,
  -55.0816,
  -55.1234,
  -55.164,
  -55.2036,
  -55.2425,
  -55.2814,
  -55.3207,
  -55.3607,
  -55.4016,
  -55.4436,
  -55.4864,
  -55.5298,
  -55.5733,
  -55.6165,
  -55.659,
  -55.6997,
  -55.7404,
  -55.7802,
  -55.8194,
  -55.8584,
  -55.8978,
  -55.9384,
  -55.9808,
  -56.0254,
  -56.0723,
  -56.1213,
  -56.1719,
  -56.2237,
  -56.2764,
  -56.3295,
  -56.3828,
  -56.4357,
  -56.4878,
  -56.5386,
  -56.5875,
  -56.6344,
  -56.6795,
  -56.7234,
  -56.7655,
  -56.8081,
  -56.8502,
  -56.8918,
  -56.9326,
  -56.9731,
  -57.0135,
  -57.0541,
  -57.095,
  -57.1363,
  -57.1783,
  -57.2206,
  -57.2626,
  -57.3033,
  -57.3419,
  -57.378,
  -57.4119,
  -57.4439,
  -57.4743,
  -57.5031,
  -57.5302,
  -57.5554,
  -57.5784,
  -57.5991,
  -57.6171,
  -57.6324,
  -57.6437,
  -57.6532,
  -57.6598,
  -57.6633,
  -57.6641,
  -57.6624,
  -57.659,
  -57.6544,
  -57.6492,
  -57.6434,
  -57.6368,
  -57.6289,
  -57.619,
  -57.6062,
  -57.5901,
  -57.5706,
  -57.5479,
  -57.5224,
  -57.4946,
  -57.4651,
  -57.4342,
  -57.4026,
  -57.3703,
  -57.3369,
  -57.3022,
  -57.2655,
  -57.2267,
  -57.1855,
  -57.1421,
  -57.0953,
  -57.0471,
  -56.9965,
  -56.9435,
  -56.8884,
  -56.8314,
  -56.7725,
  -56.7119,
  -56.6501,
  -56.5871,
  -56.5231,
  -56.4581,
  -56.3922,
  -56.3258,
  -56.2592,
  -56.1928,
  -56.1266,
  -56.0607,
  -55.995,
  -55.9293,
  -55.8636,
  -55.798,
  -55.7324,
  -55.667,
  -55.6012,
  -55.535,
  -55.468,
  -55.4003,
  -55.3322,
  -55.264,
  -55.1962,
  -55.1292,
  -55.0638,
  -55.0003,
  -54.9384,
  -54.8765,
  -54.8158,
  -54.7543,
  -54.6916,
  -54.6277,
  -54.5632,
  -54.4988,
  -54.4355,
  -54.3738,
  -54.3136,
  -54.2546,
  -54.1962,
  -54.1381,
  -54.0801,
  -54.0218,
  -53.9633,
  -53.9047,
  -53.8462,
  -53.7881,
  -53.7305,
  -53.6738,
  -53.6182,
  -53.5639,
  -53.5112,
  -53.4605,
  -53.4122,
  -53.3662,
  -53.3226,
  -53.281,
  -53.2408,
  -53.2018,
  -53.1639,
  -53.1271,
  -53.0918,
  -53.0584,
  -53.0273,
  -52.9987,
  -52.973,
  -52.9503,
  -52.9305,
  -52.9135,
  -52.899,
  -52.8868,
  -52.8763,
  -52.867,
  -48.1999,
  -48.196,
  -48.1758,
  -48.1416,
  -48.0961,
  -48.0433,
  -47.9882,
  -47.9373,
  -47.8975,
  -47.8761,
  -47.8796,
  -47.9144,
  -47.9835,
  -48.0902,
  -48.2321,
  -48.4054,
  -48.6031,
  -48.8175,
  -49.0394,
  -49.2606,
  -49.4735,
  -49.6727,
  -49.855,
  -50.0193,
  -50.1661,
  -50.2975,
  -50.416,
  -50.5234,
  -50.6243,
  -50.7199,
  -50.8117,
  -50.9007,
  -50.9873,
  -51.0712,
  -51.1519,
  -51.2292,
  -51.3025,
  -51.3718,
  -51.4377,
  -51.5005,
  -51.5602,
  -51.617,
  -51.6714,
  -51.7225,
  -51.7723,
  -51.8195,
  -51.8645,
  -51.9073,
  -51.9486,
  -51.9886,
  -52.0274,
  -52.0652,
  -52.1024,
  -52.1393,
  -52.1762,
  -52.2131,
  -52.2496,
  -52.2852,
  -52.3201,
  -52.3534,
  -52.387,
  -52.4202,
  -52.453,
  -52.4853,
  -52.517,
  -52.5478,
  -52.578,
  -52.6075,
  -52.6361,
  -52.6642,
  -52.6916,
  -52.7186,
  -52.7456,
  -52.7732,
  -52.8023,
  -52.8339,
  -52.8679,
  -52.9069,
  -52.9496,
  -52.9953,
  -53.0429,
  -53.0912,
  -53.1389,
  -53.185,
  -53.2289,
  -53.2701,
  -53.3087,
  -53.3447,
  -53.3781,
  -53.409,
  -53.4372,
  -53.4631,
  -53.4872,
  -53.5101,
  -53.5328,
  -53.5552,
  -53.5803,
  -53.6084,
  -53.6402,
  -53.6767,
  -53.7182,
  -53.7653,
  -53.8182,
  -53.8766,
  -53.9398,
  -54.0066,
  -54.076,
  -54.1471,
  -54.2193,
  -54.2924,
  -54.3656,
  -54.4386,
  -54.5107,
  -54.581,
  -54.6482,
  -54.7134,
  -54.7754,
  -54.834,
  -54.889,
  -54.9408,
  -54.9895,
  -55.0362,
  -55.0815,
  -55.1261,
  -55.1709,
  -55.2159,
  -55.2611,
  -55.3059,
  -55.3497,
  -55.392,
  -55.4326,
  -55.472,
  -55.5106,
  -55.5491,
  -55.5883,
  -55.6273,
  -55.6683,
  -55.7103,
  -55.7532,
  -55.7967,
  -55.8403,
  -55.8836,
  -55.9261,
  -55.9676,
  -56.0082,
  -56.0479,
  -56.087,
  -56.1259,
  -56.1653,
  -56.206,
  -56.2487,
  -56.2937,
  -56.341,
  -56.3906,
  -56.4419,
  -56.4947,
  -56.5485,
  -56.6019,
  -56.6568,
  -56.7115,
  -56.7654,
  -56.8179,
  -56.8684,
  -56.9167,
  -56.9633,
  -57.0085,
  -57.0531,
  -57.0971,
  -57.1404,
  -57.183,
  -57.2248,
  -57.2662,
  -57.3076,
  -57.3491,
  -57.391,
  -57.4333,
  -57.4764,
  -57.52,
  -57.5634,
  -57.6056,
  -57.6459,
  -57.6838,
  -57.7185,
  -57.752,
  -57.7835,
  -57.8131,
  -57.8409,
  -57.8667,
  -57.8902,
  -57.9113,
  -57.9295,
  -57.9449,
  -57.9574,
  -57.9673,
  -57.9746,
  -57.9791,
  -57.9811,
  -57.9809,
  -57.9791,
  -57.9761,
  -57.9723,
  -57.9678,
  -57.9622,
  -57.9549,
  -57.9452,
  -57.9324,
  -57.9161,
  -57.8963,
  -57.8734,
  -57.8478,
  -57.819,
  -57.7894,
  -57.7586,
  -57.7268,
  -57.694,
  -57.66,
  -57.6244,
  -57.587,
  -57.5474,
  -57.5054,
  -57.4609,
  -57.4137,
  -57.3637,
  -57.3109,
  -57.2555,
  -57.1977,
  -57.1382,
  -57.0773,
  -57.0151,
  -56.952,
  -56.8878,
  -56.8229,
  -56.7571,
  -56.6905,
  -56.6234,
  -56.5561,
  -56.489,
  -56.4224,
  -56.3559,
  -56.2894,
  -56.2225,
  -56.1555,
  -56.0872,
  -56.0199,
  -55.9526,
  -55.8851,
  -55.817,
  -55.7483,
  -55.6789,
  -55.609,
  -55.5387,
  -55.4686,
  -55.3993,
  -55.3314,
  -55.2655,
  -55.2012,
  -55.1381,
  -55.0751,
  -55.0115,
  -54.9468,
  -54.881,
  -54.8147,
  -54.7488,
  -54.684,
  -54.6206,
  -54.5584,
  -54.4972,
  -54.4365,
  -54.3761,
  -54.3157,
  -54.2553,
  -54.1949,
  -54.1346,
  -54.0746,
  -54.015,
  -53.9562,
  -53.8984,
  -53.8418,
  -53.7866,
  -53.7332,
  -53.682,
  -53.6332,
  -53.5868,
  -53.5415,
  -53.4988,
  -53.4572,
  -53.4167,
  -53.377,
  -53.3387,
  -53.302,
  -53.2675,
  -53.2353,
  -53.2059,
  -53.1794,
  -53.1559,
  -53.1354,
  -53.1177,
  -53.1026,
  -53.0898,
  -53.0786,
  -53.0687,
  -48.1626,
  -48.1387,
  -48.0977,
  -48.043,
  -47.9781,
  -47.9082,
  -47.8386,
  -47.7795,
  -47.7381,
  -47.723,
  -47.7402,
  -47.7954,
  -47.8906,
  -48.0245,
  -48.193,
  -48.39,
  -48.6072,
  -48.8366,
  -49.069,
  -49.2965,
  -49.5132,
  -49.7137,
  -49.898,
  -50.0648,
  -50.2152,
  -50.3512,
  -50.4755,
  -50.5905,
  -50.6984,
  -50.8005,
  -50.8983,
  -50.9926,
  -51.0836,
  -51.1716,
  -51.256,
  -51.3368,
  -51.4136,
  -51.4858,
  -51.556,
  -51.6224,
  -51.6864,
  -51.7476,
  -51.8064,
  -51.8619,
  -51.9147,
  -51.9643,
  -52.011,
  -52.0555,
  -52.0984,
  -52.1403,
  -52.1809,
  -52.221,
  -52.2606,
  -52.2987,
  -52.3378,
  -52.3767,
  -52.4156,
  -52.4537,
  -52.4911,
  -52.5276,
  -52.5634,
  -52.5988,
  -52.6339,
  -52.6685,
  -52.7027,
  -52.7359,
  -52.7682,
  -52.7994,
  -52.8294,
  -52.8585,
  -52.8857,
  -52.9135,
  -52.9415,
  -52.9702,
  -53.0005,
  -53.0332,
  -53.0696,
  -53.1099,
  -53.154,
  -53.2012,
  -53.2504,
  -53.3007,
  -53.3504,
  -53.3988,
  -53.4453,
  -53.4891,
  -53.5305,
  -53.5691,
  -53.6039,
  -53.6367,
  -53.6665,
  -53.6936,
  -53.7184,
  -53.7415,
  -53.7639,
  -53.7867,
  -53.8112,
  -53.8385,
  -53.8693,
  -53.9045,
  -53.9444,
  -53.9898,
  -54.041,
  -54.0979,
  -54.16,
  -54.2264,
  -54.2963,
  -54.3678,
  -54.4421,
  -54.5177,
  -54.5942,
  -54.6709,
  -54.7468,
  -54.8209,
  -54.8927,
  -54.9613,
  -55.0263,
  -55.0875,
  -55.1447,
  -55.1983,
  -55.249,
  -55.2978,
  -55.3454,
  -55.3925,
  -55.4398,
  -55.4871,
  -55.5344,
  -55.5797,
  -55.6243,
  -55.667,
  -55.7076,
  -55.7469,
  -55.7853,
  -55.8238,
  -55.8631,
  -55.9032,
  -55.9443,
  -55.9864,
  -56.0292,
  -56.0727,
  -56.1162,
  -56.1593,
  -56.2016,
  -56.2429,
  -56.2832,
  -56.323,
  -56.3618,
  -56.4007,
  -56.4405,
  -56.4798,
  -56.5226,
  -56.5679,
  -56.6156,
  -56.6656,
  -56.7174,
  -56.7708,
  -56.8254,
  -56.881,
  -56.9372,
  -56.9935,
  -57.0492,
  -57.1032,
  -57.1553,
  -57.2052,
  -57.2534,
  -57.3004,
  -57.3466,
  -57.3921,
  -57.4368,
  -57.4806,
  -57.5236,
  -57.5663,
  -57.6088,
  -57.6504,
  -57.6933,
  -57.7367,
  -57.7807,
  -57.825,
  -57.8691,
  -57.9122,
  -57.9538,
  -57.9934,
  -58.0306,
  -58.0655,
  -58.098,
  -58.1283,
  -58.1568,
  -58.1832,
  -58.2071,
  -58.2285,
  -58.2469,
  -58.2625,
  -58.2754,
  -58.2856,
  -58.2936,
  -58.2992,
  -58.3024,
  -58.3036,
  -58.303,
  -58.3003,
  -58.2978,
  -58.2944,
  -58.2895,
  -58.2826,
  -58.273,
  -58.2602,
  -58.2441,
  -58.2245,
  -58.2017,
  -58.1763,
  -58.1487,
  -58.1195,
  -58.089,
  -58.0571,
  -58.0239,
  -57.9891,
  -57.9527,
  -57.9143,
  -57.8736,
  -57.8305,
  -57.7846,
  -57.7358,
  -57.6838,
  -57.6285,
  -57.5704,
  -57.5101,
  -57.4478,
  -57.3847,
  -57.3208,
  -57.2564,
  -57.1902,
  -57.1246,
  -57.0583,
  -56.9911,
  -56.9235,
  -56.8558,
  -56.7884,
  -56.7213,
  -56.6543,
  -56.5872,
  -56.5198,
  -56.4518,
  -56.3833,
  -56.3145,
  -56.2453,
  -56.1761,
  -56.1063,
  -56.0358,
  -55.9647,
  -55.893,
  -55.8208,
  -55.7487,
  -55.6772,
  -55.6069,
  -55.5383,
  -55.4713,
  -55.4054,
  -55.3398,
  -55.2736,
  -55.2067,
  -55.1391,
  -55.0713,
  -55.0037,
  -54.9373,
  -54.8723,
  -54.808,
  -54.7447,
  -54.6806,
  -54.6177,
  -54.5551,
  -54.4926,
  -54.4303,
  -54.3682,
  -54.3066,
  -54.2456,
  -54.1857,
  -54.127,
  -54.0695,
  -54.0136,
  -53.9596,
  -53.908,
  -53.8588,
  -53.8117,
  -53.7662,
  -53.722,
  -53.6789,
  -53.6365,
  -53.5952,
  -53.5553,
  -53.5174,
  -53.4816,
  -53.4486,
  -53.4184,
  -53.3912,
  -53.3669,
  -53.3455,
  -53.327,
  -53.3112,
  -53.2976,
  -53.286,
  -53.2757,
  -48.1146,
  -48.071,
  -48.0112,
  -47.9377,
  -47.8553,
  -47.7706,
  -47.6911,
  -47.6264,
  -47.5859,
  -47.5782,
  -47.6103,
  -47.6855,
  -47.8043,
  -47.9637,
  -48.1571,
  -48.3763,
  -48.611,
  -48.8543,
  -49.0965,
  -49.3306,
  -49.5512,
  -49.7555,
  -49.9422,
  -50.1121,
  -50.2667,
  -50.4081,
  -50.5387,
  -50.6605,
  -50.7753,
  -50.8842,
  -50.9882,
  -51.0869,
  -51.1827,
  -51.2746,
  -51.3625,
  -51.4467,
  -51.5274,
  -51.6046,
  -51.6787,
  -51.7495,
  -51.8176,
  -51.883,
  -51.9455,
  -52.0048,
  -52.0604,
  -52.1126,
  -52.1617,
  -52.207,
  -52.2518,
  -52.2957,
  -52.3387,
  -52.3811,
  -52.4228,
  -52.4641,
  -52.5051,
  -52.5459,
  -52.587,
  -52.6276,
  -52.6674,
  -52.7064,
  -52.7448,
  -52.7829,
  -52.8207,
  -52.8582,
  -52.8942,
  -52.9302,
  -52.9651,
  -52.9985,
  -53.0306,
  -53.0613,
  -53.091,
  -53.1204,
  -53.15,
  -53.1805,
  -53.2124,
  -53.2468,
  -53.2847,
  -53.3263,
  -53.3716,
  -53.4198,
  -53.47,
  -53.5204,
  -53.5717,
  -53.6218,
  -53.6701,
  -53.716,
  -53.7595,
  -53.8003,
  -53.8382,
  -53.873,
  -53.9045,
  -53.9332,
  -53.9592,
  -53.9834,
  -54.0064,
  -54.0294,
  -54.0539,
  -54.081,
  -54.1114,
  -54.1457,
  -54.1832,
  -54.2271,
  -54.2765,
  -54.3316,
  -54.3921,
  -54.4572,
  -54.5265,
  -54.5991,
  -54.6746,
  -54.7522,
  -54.8311,
  -54.9109,
  -54.9901,
  -55.0677,
  -55.1428,
  -55.2145,
  -55.2827,
  -55.3467,
  -55.4065,
  -55.4614,
  -55.5143,
  -55.5655,
  -55.6155,
  -55.6652,
  -55.7148,
  -55.7641,
  -55.813,
  -55.8606,
  -55.9062,
  -55.9494,
  -55.9903,
  -56.0299,
  -56.0687,
  -56.1078,
  -56.1475,
  -56.1881,
  -56.2297,
  -56.2721,
  -56.3151,
  -56.3585,
  -56.4018,
  -56.4437,
  -56.4856,
  -56.5266,
  -56.5667,
  -56.6061,
  -56.6449,
  -56.6837,
  -56.7231,
  -56.7638,
  -56.8066,
  -56.8518,
  -56.8996,
  -56.9496,
  -57.0016,
  -57.0553,
  -57.1103,
  -57.1666,
  -57.2237,
  -57.2811,
  -57.338,
  -57.3934,
  -57.447,
  -57.4985,
  -57.5473,
  -57.5959,
  -57.6437,
  -57.6908,
  -57.7371,
  -57.7824,
  -57.8268,
  -57.871,
  -57.915,
  -57.9591,
  -58.0032,
  -58.0475,
  -58.0922,
  -58.137,
  -58.1816,
  -58.2253,
  -58.2675,
  -58.3079,
  -58.3461,
  -58.3818,
  -58.4152,
  -58.4463,
  -58.4753,
  -58.5022,
  -58.5266,
  -58.5474,
  -58.5662,
  -58.5822,
  -58.5955,
  -58.6064,
  -58.6151,
  -58.6216,
  -58.6261,
  -58.6285,
  -58.6292,
  -58.6286,
  -58.6269,
  -58.6241,
  -58.6196,
  -58.613,
  -58.6036,
  -58.5909,
  -58.575,
  -58.5557,
  -58.5334,
  -58.5084,
  -58.4813,
  -58.4527,
  -58.4226,
  -58.3909,
  -58.3574,
  -58.3219,
  -58.2847,
  -58.2453,
  -58.2026,
  -58.1581,
  -58.1107,
  -58.0602,
  -58.0062,
  -57.9488,
  -57.8882,
  -57.8253,
  -57.7611,
  -57.696,
  -57.6304,
  -57.5644,
  -57.4981,
  -57.4317,
  -57.3648,
  -57.2973,
  -57.2294,
  -57.1612,
  -57.0934,
  -57.0258,
  -56.9583,
  -56.8905,
  -56.8221,
  -56.7531,
  -56.6834,
  -56.6133,
  -56.5427,
  -56.4716,
  -56.4002,
  -56.3281,
  -56.2555,
  -56.1822,
  -56.1083,
  -56.0344,
  -55.9599,
  -55.8873,
  -55.8161,
  -55.7463,
  -55.6775,
  -55.6091,
  -55.5405,
  -55.4713,
  -55.4017,
  -55.3322,
  -55.2632,
  -55.1953,
  -55.1285,
  -55.0625,
  -54.997,
  -54.9318,
  -54.8667,
  -54.8017,
  -54.7368,
  -54.6722,
  -54.6082,
  -54.5448,
  -54.4825,
  -54.4213,
  -54.3617,
  -54.3036,
  -54.2473,
  -54.1929,
  -54.1408,
  -54.0908,
  -54.0426,
  -53.9958,
  -53.95,
  -53.905,
  -53.861,
  -53.8182,
  -53.777,
  -53.7378,
  -53.7011,
  -53.6671,
  -53.6362,
  -53.6083,
  -53.5833,
  -53.5612,
  -53.5418,
  -53.5242,
  -53.51,
  -53.4977,
  -53.4869,
  -48.0584,
  -47.9983,
  -47.9212,
  -47.831,
  -47.7337,
  -47.6368,
  -47.5492,
  -47.4812,
  -47.443,
  -47.4439,
  -47.4895,
  -47.5839,
  -47.7251,
  -47.9075,
  -48.1227,
  -48.3615,
  -48.6132,
  -48.8686,
  -49.12,
  -49.3606,
  -49.5861,
  -49.7943,
  -49.9851,
  -50.1594,
  -50.3196,
  -50.4663,
  -50.6041,
  -50.7332,
  -50.8551,
  -50.9706,
  -51.0805,
  -51.1856,
  -51.2861,
  -51.3822,
  -51.474,
  -51.5619,
  -51.6462,
  -51.7273,
  -51.8052,
  -51.8802,
  -51.9524,
  -52.0206,
  -52.0867,
  -52.1492,
  -52.208,
  -52.263,
  -52.3147,
  -52.3638,
  -52.4111,
  -52.4574,
  -52.5028,
  -52.5474,
  -52.5914,
  -52.6345,
  -52.6771,
  -52.7199,
  -52.7627,
  -52.8056,
  -52.8471,
  -52.8889,
  -52.9302,
  -52.9714,
  -53.0124,
  -53.053,
  -53.0931,
  -53.1322,
  -53.17,
  -53.2063,
  -53.2408,
  -53.2738,
  -53.3057,
  -53.3375,
  -53.3693,
  -53.4019,
  -53.4362,
  -53.4718,
  -53.5114,
  -53.5544,
  -53.6004,
  -53.6493,
  -53.7001,
  -53.7521,
  -53.8041,
  -53.8552,
  -53.9047,
  -53.9521,
  -53.9973,
  -54.0399,
  -54.0796,
  -54.1163,
  -54.15,
  -54.1808,
  -54.2089,
  -54.2338,
  -54.2585,
  -54.2828,
  -54.3084,
  -54.336,
  -54.3664,
  -54.4003,
  -54.438,
  -54.4806,
  -54.528,
  -54.5806,
  -54.6386,
  -54.7014,
  -54.7691,
  -54.8407,
  -54.9161,
  -54.9949,
  -55.0759,
  -55.1582,
  -55.2391,
  -55.3196,
  -55.3978,
  -55.4727,
  -55.5441,
  -55.6109,
  -55.6733,
  -55.7319,
  -55.7874,
  -55.8412,
  -55.8938,
  -55.9457,
  -55.9973,
  -56.0483,
  -56.0987,
  -56.1473,
  -56.1936,
  -56.2375,
  -56.2792,
  -56.3197,
  -56.3594,
  -56.3983,
  -56.439,
  -56.4805,
  -56.523,
  -56.5658,
  -56.6088,
  -56.6521,
  -56.6952,
  -56.7377,
  -56.7792,
  -56.8197,
  -56.8594,
  -56.8985,
  -56.9372,
  -56.9759,
  -57.0153,
  -57.0561,
  -57.0993,
  -57.1441,
  -57.1917,
  -57.2417,
  -57.2939,
  -57.3466,
  -57.4018,
  -57.4582,
  -57.5155,
  -57.5733,
  -57.6308,
  -57.6871,
  -57.7418,
  -57.7947,
  -57.8461,
  -57.8965,
  -57.9461,
  -57.9948,
  -58.0427,
  -58.0897,
  -58.136,
  -58.182,
  -58.2278,
  -58.2734,
  -58.3189,
  -58.3643,
  -58.4097,
  -58.4548,
  -58.4994,
  -58.5431,
  -58.5845,
  -58.6254,
  -58.6641,
  -58.7004,
  -58.7342,
  -58.766,
  -58.7957,
  -58.823,
  -58.8477,
  -58.8699,
  -58.8891,
  -58.9054,
  -58.9192,
  -58.9307,
  -58.9402,
  -58.9476,
  -58.9532,
  -58.957,
  -58.9584,
  -58.9585,
  -58.9574,
  -58.9551,
  -58.9507,
  -58.9441,
  -58.9348,
  -58.9223,
  -58.9068,
  -58.887,
  -58.8651,
  -58.8407,
  -58.8143,
  -58.7865,
  -58.7569,
  -58.7255,
  -58.6919,
  -58.6562,
  -58.6182,
  -58.5778,
  -58.5349,
  -58.4892,
  -58.4403,
  -58.3883,
  -58.3325,
  -58.2731,
  -58.2106,
  -58.1458,
  -58.0798,
  -58.0129,
  -57.9456,
  -57.8784,
  -57.8112,
  -57.744,
  -57.6767,
  -57.609,
  -57.5409,
  -57.4723,
  -57.404,
  -57.3356,
  -57.2671,
  -57.1974,
  -57.128,
  -57.0579,
  -56.9871,
  -56.9155,
  -56.8434,
  -56.7707,
  -56.6976,
  -56.624,
  -56.5498,
  -56.4753,
  -56.4,
  -56.3246,
  -56.2493,
  -56.1746,
  -56.101,
  -56.0284,
  -55.9568,
  -55.8856,
  -55.8144,
  -55.7431,
  -55.6715,
  -55.6004,
  -55.5299,
  -55.4604,
  -55.3918,
  -55.324,
  -55.2567,
  -55.1894,
  -55.122,
  -55.0546,
  -54.9873,
  -54.9205,
  -54.8544,
  -54.7893,
  -54.7255,
  -54.6633,
  -54.6029,
  -54.5443,
  -54.4877,
  -54.432,
  -54.3792,
  -54.3284,
  -54.2788,
  -54.2304,
  -54.1827,
  -54.1359,
  -54.0904,
  -54.0462,
  -54.0038,
  -53.9633,
  -53.9254,
  -53.8905,
  -53.8588,
  -53.8302,
  -53.8047,
  -53.7819,
  -53.7618,
  -53.7444,
  -53.7294,
  -53.7166,
  -53.7052,
  -47.9951,
  -47.9188,
  -47.8265,
  -47.7224,
  -47.6135,
  -47.5069,
  -47.4147,
  -47.3467,
  -47.3131,
  -47.3233,
  -47.3832,
  -47.4944,
  -47.6543,
  -47.8557,
  -48.0893,
  -48.3443,
  -48.6099,
  -48.8767,
  -49.1367,
  -49.3846,
  -49.6151,
  -49.8289,
  -50.0251,
  -50.2056,
  -50.3724,
  -50.5277,
  -50.6731,
  -50.81,
  -50.9393,
  -51.0616,
  -51.1778,
  -51.2881,
  -51.3933,
  -51.4939,
  -51.5899,
  -51.6807,
  -51.7688,
  -51.8535,
  -51.9353,
  -52.0144,
  -52.0904,
  -52.1633,
  -52.2328,
  -52.2985,
  -52.3602,
  -52.4182,
  -52.4729,
  -52.5253,
  -52.5756,
  -52.6249,
  -52.673,
  -52.719,
  -52.7648,
  -52.8097,
  -52.8541,
  -52.8982,
  -52.9427,
  -52.9874,
  -53.0323,
  -53.0772,
  -53.1217,
  -53.1662,
  -53.2104,
  -53.2545,
  -53.2978,
  -53.3402,
  -53.3812,
  -53.4206,
  -53.457,
  -53.493,
  -53.5278,
  -53.5622,
  -53.5969,
  -53.6321,
  -53.669,
  -53.7079,
  -53.7494,
  -53.7937,
  -53.8409,
  -53.8904,
  -53.9417,
  -53.994,
  -54.0463,
  -54.098,
  -54.1484,
  -54.197,
  -54.2425,
  -54.2867,
  -54.3283,
  -54.3671,
  -54.403,
  -54.4362,
  -54.4667,
  -54.4954,
  -54.5225,
  -54.549,
  -54.5763,
  -54.6052,
  -54.6366,
  -54.6707,
  -54.708,
  -54.7492,
  -54.7946,
  -54.8449,
  -54.9,
  -54.9589,
  -55.0238,
  -55.0934,
  -55.1678,
  -55.2467,
  -55.3285,
  -55.4122,
  -55.4962,
  -55.5793,
  -55.6602,
  -55.7381,
  -55.8123,
  -55.8821,
  -55.9475,
  -56.009,
  -56.0672,
  -56.1235,
  -56.1783,
  -56.2324,
  -56.2857,
  -56.3371,
  -56.3885,
  -56.4379,
  -56.4853,
  -56.5302,
  -56.573,
  -56.6145,
  -56.6555,
  -56.6969,
  -56.739,
  -56.7818,
  -56.8251,
  -56.8683,
  -56.9116,
  -56.9549,
  -56.9977,
  -57.0399,
  -57.0812,
  -57.1216,
  -57.1611,
  -57.2002,
  -57.239,
  -57.2771,
  -57.3168,
  -57.3578,
  -57.4006,
  -57.4457,
  -57.4932,
  -57.5428,
  -57.5944,
  -57.6478,
  -57.7028,
  -57.7589,
  -57.8156,
  -57.8729,
  -57.9303,
  -57.9869,
  -58.0422,
  -58.0961,
  -58.1489,
  -58.2009,
  -58.2523,
  -58.3028,
  -58.3526,
  -58.4017,
  -58.4491,
  -58.4971,
  -58.5447,
  -58.592,
  -58.6389,
  -58.6853,
  -58.7312,
  -58.7765,
  -58.8211,
  -58.8646,
  -58.9068,
  -58.9475,
  -58.986,
  -59.0225,
  -59.0566,
  -59.0887,
  -59.1187,
  -59.1463,
  -59.1715,
  -59.1938,
  -59.2133,
  -59.2301,
  -59.2446,
  -59.257,
  -59.2673,
  -59.2762,
  -59.2827,
  -59.2863,
  -59.2886,
  -59.2892,
  -59.2883,
  -59.2856,
  -59.2809,
  -59.274,
  -59.2645,
  -59.2522,
  -59.2368,
  -59.2184,
  -59.1972,
  -59.1736,
  -59.148,
  -59.1209,
  -59.0918,
  -59.0608,
  -59.0273,
  -58.9913,
  -58.9528,
  -58.9116,
  -58.8679,
  -58.821,
  -58.7711,
  -58.718,
  -58.6612,
  -58.6009,
  -58.5374,
  -58.4717,
  -58.4044,
  -58.3352,
  -58.2668,
  -58.1983,
  -58.1301,
  -58.0621,
  -57.9941,
  -57.926,
  -57.8575,
  -57.7887,
  -57.7194,
  -57.6501,
  -57.5805,
  -57.5105,
  -57.4397,
  -57.3682,
  -57.2959,
  -57.223,
  -57.1493,
  -57.075,
  -57.0005,
  -56.9254,
  -56.8502,
  -56.7744,
  -56.698,
  -56.6213,
  -56.5446,
  -56.4682,
  -56.3924,
  -56.3175,
  -56.2434,
  -56.1697,
  -56.0962,
  -56.0227,
  -55.9491,
  -55.876,
  -55.8036,
  -55.7312,
  -55.6608,
  -55.591,
  -55.5218,
  -55.4524,
  -55.3829,
  -55.3132,
  -55.2436,
  -55.1745,
  -55.1064,
  -55.0396,
  -54.9745,
  -54.9112,
  -54.85,
  -54.7908,
  -54.7335,
  -54.6782,
  -54.6247,
  -54.5728,
  -54.5219,
  -54.4717,
  -54.4224,
  -54.3741,
  -54.3272,
  -54.282,
  -54.2384,
  -54.1967,
  -54.1577,
  -54.1217,
  -54.0892,
  -54.0598,
  -54.0335,
  -54.01,
  -53.9892,
  -53.971,
  -53.9553,
  -53.942,
  -53.9299,
  -47.9244,
  -47.8333,
  -47.7274,
  -47.6121,
  -47.4953,
  -47.385,
  -47.292,
  -47.2268,
  -47.1999,
  -47.2197,
  -47.2918,
  -47.4171,
  -47.5919,
  -47.808,
  -48.0544,
  -48.3221,
  -48.5991,
  -48.8756,
  -49.1446,
  -49.4,
  -49.639,
  -49.8601,
  -50.0638,
  -50.2521,
  -50.4271,
  -50.5907,
  -50.7445,
  -50.8894,
  -51.0262,
  -51.1556,
  -51.2771,
  -51.3931,
  -51.5033,
  -51.6086,
  -51.709,
  -51.8052,
  -51.8975,
  -51.9862,
  -52.0719,
  -52.1545,
  -52.2342,
  -52.3106,
  -52.3833,
  -52.452,
  -52.5167,
  -52.5776,
  -52.6347,
  -52.6903,
  -52.7443,
  -52.7968,
  -52.8479,
  -52.8974,
  -52.9453,
  -52.9919,
  -53.0378,
  -53.0831,
  -53.1289,
  -53.1754,
  -53.2226,
  -53.2702,
  -53.3181,
  -53.3662,
  -53.413,
  -53.4604,
  -53.5072,
  -53.5529,
  -53.597,
  -53.6398,
  -53.6807,
  -53.72,
  -53.7582,
  -53.7958,
  -53.8334,
  -53.8716,
  -53.9112,
  -53.9526,
  -53.9962,
  -54.042,
  -54.0903,
  -54.1405,
  -54.1913,
  -54.2438,
  -54.2964,
  -54.3484,
  -54.3993,
  -54.4488,
  -54.4966,
  -54.5422,
  -54.5856,
  -54.6266,
  -54.6651,
  -54.7013,
  -54.735,
  -54.7668,
  -54.797,
  -54.8267,
  -54.8566,
  -54.8875,
  -54.9192,
  -54.9541,
  -54.9916,
  -55.0318,
  -55.0754,
  -55.1231,
  -55.175,
  -55.2316,
  -55.2931,
  -55.3599,
  -55.4323,
  -55.51,
  -55.5919,
  -55.6763,
  -55.7617,
  -55.8467,
  -55.93,
  -56.0106,
  -56.0875,
  -56.16,
  -56.2272,
  -56.2914,
  -56.3525,
  -56.4112,
  -56.4681,
  -56.5239,
  -56.5786,
  -56.6323,
  -56.6846,
  -56.7349,
  -56.783,
  -56.8291,
  -56.8734,
  -56.9164,
  -56.9589,
  -57.0018,
  -57.0455,
  -57.0896,
  -57.1338,
  -57.1776,
  -57.2212,
  -57.2636,
  -57.3066,
  -57.3487,
  -57.3898,
  -57.4299,
  -57.4696,
  -57.5088,
  -57.5482,
  -57.588,
  -57.6285,
  -57.6701,
  -57.7132,
  -57.7582,
  -57.8053,
  -57.8545,
  -57.9057,
  -57.9586,
  -58.0128,
  -58.0681,
  -58.1238,
  -58.1801,
  -58.2365,
  -58.2915,
  -58.3469,
  -58.4014,
  -58.4553,
  -58.5087,
  -58.5618,
  -58.6143,
  -58.6663,
  -58.7175,
  -58.7683,
  -58.8184,
  -58.8679,
  -58.9167,
  -58.9647,
  -59.012,
  -59.0585,
  -59.1039,
  -59.1483,
  -59.1911,
  -59.2326,
  -59.2726,
  -59.3107,
  -59.3468,
  -59.3809,
  -59.413,
  -59.4432,
  -59.4699,
  -59.495,
  -59.5173,
  -59.5369,
  -59.5541,
  -59.5695,
  -59.583,
  -59.5948,
  -59.6045,
  -59.6123,
  -59.6175,
  -59.6204,
  -59.6209,
  -59.6197,
  -59.6163,
  -59.6109,
  -59.6032,
  -59.5933,
  -59.5809,
  -59.5655,
  -59.5474,
  -59.5268,
  -59.504,
  -59.4793,
  -59.4528,
  -59.4242,
  -59.3935,
  -59.3602,
  -59.3235,
  -59.2846,
  -59.2429,
  -59.1983,
  -59.1508,
  -59.1005,
  -59.047,
  -58.9901,
  -58.9298,
  -58.8664,
  -58.8005,
  -58.7329,
  -58.664,
  -58.5947,
  -58.5255,
  -58.4566,
  -58.388,
  -58.3193,
  -58.2507,
  -58.1816,
  -58.1123,
  -58.0421,
  -57.9716,
  -57.9007,
  -57.8291,
  -57.7568,
  -57.6837,
  -57.6096,
  -57.5349,
  -57.4596,
  -57.384,
  -57.308,
  -57.2317,
  -57.1551,
  -57.0774,
  -57.0002,
  -56.9224,
  -56.8445,
  -56.7667,
  -56.6893,
  -56.6126,
  -56.5365,
  -56.4607,
  -56.385,
  -56.3093,
  -56.2338,
  -56.1585,
  -56.0839,
  -56.0103,
  -55.9376,
  -55.8657,
  -55.7944,
  -55.723,
  -55.6517,
  -55.5798,
  -55.5082,
  -55.4372,
  -55.367,
  -55.2986,
  -55.232,
  -55.1677,
  -55.1055,
  -55.0453,
  -54.9873,
  -54.9312,
  -54.8767,
  -54.8235,
  -54.7712,
  -54.7195,
  -54.6686,
  -54.6191,
  -54.5712,
  -54.525,
  -54.4809,
  -54.4386,
  -54.3982,
  -54.3609,
  -54.326,
  -54.2957,
  -54.2688,
  -54.2446,
  -54.2232,
  -54.2041,
  -54.1876,
  -54.1733,
  -54.1608,
  -47.8487,
  -47.7439,
  -47.6266,
  -47.5038,
  -47.382,
  -47.2709,
  -47.1809,
  -47.1221,
  -47.1038,
  -47.1327,
  -47.2154,
  -47.3515,
  -47.5366,
  -47.7632,
  -48.0202,
  -48.2969,
  -48.583,
  -48.8683,
  -49.1458,
  -49.4099,
  -49.6573,
  -49.8874,
  -50.1004,
  -50.298,
  -50.4814,
  -50.6543,
  -50.8169,
  -50.97,
  -51.1146,
  -51.2509,
  -51.3798,
  -51.5018,
  -51.6174,
  -51.7277,
  -51.8332,
  -51.9339,
  -52.0309,
  -52.1241,
  -52.2139,
  -52.3003,
  -52.3824,
  -52.4618,
  -52.5374,
  -52.6092,
  -52.677,
  -52.7412,
  -52.8026,
  -52.8618,
  -52.9194,
  -52.9753,
  -53.0294,
  -53.0816,
  -53.1317,
  -53.1802,
  -53.2275,
  -53.2744,
  -53.3204,
  -53.3684,
  -53.4174,
  -53.4678,
  -53.5191,
  -53.5708,
  -53.6222,
  -53.6732,
  -53.7234,
  -53.7724,
  -53.8201,
  -53.8661,
  -53.9104,
  -53.9535,
  -53.9952,
  -54.0362,
  -54.0771,
  -54.1175,
  -54.1597,
  -54.2036,
  -54.2493,
  -54.2968,
  -54.3463,
  -54.3973,
  -54.4497,
  -54.5027,
  -54.5556,
  -54.6079,
  -54.6593,
  -54.7096,
  -54.7585,
  -54.8057,
  -54.8511,
  -54.8944,
  -54.9358,
  -54.9742,
  -55.0115,
  -55.047,
  -55.081,
  -55.1143,
  -55.1474,
  -55.181,
  -55.2157,
  -55.2517,
  -55.2895,
  -55.3292,
  -55.3714,
  -55.4168,
  -55.4657,
  -55.5188,
  -55.5768,
  -55.6404,
  -55.7102,
  -55.7858,
  -55.8656,
  -55.9498,
  -56.0359,
  -56.1223,
  -56.2076,
  -56.2904,
  -56.3697,
  -56.4447,
  -56.5155,
  -56.5822,
  -56.6456,
  -56.7064,
  -56.7652,
  -56.8226,
  -56.8786,
  -56.9334,
  -56.9866,
  -57.0378,
  -57.0871,
  -57.1343,
  -57.1798,
  -57.2233,
  -57.2673,
  -57.3119,
  -57.357,
  -57.4022,
  -57.4473,
  -57.4916,
  -57.5354,
  -57.5788,
  -57.622,
  -57.6645,
  -57.7054,
  -57.7459,
  -57.786,
  -57.826,
  -57.8666,
  -57.9074,
  -57.9489,
  -57.9916,
  -58.0354,
  -58.0806,
  -58.1274,
  -58.1753,
  -58.226,
  -58.2782,
  -58.3317,
  -58.3856,
  -58.44,
  -58.4948,
  -58.5495,
  -58.6044,
  -58.6592,
  -58.7138,
  -58.7684,
  -58.8231,
  -58.8777,
  -58.9322,
  -58.9863,
  -59.0397,
  -59.0927,
  -59.1449,
  -59.1961,
  -59.2461,
  -59.295,
  -59.343,
  -59.3899,
  -59.4344,
  -59.4782,
  -59.5203,
  -59.5606,
  -59.5994,
  -59.6365,
  -59.6719,
  -59.7055,
  -59.7374,
  -59.7674,
  -59.7949,
  -59.8197,
  -59.8417,
  -59.8614,
  -59.8791,
  -59.8952,
  -59.9099,
  -59.923,
  -59.934,
  -59.9425,
  -59.9483,
  -59.9514,
  -59.9518,
  -59.9496,
  -59.9452,
  -59.9385,
  -59.9299,
  -59.918,
  -59.9048,
  -59.8893,
  -59.8713,
  -59.8513,
  -59.8292,
  -59.8052,
  -59.7792,
  -59.751,
  -59.7204,
  -59.6874,
  -59.6516,
  -59.6129,
  -59.5711,
  -59.5263,
  -59.4787,
  -59.4285,
  -59.3756,
  -59.3196,
  -59.2604,
  -59.198,
  -59.1329,
  -59.0658,
  -58.9969,
  -58.9275,
  -58.8579,
  -58.7887,
  -58.7196,
  -58.6505,
  -58.5813,
  -58.5116,
  -58.4414,
  -58.3696,
  -58.2979,
  -58.2256,
  -58.1524,
  -58.0783,
  -58.0033,
  -57.9274,
  -57.8509,
  -57.7739,
  -57.6967,
  -57.6193,
  -57.5417,
  -57.4643,
  -57.3865,
  -57.3084,
  -57.2299,
  -57.1511,
  -57.0723,
  -56.9938,
  -56.9157,
  -56.838,
  -56.7605,
  -56.6828,
  -56.6051,
  -56.5273,
  -56.4499,
  -56.3727,
  -56.2966,
  -56.2213,
  -56.1471,
  -56.0736,
  -56.0004,
  -55.9271,
  -55.8536,
  -55.7801,
  -55.7072,
  -55.6355,
  -55.5654,
  -55.4973,
  -55.4307,
  -55.3673,
  -55.3061,
  -55.2473,
  -55.19,
  -55.1342,
  -55.0796,
  -55.0257,
  -54.973,
  -54.9211,
  -54.8705,
  -54.8218,
  -54.775,
  -54.7301,
  -54.6866,
  -54.6453,
  -54.6069,
  -54.5719,
  -54.5405,
  -54.5126,
  -54.4877,
  -54.4655,
  -54.4458,
  -54.4286,
  -54.4131,
  -54.3993,
  -47.768,
  -47.6506,
  -47.5242,
  -47.3968,
  -47.2731,
  -47.1649,
  -47.0816,
  -47.0319,
  -47.024,
  -47.0641,
  -47.156,
  -47.2998,
  -47.4914,
  -47.7237,
  -47.9864,
  -48.2691,
  -48.5618,
  -48.8549,
  -49.1409,
  -49.4134,
  -49.6706,
  -49.9109,
  -50.1346,
  -50.3429,
  -50.5376,
  -50.7203,
  -50.8919,
  -51.0535,
  -51.2056,
  -51.3489,
  -51.4843,
  -51.6125,
  -51.7342,
  -51.8501,
  -51.9598,
  -52.0659,
  -52.1677,
  -52.2657,
  -52.36,
  -52.4504,
  -52.5369,
  -52.6193,
  -52.6976,
  -52.7723,
  -52.8433,
  -52.911,
  -52.9762,
  -53.0392,
  -53.1003,
  -53.1598,
  -53.2158,
  -53.2708,
  -53.3233,
  -53.3738,
  -53.4228,
  -53.4712,
  -53.5201,
  -53.5698,
  -53.6208,
  -53.6734,
  -53.7276,
  -53.7828,
  -53.8379,
  -53.8926,
  -53.9461,
  -53.9984,
  -54.0493,
  -54.0977,
  -54.1457,
  -54.1924,
  -54.2377,
  -54.2821,
  -54.3262,
  -54.3707,
  -54.4159,
  -54.4622,
  -54.5099,
  -54.5592,
  -54.6101,
  -54.6621,
  -54.7151,
  -54.7685,
  -54.8219,
  -54.8748,
  -54.927,
  -54.9772,
  -55.0272,
  -55.0762,
  -55.1239,
  -55.1698,
  -55.2141,
  -55.2569,
  -55.298,
  -55.3376,
  -55.3758,
  -55.413,
  -55.4497,
  -55.4863,
  -55.5234,
  -55.5609,
  -55.5993,
  -55.6388,
  -55.6801,
  -55.7228,
  -55.7692,
  -55.8194,
  -55.8742,
  -55.9347,
  -56.0014,
  -56.0742,
  -56.1529,
  -56.2361,
  -56.3222,
  -56.4095,
  -56.496,
  -56.5806,
  -56.6618,
  -56.739,
  -56.812,
  -56.8808,
  -56.9461,
  -57.0087,
  -57.0692,
  -57.1271,
  -57.1845,
  -57.2404,
  -57.2946,
  -57.3469,
  -57.3973,
  -57.4453,
  -57.4918,
  -57.5375,
  -57.5829,
  -57.6288,
  -57.6748,
  -57.721,
  -57.7666,
  -57.8113,
  -57.8554,
  -57.8989,
  -57.9421,
  -57.9847,
  -58.0267,
  -58.068,
  -58.1089,
  -58.1489,
  -58.1907,
  -58.2333,
  -58.2766,
  -58.3209,
  -58.3653,
  -58.411,
  -58.4582,
  -58.5067,
  -58.557,
  -58.6087,
  -58.661,
  -58.7137,
  -58.7665,
  -58.8196,
  -58.8725,
  -58.9258,
  -58.9795,
  -59.0338,
  -59.0886,
  -59.1441,
  -59.1999,
  -59.2559,
  -59.3109,
  -59.3666,
  -59.4215,
  -59.4756,
  -59.5282,
  -59.5792,
  -59.6288,
  -59.6771,
  -59.724,
  -59.7692,
  -59.8123,
  -59.8531,
  -59.892,
  -59.9292,
  -59.965,
  -59.9994,
  -60.0322,
  -60.0635,
  -60.0929,
  -60.1199,
  -60.1442,
  -60.1658,
  -60.1854,
  -60.2035,
  -60.2204,
  -60.2361,
  -60.2492,
  -60.261,
  -60.2702,
  -60.2764,
  -60.2794,
  -60.2792,
  -60.276,
  -60.27,
  -60.2618,
  -60.2517,
  -60.2395,
  -60.2252,
  -60.2088,
  -60.191,
  -60.1713,
  -60.1496,
  -60.1261,
  -60.1004,
  -60.0723,
  -60.0418,
  -60.0088,
  -59.9731,
  -59.9345,
  -59.8929,
  -59.8486,
  -59.8016,
  -59.7523,
  -59.7007,
  -59.6465,
  -59.5893,
  -59.5278,
  -59.4642,
  -59.3982,
  -59.3305,
  -59.2616,
  -59.1923,
  -59.1231,
  -59.0539,
  -58.9845,
  -58.915,
  -58.8449,
  -58.7744,
  -58.7028,
  -58.6303,
  -58.5567,
  -58.482,
  -58.4061,
  -58.3292,
  -58.2514,
  -58.1732,
  -58.0945,
  -58.0157,
  -57.9368,
  -57.858,
  -57.7793,
  -57.7004,
  -57.6214,
  -57.5423,
  -57.4629,
  -57.3835,
  -57.3042,
  -57.2252,
  -57.1462,
  -57.0669,
  -56.9874,
  -56.9067,
  -56.8268,
  -56.747,
  -56.6674,
  -56.5887,
  -56.5108,
  -56.4341,
  -56.3584,
  -56.2832,
  -56.2083,
  -56.1332,
  -56.0583,
  -55.9838,
  -55.9106,
  -55.8389,
  -55.7694,
  -55.7022,
  -55.6374,
  -55.5753,
  -55.5152,
  -55.4567,
  -55.3995,
  -55.3436,
  -55.2886,
  -55.2346,
  -55.1818,
  -55.1306,
  -55.081,
  -55.0337,
  -54.988,
  -54.9439,
  -54.9017,
  -54.8622,
  -54.8259,
  -54.7933,
  -54.7643,
  -54.7385,
  -54.7155,
  -54.695,
  -54.6766,
  -54.66,
  -54.645,
  -47.685,
  -47.5571,
  -47.4237,
  -47.2938,
  -47.1734,
  -47.0718,
  -46.9978,
  -46.9593,
  -46.9626,
  -47.0127,
  -47.1119,
  -47.2605,
  -47.4551,
  -47.688,
  -47.9527,
  -48.2388,
  -48.5363,
  -48.8362,
  -49.1307,
  -49.4139,
  -49.6823,
  -49.9339,
  -50.1694,
  -50.3892,
  -50.595,
  -50.7876,
  -50.9685,
  -51.1383,
  -51.297,
  -51.4475,
  -51.5897,
  -51.7243,
  -51.8522,
  -51.9741,
  -52.0906,
  -52.2024,
  -52.3095,
  -52.4127,
  -52.5118,
  -52.6064,
  -52.6967,
  -52.7822,
  -52.8634,
  -52.941,
  -53.0142,
  -53.0854,
  -53.1546,
  -53.2214,
  -53.2864,
  -53.3492,
  -53.4095,
  -53.4674,
  -53.5225,
  -53.5753,
  -53.6264,
  -53.6767,
  -53.7275,
  -53.7792,
  -53.8326,
  -53.8875,
  -53.9441,
  -54.0012,
  -54.0597,
  -54.1179,
  -54.1748,
  -54.2304,
  -54.2845,
  -54.3374,
  -54.3887,
  -54.4388,
  -54.4875,
  -54.5353,
  -54.5827,
  -54.6302,
  -54.6782,
  -54.727,
  -54.7768,
  -54.8281,
  -54.8793,
  -54.9323,
  -54.9861,
  -55.0401,
  -55.0941,
  -55.1477,
  -55.2007,
  -55.2533,
  -55.3048,
  -55.3556,
  -55.4056,
  -55.4544,
  -55.502,
  -55.5483,
  -55.5931,
  -55.6368,
  -55.6793,
  -55.7205,
  -55.7599,
  -55.7998,
  -55.8393,
  -55.8787,
  -55.9181,
  -55.9579,
  -55.9988,
  -56.0414,
  -56.0865,
  -56.1345,
  -56.1868,
  -56.244,
  -56.3075,
  -56.3775,
  -56.4537,
  -56.5352,
  -56.6204,
  -56.7077,
  -56.7951,
  -56.8809,
  -56.9624,
  -57.0412,
  -57.1159,
  -57.1865,
  -57.2535,
  -57.3176,
  -57.3796,
  -57.44,
  -57.4987,
  -57.556,
  -57.6113,
  -57.6646,
  -57.7157,
  -57.7646,
  -57.812,
  -57.8583,
  -57.9044,
  -57.9509,
  -57.9976,
  -58.0443,
  -58.0901,
  -58.1343,
  -58.1786,
  -58.2226,
  -58.2662,
  -58.3094,
  -58.3521,
  -58.3942,
  -58.4365,
  -58.4794,
  -58.5229,
  -58.5674,
  -58.6128,
  -58.6584,
  -58.7044,
  -58.7509,
  -58.7986,
  -58.8472,
  -58.8971,
  -58.9482,
  -58.9994,
  -59.051,
  -59.1023,
  -59.1524,
  -59.2037,
  -59.2554,
  -59.3079,
  -59.3615,
  -59.4161,
  -59.4717,
  -59.5283,
  -59.5853,
  -59.6426,
  -59.6998,
  -59.7563,
  -59.8115,
  -59.865,
  -59.9167,
  -59.9667,
  -60.015,
  -60.0617,
  -60.1063,
  -60.1483,
  -60.1877,
  -60.225,
  -60.2606,
  -60.2949,
  -60.3281,
  -60.3589,
  -60.3893,
  -60.4178,
  -60.4438,
  -60.4673,
  -60.4885,
  -60.508,
  -60.5261,
  -60.5434,
  -60.5597,
  -60.5741,
  -60.5863,
  -60.5956,
  -60.6018,
  -60.6044,
  -60.6034,
  -60.5991,
  -60.5914,
  -60.5814,
  -60.5694,
  -60.5556,
  -60.5401,
  -60.5229,
  -60.5046,
  -60.4849,
  -60.4636,
  -60.4403,
  -60.4145,
  -60.3862,
  -60.3545,
  -60.3213,
  -60.2856,
  -60.2472,
  -60.206,
  -60.1624,
  -60.1166,
  -60.0689,
  -60.0192,
  -59.9673,
  -59.9125,
  -59.8545,
  -59.7934,
  -59.7293,
  -59.6632,
  -59.5957,
  -59.5273,
  -59.4587,
  -59.3898,
  -59.3208,
  -59.2514,
  -59.1815,
  -59.1108,
  -59.0392,
  -58.966,
  -58.8916,
  -58.8158,
  -58.7384,
  -58.6598,
  -58.5804,
  -58.5005,
  -58.4202,
  -58.3398,
  -58.2584,
  -58.1781,
  -58.0979,
  -58.0178,
  -57.9378,
  -57.8578,
  -57.7779,
  -57.6981,
  -57.6185,
  -57.5386,
  -57.4584,
  -57.3777,
  -57.2964,
  -57.2147,
  -57.1328,
  -57.0508,
  -56.9691,
  -56.8879,
  -56.8077,
  -56.7288,
  -56.6508,
  -56.5737,
  -56.497,
  -56.4205,
  -56.3442,
  -56.2685,
  -56.1937,
  -56.1205,
  -56.0493,
  -55.9806,
  -55.9143,
  -55.851,
  -55.7895,
  -55.7303,
  -55.6723,
  -55.6153,
  -55.5593,
  -55.5043,
  -55.4504,
  -55.3983,
  -55.348,
  -55.2988,
  -55.2523,
  -55.2078,
  -55.1649,
  -55.1245,
  -55.0872,
  -55.0534,
  -55.0232,
  -54.9963,
  -54.9722,
  -54.9505,
  -54.9309,
  -54.9129,
  -54.8962,
  -47.6052,
  -47.4684,
  -47.3313,
  -47.2011,
  -47.0857,
  -46.9932,
  -46.9308,
  -46.9044,
  -46.9182,
  -46.9772,
  -47.0822,
  -47.2329,
  -47.4267,
  -47.6591,
  -47.923,
  -48.21,
  -48.5108,
  -48.8167,
  -49.1195,
  -49.413,
  -49.6928,
  -49.9567,
  -50.2045,
  -50.4356,
  -50.6525,
  -50.8555,
  -51.0454,
  -51.2235,
  -51.3905,
  -51.548,
  -51.6972,
  -51.8385,
  -51.973,
  -52.1013,
  -52.2241,
  -52.342,
  -52.455,
  -52.5636,
  -52.6666,
  -52.7658,
  -52.8602,
  -52.9493,
  -53.0339,
  -53.1144,
  -53.1919,
  -53.2671,
  -53.34,
  -53.4109,
  -53.4798,
  -53.5463,
  -53.6099,
  -53.6707,
  -53.7287,
  -53.7842,
  -53.8379,
  -53.8896,
  -53.9427,
  -53.9968,
  -54.0523,
  -54.1096,
  -54.1687,
  -54.2293,
  -54.2907,
  -54.3518,
  -54.4119,
  -54.4707,
  -54.5281,
  -54.584,
  -54.6387,
  -54.6919,
  -54.7439,
  -54.795,
  -54.8446,
  -54.895,
  -54.9457,
  -54.997,
  -55.0491,
  -55.1021,
  -55.1557,
  -55.2099,
  -55.2644,
  -55.3191,
  -55.374,
  -55.4285,
  -55.4826,
  -55.5366,
  -55.59,
  -55.643,
  -55.6955,
  -55.7472,
  -55.797,
  -55.8468,
  -55.8953,
  -55.9428,
  -55.9889,
  -56.0342,
  -56.0784,
  -56.1215,
  -56.1636,
  -56.2048,
  -56.2458,
  -56.2866,
  -56.3282,
  -56.3707,
  -56.415,
  -56.462,
  -56.512,
  -56.5672,
  -56.6278,
  -56.6936,
  -56.7669,
  -56.8461,
  -56.93,
  -57.0165,
  -57.1038,
  -57.19,
  -57.2735,
  -57.3536,
  -57.4295,
  -57.5014,
  -57.5699,
  -57.6355,
  -57.699,
  -57.7606,
  -57.8206,
  -57.879,
  -57.9356,
  -57.9901,
  -58.042,
  -58.0904,
  -58.138,
  -58.1847,
  -58.2311,
  -58.2777,
  -58.3245,
  -58.3711,
  -58.4171,
  -58.4626,
  -58.5076,
  -58.5521,
  -58.5965,
  -58.6405,
  -58.6841,
  -58.7276,
  -58.7715,
  -58.8163,
  -58.8621,
  -58.9086,
  -58.9558,
  -59.0032,
  -59.0507,
  -59.0975,
  -59.1457,
  -59.1945,
  -59.244,
  -59.2942,
  -59.3446,
  -59.395,
  -59.4452,
  -59.4953,
  -59.5455,
  -59.596,
  -59.6474,
  -59.6999,
  -59.7538,
  -59.809,
  -59.8655,
  -59.9226,
  -59.9803,
  -60.038,
  -60.0951,
  -60.1508,
  -60.2047,
  -60.2566,
  -60.3065,
  -60.3537,
  -60.3998,
  -60.4435,
  -60.4843,
  -60.5223,
  -60.5582,
  -60.5923,
  -60.6252,
  -60.657,
  -60.6874,
  -60.7164,
  -60.7435,
  -60.7684,
  -60.791,
  -60.8116,
  -60.8307,
  -60.8488,
  -60.8655,
  -60.8818,
  -60.896,
  -60.9078,
  -60.9167,
  -60.9223,
  -60.9241,
  -60.9221,
  -60.9164,
  -60.9072,
  -60.8942,
  -60.8802,
  -60.8645,
  -60.8476,
  -60.8295,
  -60.8107,
  -60.7908,
  -60.7695,
  -60.7461,
  -60.7201,
  -60.6913,
  -60.6601,
  -60.6265,
  -60.5906,
  -60.5524,
  -60.5118,
  -60.469,
  -60.4246,
  -60.3786,
  -60.3311,
  -60.2817,
  -60.2295,
  -60.1741,
  -60.1157,
  -60.0542,
  -59.9905,
  -59.9251,
  -59.8585,
  -59.7911,
  -59.7234,
  -59.6551,
  -59.5855,
  -59.5163,
  -59.4462,
  -59.3749,
  -59.302,
  -59.2271,
  -59.1507,
  -59.0724,
  -58.9927,
  -58.9119,
  -58.8304,
  -58.7485,
  -58.6667,
  -58.5848,
  -58.503,
  -58.4213,
  -58.3397,
  -58.2583,
  -58.1773,
  -58.0968,
  -58.0167,
  -57.9366,
  -57.8561,
  -57.7748,
  -57.6927,
  -57.6098,
  -57.5264,
  -57.4428,
  -57.3591,
  -57.2755,
  -57.1925,
  -57.1103,
  -57.0292,
  -56.9494,
  -56.8703,
  -56.7919,
  -56.7139,
  -56.6364,
  -56.5583,
  -56.4822,
  -56.4073,
  -56.3344,
  -56.264,
  -56.1964,
  -56.1318,
  -56.0697,
  -56.0095,
  -55.9508,
  -55.8931,
  -55.8362,
  -55.7802,
  -55.7254,
  -55.6721,
  -55.6208,
  -55.5716,
  -55.5246,
  -55.4798,
  -55.4366,
  -55.3958,
  -55.3578,
  -55.3232,
  -55.2918,
  -55.2633,
  -55.2377,
  -55.2144,
  -55.1931,
  -55.1736,
  -55.1549,
  -47.5332,
  -47.3899,
  -47.2505,
  -47.122,
  -47.0138,
  -46.9317,
  -46.881,
  -46.8671,
  -46.8924,
  -46.9593,
  -47.0682,
  -47.2191,
  -47.4107,
  -47.6395,
  -47.8998,
  -48.1856,
  -48.4879,
  -48.7973,
  -49.1077,
  -49.411,
  -49.7023,
  -49.9792,
  -50.2398,
  -50.4842,
  -50.7128,
  -50.926,
  -51.1251,
  -51.3112,
  -51.4857,
  -51.6502,
  -51.8059,
  -51.9542,
  -52.0957,
  -52.2297,
  -52.3592,
  -52.4834,
  -52.6027,
  -52.7172,
  -52.8266,
  -52.9306,
  -53.0294,
  -53.1224,
  -53.2108,
  -53.295,
  -53.3762,
  -53.4549,
  -53.5318,
  -53.6068,
  -53.6797,
  -53.7491,
  -53.8164,
  -53.8804,
  -53.9413,
  -53.9998,
  -54.0565,
  -54.1123,
  -54.1681,
  -54.2246,
  -54.2826,
  -54.3422,
  -54.4036,
  -54.4666,
  -54.5306,
  -54.5944,
  -54.6573,
  -54.7178,
  -54.7781,
  -54.8368,
  -54.8944,
  -54.9507,
  -55.0059,
  -55.06,
  -55.1136,
  -55.167,
  -55.2205,
  -55.2743,
  -55.3284,
  -55.3829,
  -55.4379,
  -55.493,
  -55.5485,
  -55.604,
  -55.6598,
  -55.7146,
  -55.7701,
  -55.8256,
  -55.8807,
  -55.936,
  -55.9911,
  -56.0456,
  -56.0993,
  -56.1525,
  -56.2045,
  -56.2556,
  -56.3056,
  -56.3546,
  -56.4021,
  -56.4485,
  -56.4936,
  -56.5374,
  -56.5804,
  -56.6228,
  -56.6644,
  -56.7077,
  -56.7523,
  -56.7988,
  -56.8478,
  -56.9011,
  -56.9593,
  -57.0235,
  -57.094,
  -57.1706,
  -57.2524,
  -57.3376,
  -57.4242,
  -57.5102,
  -57.594,
  -57.6747,
  -57.7517,
  -57.8248,
  -57.8946,
  -57.9604,
  -58.0249,
  -58.0876,
  -58.1488,
  -58.2085,
  -58.2662,
  -58.3214,
  -58.3739,
  -58.4237,
  -58.4715,
  -58.5184,
  -58.5649,
  -58.6114,
  -58.6579,
  -58.7043,
  -58.7504,
  -58.7962,
  -58.842,
  -58.8875,
  -58.9327,
  -58.9777,
  -59.0226,
  -59.0666,
  -59.1124,
  -59.1591,
  -59.2069,
  -59.2555,
  -59.3046,
  -59.3537,
  -59.4028,
  -59.4517,
  -59.5006,
  -59.5496,
  -59.5989,
  -59.6483,
  -59.6979,
  -59.7479,
  -59.7971,
  -59.8468,
  -59.8966,
  -59.9464,
  -59.9969,
  -60.0484,
  -60.1012,
  -60.1553,
  -60.2097,
  -60.266,
  -60.3228,
  -60.3797,
  -60.4362,
  -60.4915,
  -60.545,
  -60.5965,
  -60.646,
  -60.6937,
  -60.7388,
  -60.7815,
  -60.8212,
  -60.8581,
  -60.8927,
  -60.9254,
  -60.957,
  -60.9872,
  -61.016,
  -61.0432,
  -61.0685,
  -61.0919,
  -61.1134,
  -61.1333,
  -61.1518,
  -61.1689,
  -61.1842,
  -61.1993,
  -61.2122,
  -61.2229,
  -61.2304,
  -61.2347,
  -61.2355,
  -61.2324,
  -61.2254,
  -61.2148,
  -61.2013,
  -61.1857,
  -61.1686,
  -61.1505,
  -61.1315,
  -61.112,
  -61.0916,
  -61.0698,
  -61.0457,
  -61.019,
  -60.9897,
  -60.9579,
  -60.9238,
  -60.8876,
  -60.8493,
  -60.8091,
  -60.7672,
  -60.724,
  -60.6797,
  -60.6331,
  -60.5859,
  -60.5361,
  -60.4833,
  -60.4274,
  -60.3687,
  -60.3077,
  -60.2449,
  -60.1806,
  -60.1153,
  -60.0492,
  -59.9825,
  -59.9153,
  -59.8474,
  -59.7787,
  -59.7085,
  -59.6365,
  -59.5622,
  -59.4857,
  -59.4071,
  -59.3267,
  -59.2451,
  -59.1625,
  -59.0794,
  -58.9961,
  -58.9129,
  -58.8298,
  -58.7467,
  -58.6636,
  -58.5808,
  -58.4986,
  -58.4172,
  -58.3365,
  -58.2559,
  -58.1747,
  -58.0915,
  -58.0081,
  -57.924,
  -57.8392,
  -57.7541,
  -57.669,
  -57.5838,
  -57.4992,
  -57.4156,
  -57.333,
  -57.2515,
  -57.1709,
  -57.0911,
  -57.0118,
  -56.933,
  -56.8547,
  -56.7772,
  -56.7009,
  -56.6264,
  -56.5545,
  -56.4857,
  -56.42,
  -56.3568,
  -56.2957,
  -56.2363,
  -56.1778,
  -56.1201,
  -56.0633,
  -56.0077,
  -55.9535,
  -55.9013,
  -55.8512,
  -55.8038,
  -55.7589,
  -55.7158,
  -55.6751,
  -55.6368,
  -55.6014,
  -55.5688,
  -55.5389,
  -55.5114,
  -55.486,
  -55.4627,
  -55.441,
  -55.4202,
  -47.4722,
  -47.3246,
  -47.1852,
  -47.0623,
  -46.9627,
  -46.8916,
  -46.8531,
  -46.8506,
  -46.8851,
  -46.958,
  -47.0694,
  -47.219,
  -47.4055,
  -47.6289,
  -47.8841,
  -48.1666,
  -48.4689,
  -48.7826,
  -49.0994,
  -49.4123,
  -49.7153,
  -50.0045,
  -50.2781,
  -50.535,
  -50.7751,
  -50.9984,
  -51.2064,
  -51.3995,
  -51.5814,
  -51.7528,
  -51.9155,
  -52.0708,
  -52.2192,
  -52.3614,
  -52.4976,
  -52.6287,
  -52.7545,
  -52.875,
  -52.9902,
  -53.0996,
  -53.2031,
  -53.3008,
  -53.3934,
  -53.4808,
  -53.566,
  -53.6489,
  -53.7298,
  -53.8089,
  -53.8859,
  -53.9599,
  -54.0309,
  -54.0987,
  -54.1631,
  -54.2248,
  -54.2846,
  -54.3435,
  -54.4023,
  -54.4616,
  -54.5223,
  -54.5835,
  -54.6473,
  -54.7126,
  -54.7788,
  -54.8449,
  -54.9104,
  -54.9743,
  -55.0367,
  -55.098,
  -55.1583,
  -55.2172,
  -55.2753,
  -55.3326,
  -55.3889,
  -55.4452,
  -55.5011,
  -55.5571,
  -55.613,
  -55.6681,
  -55.7244,
  -55.7804,
  -55.8368,
  -55.8936,
  -55.9507,
  -56.0079,
  -56.065,
  -56.1221,
  -56.1792,
  -56.2365,
  -56.2938,
  -56.3506,
  -56.4071,
  -56.4633,
  -56.5185,
  -56.573,
  -56.6266,
  -56.6781,
  -56.7293,
  -56.7792,
  -56.8275,
  -56.8741,
  -56.9197,
  -56.9643,
  -57.0087,
  -57.0534,
  -57.0985,
  -57.1452,
  -57.194,
  -57.2462,
  -57.3028,
  -57.3648,
  -57.4329,
  -57.5071,
  -57.5867,
  -57.6702,
  -57.7543,
  -57.8394,
  -57.9231,
  -58.0041,
  -58.0818,
  -58.1557,
  -58.2262,
  -58.2939,
  -58.3592,
  -58.4226,
  -58.4845,
  -58.5451,
  -58.6037,
  -58.6598,
  -58.713,
  -58.7632,
  -58.8115,
  -58.8586,
  -58.9053,
  -58.9517,
  -58.9979,
  -59.0431,
  -59.0893,
  -59.1356,
  -59.1821,
  -59.2286,
  -59.2751,
  -59.3215,
  -59.3678,
  -59.4145,
  -59.4621,
  -59.5109,
  -59.5606,
  -59.6111,
  -59.6619,
  -59.7125,
  -59.7627,
  -59.8126,
  -59.8621,
  -59.9114,
  -59.9606,
  -60.0096,
  -60.0591,
  -60.1068,
  -60.1562,
  -60.206,
  -60.2557,
  -60.3052,
  -60.355,
  -60.4054,
  -60.4567,
  -60.5091,
  -60.5624,
  -60.6166,
  -60.6717,
  -60.7264,
  -60.7812,
  -60.8348,
  -60.887,
  -60.9375,
  -60.9862,
  -61.0327,
  -61.077,
  -61.1185,
  -61.1572,
  -61.1931,
  -61.2266,
  -61.2583,
  -61.2875,
  -61.3161,
  -61.3431,
  -61.3683,
  -61.3916,
  -61.4131,
  -61.4332,
  -61.4519,
  -61.4693,
  -61.4856,
  -61.5005,
  -61.5136,
  -61.5247,
  -61.5334,
  -61.5391,
  -61.5417,
  -61.5409,
  -61.5363,
  -61.5279,
  -61.5162,
  -61.5017,
  -61.485,
  -61.4669,
  -61.4477,
  -61.428,
  -61.4076,
  -61.3864,
  -61.3635,
  -61.3375,
  -61.3099,
  -61.2796,
  -61.2472,
  -61.2125,
  -61.1759,
  -61.1375,
  -61.0975,
  -61.0561,
  -61.0138,
  -60.9708,
  -60.9269,
  -60.8814,
  -60.8336,
  -60.7828,
  -60.7291,
  -60.6729,
  -60.6148,
  -60.5549,
  -60.4933,
  -60.4304,
  -60.3665,
  -60.3019,
  -60.2368,
  -60.1708,
  -60.1039,
  -60.0355,
  -59.9649,
  -59.8919,
  -59.8162,
  -59.7381,
  -59.6578,
  -59.5749,
  -59.4918,
  -59.4078,
  -59.3236,
  -59.2394,
  -59.1553,
  -59.0709,
  -58.9865,
  -58.9023,
  -58.8189,
  -58.7364,
  -58.6549,
  -58.5735,
  -58.4916,
  -58.4085,
  -58.3243,
  -58.2391,
  -58.1532,
  -58.067,
  -57.9806,
  -57.8942,
  -57.8085,
  -57.7238,
  -57.6401,
  -57.5574,
  -57.4757,
  -57.3948,
  -57.3144,
  -57.2345,
  -57.1551,
  -57.0763,
  -56.9988,
  -56.9229,
  -56.8497,
  -56.7795,
  -56.7124,
  -56.6481,
  -56.5862,
  -56.5259,
  -56.4667,
  -56.4082,
  -56.3497,
  -56.2933,
  -56.2385,
  -56.1856,
  -56.1353,
  -56.0878,
  -56.0429,
  -56.0002,
  -55.9598,
  -55.9213,
  -55.8853,
  -55.8517,
  -55.8202,
  -55.7908,
  -55.7634,
  -55.7379,
  -55.7141,
  -55.6913,
  -47.4285,
  -47.2789,
  -47.1417,
  -47.0243,
  -46.9334,
  -46.8729,
  -46.8459,
  -46.8524,
  -46.8951,
  -46.9725,
  -47.085,
  -47.2321,
  -47.414,
  -47.6306,
  -47.8797,
  -48.1575,
  -48.4582,
  -48.7738,
  -49.0964,
  -49.418,
  -49.732,
  -50.0334,
  -50.3183,
  -50.5871,
  -50.8382,
  -51.0717,
  -51.2884,
  -51.4904,
  -51.6796,
  -51.8582,
  -52.028,
  -52.1904,
  -52.3461,
  -52.4956,
  -52.6391,
  -52.7771,
  -52.9097,
  -53.0355,
  -53.1566,
  -53.2715,
  -53.3803,
  -53.483,
  -53.5806,
  -53.6738,
  -53.7638,
  -53.8512,
  -53.9366,
  -54.0198,
  -54.1008,
  -54.179,
  -54.2539,
  -54.3251,
  -54.3931,
  -54.4574,
  -54.5206,
  -54.5827,
  -54.6447,
  -54.707,
  -54.7705,
  -54.8354,
  -54.9019,
  -54.9695,
  -55.0377,
  -55.1059,
  -55.1734,
  -55.2395,
  -55.3039,
  -55.3671,
  -55.4295,
  -55.491,
  -55.5507,
  -55.6105,
  -55.6695,
  -55.728,
  -55.7861,
  -55.8439,
  -55.9016,
  -55.9591,
  -56.0164,
  -56.0738,
  -56.1314,
  -56.1895,
  -56.2482,
  -56.3071,
  -56.366,
  -56.4249,
  -56.4839,
  -56.5428,
  -56.601,
  -56.66,
  -56.7189,
  -56.7776,
  -56.8357,
  -56.8934,
  -56.9504,
  -57.0065,
  -57.0614,
  -57.1147,
  -57.1664,
  -57.2164,
  -57.2648,
  -57.3122,
  -57.3587,
  -57.405,
  -57.4515,
  -57.4989,
  -57.5481,
  -57.5989,
  -57.6546,
  -57.7152,
  -57.7815,
  -57.8537,
  -57.9311,
  -58.0124,
  -58.096,
  -58.18,
  -58.263,
  -58.3436,
  -58.4212,
  -58.4954,
  -58.5662,
  -58.6342,
  -58.6996,
  -58.7634,
  -58.826,
  -58.8873,
  -58.9468,
  -59.0027,
  -59.0567,
  -59.1079,
  -59.1571,
  -59.205,
  -59.2519,
  -59.2985,
  -59.3447,
  -59.3908,
  -59.4372,
  -59.4839,
  -59.5312,
  -59.5789,
  -59.6268,
  -59.6748,
  -59.7229,
  -59.7714,
  -59.8208,
  -59.8713,
  -59.9229,
  -59.975,
  -60.0271,
  -60.0778,
  -60.1289,
  -60.1794,
  -60.2295,
  -60.2791,
  -60.3284,
  -60.3774,
  -60.4264,
  -60.4755,
  -60.525,
  -60.5748,
  -60.6244,
  -60.6736,
  -60.7225,
  -60.7716,
  -60.8211,
  -60.8712,
  -60.9218,
  -60.973,
  -61.0246,
  -61.0765,
  -61.1282,
  -61.1794,
  -61.2294,
  -61.2769,
  -61.3239,
  -61.369,
  -61.4119,
  -61.4523,
  -61.49,
  -61.5251,
  -61.558,
  -61.5888,
  -61.6178,
  -61.645,
  -61.6702,
  -61.6933,
  -61.7146,
  -61.7342,
  -61.7525,
  -61.7696,
  -61.7855,
  -61.8001,
  -61.813,
  -61.8239,
  -61.8326,
  -61.8387,
  -61.8421,
  -61.8424,
  -61.8396,
  -61.8324,
  -61.8228,
  -61.8102,
  -61.7949,
  -61.7775,
  -61.7587,
  -61.7387,
  -61.7181,
  -61.6968,
  -61.6744,
  -61.6503,
  -61.624,
  -61.5953,
  -61.5641,
  -61.5307,
  -61.4953,
  -61.4583,
  -61.4197,
  -61.3797,
  -61.3387,
  -61.297,
  -61.2549,
  -61.212,
  -61.1677,
  -61.1212,
  -61.072,
  -61.0202,
  -60.9663,
  -60.9104,
  -60.853,
  -60.7942,
  -60.733,
  -60.6718,
  -60.6097,
  -60.5469,
  -60.4833,
  -60.4186,
  -60.3522,
  -60.2835,
  -60.2121,
  -60.1379,
  -60.061,
  -59.9817,
  -59.9002,
  -59.8171,
  -59.7331,
  -59.6485,
  -59.5638,
  -59.4789,
  -59.3936,
  -59.3081,
  -59.2228,
  -59.1383,
  -59.0548,
  -58.9723,
  -58.89,
  -58.8074,
  -58.7236,
  -58.6387,
  -58.5528,
  -58.4661,
  -58.3789,
  -58.2915,
  -58.2041,
  -58.1175,
  -58.0319,
  -57.9474,
  -57.864,
  -57.7805,
  -57.6988,
  -57.6176,
  -57.5368,
  -57.4564,
  -57.3766,
  -57.298,
  -57.2211,
  -57.1466,
  -57.0751,
  -57.0066,
  -56.9411,
  -56.8779,
  -56.8167,
  -56.7567,
  -56.6977,
  -56.6397,
  -56.5828,
  -56.5276,
  -56.4747,
  -56.4244,
  -56.3769,
  -56.3321,
  -56.2898,
  -56.2494,
  -56.2109,
  -56.1744,
  -56.1398,
  -56.107,
  -56.0761,
  -56.0469,
  -56.0194,
  -55.9933,
  -55.9682,
  -47.4047,
  -47.2543,
  -47.1212,
  -47.0108,
  -46.9288,
  -46.8785,
  -46.8614,
  -46.8776,
  -46.9262,
  -47.0066,
  -47.1184,
  -47.2618,
  -47.4374,
  -47.6461,
  -47.8877,
  -48.1597,
  -48.4566,
  -48.7729,
  -49.0999,
  -49.4291,
  -49.7531,
  -50.0656,
  -50.363,
  -50.6429,
  -50.9045,
  -51.1476,
  -51.3731,
  -51.583,
  -51.7799,
  -51.9659,
  -52.143,
  -52.3117,
  -52.4748,
  -52.6318,
  -52.7829,
  -52.928,
  -53.0676,
  -53.2008,
  -53.3279,
  -53.4486,
  -53.5631,
  -53.6715,
  -53.7746,
  -53.8732,
  -53.9682,
  -54.0606,
  -54.1507,
  -54.2376,
  -54.3225,
  -54.4046,
  -54.4834,
  -54.5584,
  -54.6304,
  -54.6995,
  -54.7665,
  -54.8321,
  -54.8973,
  -54.9628,
  -55.0293,
  -55.097,
  -55.166,
  -55.2361,
  -55.3065,
  -55.3766,
  -55.4447,
  -55.5126,
  -55.5789,
  -55.644,
  -55.7079,
  -55.7715,
  -55.8342,
  -55.896,
  -55.9572,
  -56.0179,
  -56.0778,
  -56.1371,
  -56.196,
  -56.2544,
  -56.3129,
  -56.3715,
  -56.4308,
  -56.4905,
  -56.55,
  -56.611,
  -56.6719,
  -56.7327,
  -56.7934,
  -56.8541,
  -56.9148,
  -56.9755,
  -57.0361,
  -57.0971,
  -57.158,
  -57.2186,
  -57.279,
  -57.3386,
  -57.397,
  -57.4539,
  -57.509,
  -57.5623,
  -57.6128,
  -57.663,
  -57.7122,
  -57.7608,
  -57.8091,
  -57.8577,
  -57.9079,
  -57.9601,
  -58.0158,
  -58.0759,
  -58.1409,
  -58.2113,
  -58.2865,
  -58.3657,
  -58.4474,
  -58.53,
  -58.6119,
  -58.6918,
  -58.7691,
  -58.843,
  -58.9124,
  -58.9798,
  -59.0449,
  -59.1087,
  -59.1717,
  -59.2334,
  -59.2935,
  -59.3513,
  -59.4066,
  -59.4587,
  -59.5091,
  -59.5582,
  -59.6061,
  -59.6532,
  -59.6998,
  -59.7463,
  -59.793,
  -59.8403,
  -59.8886,
  -59.9377,
  -59.9871,
  -60.0357,
  -60.0856,
  -60.136,
  -60.1871,
  -60.2394,
  -60.2924,
  -60.3459,
  -60.399,
  -60.4512,
  -60.5027,
  -60.5535,
  -60.6039,
  -60.6537,
  -60.7032,
  -60.7524,
  -60.8018,
  -60.8511,
  -60.9009,
  -60.9509,
  -61.0004,
  -61.0491,
  -61.0971,
  -61.1445,
  -61.1908,
  -61.238,
  -61.2852,
  -61.3323,
  -61.3796,
  -61.4273,
  -61.4751,
  -61.523,
  -61.5697,
  -61.6156,
  -61.6602,
  -61.7034,
  -61.7444,
  -61.7834,
  -61.8203,
  -61.8548,
  -61.8872,
  -61.9175,
  -61.9457,
  -61.9717,
  -61.9954,
  -62.0167,
  -62.0357,
  -62.0532,
  -62.0696,
  -62.0842,
  -62.0982,
  -62.1108,
  -62.1215,
  -62.1298,
  -62.1355,
  -62.1386,
  -62.1391,
  -62.1368,
  -62.1316,
  -62.1234,
  -62.1127,
  -62.0993,
  -62.0837,
  -62.066,
  -62.0467,
  -62.0261,
  -62.0046,
  -61.9821,
  -61.9582,
  -61.9326,
  -61.9048,
  -61.8747,
  -61.8425,
  -61.8083,
  -61.7722,
  -61.7346,
  -61.6956,
  -61.6557,
  -61.6139,
  -61.5727,
  -61.531,
  -61.4887,
  -61.445,
  -61.3992,
  -61.3508,
  -61.3001,
  -61.2475,
  -61.1935,
  -61.1384,
  -61.082,
  -61.0243,
  -60.9654,
  -60.906,
  -60.8456,
  -60.7848,
  -60.7226,
  -60.6585,
  -60.5921,
  -60.5228,
  -60.4508,
  -60.3758,
  -60.298,
  -60.2176,
  -60.1353,
  -60.0518,
  -59.9676,
  -59.883,
  -59.7978,
  -59.7118,
  -59.6256,
  -59.5394,
  -59.454,
  -59.3695,
  -59.285,
  -59.2019,
  -59.1183,
  -59.0339,
  -58.9485,
  -58.8622,
  -58.775,
  -58.6871,
  -58.5987,
  -58.5106,
  -58.4232,
  -58.337,
  -58.2521,
  -58.1683,
  -58.0853,
  -58.0029,
  -57.921,
  -57.8393,
  -57.7582,
  -57.6774,
  -57.598,
  -57.5203,
  -57.445,
  -57.3724,
  -57.3027,
  -57.2359,
  -57.1716,
  -57.1095,
  -57.0487,
  -56.9891,
  -56.9306,
  -56.8733,
  -56.818,
  -56.765,
  -56.7148,
  -56.6675,
  -56.6229,
  -56.5807,
  -56.5404,
  -56.5018,
  -56.4649,
  -56.4295,
  -56.3956,
  -56.3634,
  -56.3316,
  -56.3023,
  -56.2741,
  -56.247,
  -47.4008,
  -47.2534,
  -47.125,
  -47.022,
  -46.9492,
  -46.9086,
  -46.9006,
  -46.924,
  -46.9774,
  -47.0593,
  -47.1693,
  -47.3071,
  -47.4755,
  -47.676,
  -47.9095,
  -48.1748,
  -48.4687,
  -48.7847,
  -49.1145,
  -49.4494,
  -49.7818,
  -50.104,
  -50.4115,
  -50.7015,
  -50.9726,
  -51.2245,
  -51.4576,
  -51.6758,
  -51.8806,
  -52.0744,
  -52.2595,
  -52.4371,
  -52.6081,
  -52.773,
  -52.9318,
  -53.0843,
  -53.2307,
  -53.3704,
  -53.5035,
  -53.6302,
  -53.7504,
  -53.8648,
  -53.9728,
  -54.0772,
  -54.1782,
  -54.2761,
  -54.3713,
  -54.4641,
  -54.5539,
  -54.6401,
  -54.7226,
  -54.8015,
  -54.8773,
  -54.9504,
  -55.0214,
  -55.0907,
  -55.1593,
  -55.2279,
  -55.2964,
  -55.3671,
  -55.4389,
  -55.5114,
  -55.5839,
  -55.6556,
  -55.7261,
  -55.7954,
  -55.8633,
  -55.9299,
  -55.9954,
  -56.0603,
  -56.1246,
  -56.188,
  -56.2507,
  -56.313,
  -56.3742,
  -56.4337,
  -56.4936,
  -56.5533,
  -56.6129,
  -56.6731,
  -56.734,
  -56.7958,
  -56.8585,
  -56.9215,
  -56.9845,
  -57.0472,
  -57.1099,
  -57.1721,
  -57.234,
  -57.2959,
  -57.3583,
  -57.4213,
  -57.4846,
  -57.5472,
  -57.6106,
  -57.6735,
  -57.7354,
  -57.7959,
  -57.8543,
  -57.9108,
  -57.9655,
  -58.0187,
  -58.0709,
  -58.1216,
  -58.1722,
  -58.2226,
  -58.274,
  -58.3275,
  -58.3839,
  -58.444,
  -58.5084,
  -58.5775,
  -58.6501,
  -58.7273,
  -58.807,
  -58.8878,
  -58.9682,
  -59.0469,
  -59.1231,
  -59.1954,
  -59.2646,
  -59.3311,
  -59.3958,
  -59.4595,
  -59.5227,
  -59.5854,
  -59.6466,
  -59.7061,
  -59.7628,
  -59.8169,
  -59.8695,
  -59.9202,
  -59.9691,
  -60.0161,
  -60.0631,
  -60.1097,
  -60.1568,
  -60.2049,
  -60.254,
  -60.3042,
  -60.355,
  -60.4065,
  -60.4582,
  -60.5105,
  -60.5633,
  -60.6169,
  -60.6713,
  -60.7255,
  -60.7792,
  -60.8318,
  -60.8835,
  -60.9343,
  -60.9848,
  -61.0347,
  -61.0845,
  -61.1332,
  -61.1828,
  -61.2325,
  -61.2823,
  -61.332,
  -61.3808,
  -61.4287,
  -61.4751,
  -61.5207,
  -61.5655,
  -61.6095,
  -61.6529,
  -61.6959,
  -61.7386,
  -61.7814,
  -61.8244,
  -61.8675,
  -61.9103,
  -61.9525,
  -61.994,
  -62.0345,
  -62.0735,
  -62.1108,
  -62.1464,
  -62.1802,
  -62.2113,
  -62.2412,
  -62.269,
  -62.2946,
  -62.3175,
  -62.3375,
  -62.355,
  -62.3707,
  -62.3853,
  -62.3987,
  -62.4106,
  -62.4207,
  -62.4287,
  -62.434,
  -62.4364,
  -62.4364,
  -62.4336,
  -62.4285,
  -62.4209,
  -62.4109,
  -62.3988,
  -62.3845,
  -62.3681,
  -62.3498,
  -62.33,
  -62.3083,
  -62.2858,
  -62.261,
  -62.2356,
  -62.2086,
  -62.1795,
  -62.1484,
  -62.1152,
  -62.0802,
  -62.0435,
  -62.0055,
  -61.9664,
  -61.9263,
  -61.8856,
  -61.8443,
  -61.8027,
  -61.7604,
  -61.7167,
  -61.6711,
  -61.6231,
  -61.5731,
  -61.5218,
  -61.4695,
  -61.416,
  -61.3614,
  -61.3058,
  -61.2491,
  -61.1914,
  -61.1335,
  -61.0752,
  -61.0152,
  -60.9533,
  -60.8889,
  -60.8217,
  -60.7507,
  -60.6778,
  -60.6019,
  -60.5233,
  -60.4425,
  -60.3602,
  -60.2768,
  -60.1928,
  -60.1077,
  -60.0218,
  -59.9353,
  -59.8488,
  -59.7629,
  -59.6778,
  -59.5935,
  -59.5095,
  -59.4252,
  -59.3403,
  -59.2544,
  -59.1677,
  -59.0802,
  -58.9919,
  -58.903,
  -58.8143,
  -58.7263,
  -58.6395,
  -58.5541,
  -58.4698,
  -58.3866,
  -58.3037,
  -58.2213,
  -58.1391,
  -58.0571,
  -57.9761,
  -57.8961,
  -57.8181,
  -57.742,
  -57.6684,
  -57.5976,
  -57.5296,
  -57.4633,
  -57.4001,
  -57.3387,
  -57.2785,
  -57.2195,
  -57.1621,
  -57.1067,
  -57.0539,
  -57.0038,
  -56.9565,
  -56.9119,
  -56.8695,
  -56.829,
  -56.7902,
  -56.7528,
  -56.7169,
  -56.6823,
  -56.649,
  -56.617,
  -56.5862,
  -56.5565,
  -56.5278,
  -47.4187,
  -47.2757,
  -47.1533,
  -47.0588,
  -46.9949,
  -46.9625,
  -46.9628,
  -46.9924,
  -47.0489,
  -47.1311,
  -47.2388,
  -47.3725,
  -47.5339,
  -47.7257,
  -47.9503,
  -48.208,
  -48.496,
  -48.8095,
  -49.1405,
  -49.4792,
  -49.8166,
  -50.1469,
  -50.463,
  -50.7616,
  -51.041,
  -51.3013,
  -51.5439,
  -51.7707,
  -51.984,
  -52.1865,
  -52.3802,
  -52.5663,
  -52.7456,
  -52.9187,
  -53.0852,
  -53.2452,
  -53.3973,
  -53.5434,
  -53.6827,
  -53.8151,
  -53.9414,
  -54.0617,
  -54.1768,
  -54.2876,
  -54.3946,
  -54.4986,
  -54.5996,
  -54.6979,
  -54.7926,
  -54.8834,
  -54.9701,
  -55.0532,
  -55.1322,
  -55.2092,
  -55.2842,
  -55.3574,
  -55.4296,
  -55.5016,
  -55.5741,
  -55.6476,
  -55.722,
  -55.7968,
  -55.8711,
  -55.9443,
  -56.0162,
  -56.0866,
  -56.1558,
  -56.2237,
  -56.2904,
  -56.3553,
  -56.4207,
  -56.4851,
  -56.549,
  -56.6121,
  -56.6746,
  -56.736,
  -56.7968,
  -56.8574,
  -56.9184,
  -56.9799,
  -57.0428,
  -57.1068,
  -57.1718,
  -57.237,
  -57.3022,
  -57.367,
  -57.4316,
  -57.4946,
  -57.5577,
  -57.6212,
  -57.6846,
  -57.7493,
  -57.815,
  -57.881,
  -57.9476,
  -58.0135,
  -58.0785,
  -58.1422,
  -58.2038,
  -58.2636,
  -58.3216,
  -58.3777,
  -58.4326,
  -58.4862,
  -58.5391,
  -58.5909,
  -58.6439,
  -58.6988,
  -58.7563,
  -58.817,
  -58.8816,
  -58.95,
  -59.0222,
  -59.0976,
  -59.1756,
  -59.2545,
  -59.3331,
  -59.4101,
  -59.484,
  -59.5546,
  -59.622,
  -59.6869,
  -59.7508,
  -59.8144,
  -59.8782,
  -59.9409,
  -60.0037,
  -60.065,
  -60.1238,
  -60.1807,
  -60.2355,
  -60.2881,
  -60.3389,
  -60.3879,
  -60.4357,
  -60.4829,
  -60.5304,
  -60.5791,
  -60.6291,
  -60.6802,
  -60.7323,
  -60.7852,
  -60.8386,
  -60.8923,
  -60.9467,
  -61.0017,
  -61.0567,
  -61.1106,
  -61.1646,
  -61.2174,
  -61.2691,
  -61.3198,
  -61.3699,
  -61.4199,
  -61.4699,
  -61.5198,
  -61.5698,
  -61.6197,
  -61.6693,
  -61.7179,
  -61.7658,
  -61.812,
  -61.8566,
  -61.9,
  -61.942,
  -61.9827,
  -62.0221,
  -62.0606,
  -62.0985,
  -62.136,
  -62.1736,
  -62.2103,
  -62.2482,
  -62.286,
  -62.3238,
  -62.3607,
  -62.3968,
  -62.432,
  -62.4657,
  -62.4988,
  -62.5309,
  -62.5609,
  -62.589,
  -62.6145,
  -62.6369,
  -62.6562,
  -62.6727,
  -62.6871,
  -62.6998,
  -62.711,
  -62.7206,
  -62.7282,
  -62.7328,
  -62.7349,
  -62.7342,
  -62.731,
  -62.7251,
  -62.716,
  -62.7059,
  -62.694,
  -62.6804,
  -62.665,
  -62.6479,
  -62.6287,
  -62.6075,
  -62.5852,
  -62.5612,
  -62.5357,
  -62.509,
  -62.4806,
  -62.4504,
  -62.4184,
  -62.3845,
  -62.3489,
  -62.3118,
  -62.2735,
  -62.2342,
  -62.1943,
  -62.1536,
  -62.1123,
  -62.0704,
  -62.0276,
  -61.9834,
  -61.9375,
  -61.8897,
  -61.8402,
  -61.7895,
  -61.737,
  -61.6847,
  -61.6312,
  -61.5769,
  -61.5215,
  -61.4657,
  -61.4097,
  -61.3531,
  -61.2949,
  -61.2347,
  -61.172,
  -61.1067,
  -61.0386,
  -60.9677,
  -60.8938,
  -60.8172,
  -60.7385,
  -60.658,
  -60.5761,
  -60.493,
  -60.4086,
  -60.3232,
  -60.2371,
  -60.151,
  -60.0652,
  -59.98,
  -59.8952,
  -59.8105,
  -59.7255,
  -59.6398,
  -59.5536,
  -59.4667,
  -59.3791,
  -59.2907,
  -59.2018,
  -59.1128,
  -59.0233,
  -58.9358,
  -58.8497,
  -58.7649,
  -58.6812,
  -58.5981,
  -58.5154,
  -58.4329,
  -58.351,
  -58.2698,
  -58.19,
  -58.1117,
  -58.0352,
  -57.9609,
  -57.8892,
  -57.8201,
  -57.7538,
  -57.6897,
  -57.6275,
  -57.5668,
  -57.5074,
  -57.4498,
  -57.3944,
  -57.3416,
  -57.2914,
  -57.244,
  -57.1991,
  -57.1563,
  -57.1155,
  -57.0763,
  -57.0385,
  -57.002,
  -56.9668,
  -56.9328,
  -56.8998,
  -56.8678,
  -56.8367,
  -56.8066,
  -47.457,
  -47.3191,
  -47.2045,
  -47.119,
  -47.0649,
  -47.0421,
  -47.0496,
  -47.0847,
  -47.1439,
  -47.226,
  -47.3308,
  -47.4589,
  -47.6127,
  -47.7956,
  -48.0112,
  -48.2596,
  -48.5411,
  -48.8501,
  -49.1799,
  -49.5203,
  -49.8623,
  -50.1976,
  -50.5199,
  -50.8253,
  -51.1117,
  -51.3797,
  -51.6306,
  -51.8661,
  -52.0887,
  -52.3009,
  -52.5033,
  -52.6988,
  -52.8872,
  -53.0686,
  -53.2431,
  -53.4104,
  -53.5703,
  -53.7227,
  -53.8677,
  -54.0061,
  -54.1381,
  -54.2644,
  -54.3858,
  -54.5029,
  -54.6166,
  -54.7268,
  -54.833,
  -54.9369,
  -55.0372,
  -55.1331,
  -55.2249,
  -55.3128,
  -55.3971,
  -55.4784,
  -55.5573,
  -55.6345,
  -55.7104,
  -55.7857,
  -55.8612,
  -55.9372,
  -56.0139,
  -56.0904,
  -56.1662,
  -56.2401,
  -56.313,
  -56.3844,
  -56.4544,
  -56.5234,
  -56.5912,
  -56.6578,
  -56.7238,
  -56.7889,
  -56.8533,
  -56.9172,
  -56.9803,
  -57.0427,
  -57.1043,
  -57.166,
  -57.2283,
  -57.2917,
  -57.3556,
  -57.4218,
  -57.489,
  -57.5565,
  -57.624,
  -57.6912,
  -57.7576,
  -57.8229,
  -57.8878,
  -57.9528,
  -58.0179,
  -58.0843,
  -58.1517,
  -58.2204,
  -58.2895,
  -58.3583,
  -58.4261,
  -58.4927,
  -58.5565,
  -58.6194,
  -58.6804,
  -58.7395,
  -58.7971,
  -58.8537,
  -58.9093,
  -58.9643,
  -59.0194,
  -59.0756,
  -59.1344,
  -59.1958,
  -59.2607,
  -59.3287,
  -59.3998,
  -59.4739,
  -59.5501,
  -59.6272,
  -59.7038,
  -59.7781,
  -59.8488,
  -59.9171,
  -59.9825,
  -60.0459,
  -60.1089,
  -60.1725,
  -60.2371,
  -60.3023,
  -60.367,
  -60.4304,
  -60.4923,
  -60.5522,
  -60.6097,
  -60.6649,
  -60.7174,
  -60.7676,
  -60.8161,
  -60.864,
  -60.912,
  -60.9613,
  -61.0119,
  -61.0629,
  -61.1159,
  -61.17,
  -61.2247,
  -61.2798,
  -61.3353,
  -61.391,
  -61.4466,
  -61.5017,
  -61.5556,
  -61.6084,
  -61.6599,
  -61.7106,
  -61.7603,
  -61.8099,
  -61.8595,
  -61.9092,
  -61.9588,
  -62.0083,
  -62.0567,
  -62.1044,
  -62.1505,
  -62.195,
  -62.2366,
  -62.2776,
  -62.3167,
  -62.354,
  -62.3895,
  -62.4235,
  -62.4565,
  -62.4889,
  -62.5209,
  -62.553,
  -62.5854,
  -62.6183,
  -62.6517,
  -62.685,
  -62.7182,
  -62.7508,
  -62.7828,
  -62.8149,
  -62.8461,
  -62.8764,
  -62.9046,
  -62.9299,
  -62.9522,
  -62.9712,
  -62.987,
  -62.9993,
  -63.0106,
  -63.0196,
  -63.0266,
  -63.0311,
  -63.0329,
  -63.0319,
  -63.0279,
  -63.0215,
  -63.0126,
  -63.0018,
  -62.9892,
  -62.9753,
  -62.9598,
  -62.943,
  -62.924,
  -62.9035,
  -62.8812,
  -62.8573,
  -62.8317,
  -62.8049,
  -62.7768,
  -62.7473,
  -62.7164,
  -62.6837,
  -62.6494,
  -62.6136,
  -62.5764,
  -62.5381,
  -62.4978,
  -62.4577,
  -62.4171,
  -62.3753,
  -62.3329,
  -62.2894,
  -62.2446,
  -62.1984,
  -62.1505,
  -62.1013,
  -62.0511,
  -62.0003,
  -61.9486,
  -61.8958,
  -61.8422,
  -61.7879,
  -61.7332,
  -61.6783,
  -61.6226,
  -61.5655,
  -61.5062,
  -61.4445,
  -61.3805,
  -61.3137,
  -61.2445,
  -61.1729,
  -61.0984,
  -61.0217,
  -60.9432,
  -60.8629,
  -60.7812,
  -60.6978,
  -60.6135,
  -60.5275,
  -60.4421,
  -60.3569,
  -60.2719,
  -60.187,
  -60.1018,
  -60.0163,
  -59.9301,
  -59.8435,
  -59.7564,
  -59.6689,
  -59.5806,
  -59.4918,
  -59.4028,
  -59.314,
  -59.2261,
  -59.1394,
  -59.0541,
  -58.9701,
  -58.887,
  -58.8043,
  -58.722,
  -58.6404,
  -58.5596,
  -58.48,
  -58.4018,
  -58.3251,
  -58.2504,
  -58.178,
  -58.1081,
  -58.0407,
  -57.9758,
  -57.9128,
  -57.8515,
  -57.7919,
  -57.7341,
  -57.6787,
  -57.6256,
  -57.5754,
  -57.5275,
  -57.4821,
  -57.4389,
  -57.3976,
  -57.3579,
  -57.3184,
  -57.2814,
  -57.2456,
  -57.2109,
  -57.1772,
  -57.1443,
  -57.1124,
  -57.0812,
  -47.5137,
  -47.3832,
  -47.2776,
  -47.2027,
  -47.1582,
  -47.1452,
  -47.16,
  -47.2002,
  -47.2618,
  -47.3439,
  -47.4447,
  -47.5676,
  -47.7142,
  -47.8883,
  -48.0945,
  -48.3349,
  -48.608,
  -48.9107,
  -49.2362,
  -49.5753,
  -49.918,
  -50.2559,
  -50.5821,
  -50.8923,
  -51.1847,
  -51.4582,
  -51.7171,
  -51.9617,
  -52.1944,
  -52.417,
  -52.6308,
  -52.8367,
  -53.0349,
  -53.2255,
  -53.4082,
  -53.5828,
  -53.7492,
  -53.9077,
  -54.0585,
  -54.2022,
  -54.3387,
  -54.4707,
  -54.5981,
  -54.7215,
  -54.8417,
  -54.9586,
  -55.0723,
  -55.1824,
  -55.2888,
  -55.3907,
  -55.4881,
  -55.5812,
  -55.6707,
  -55.7567,
  -55.8398,
  -55.9208,
  -56.0002,
  -56.0779,
  -56.1563,
  -56.2347,
  -56.3131,
  -56.391,
  -56.4681,
  -56.5437,
  -56.6177,
  -56.69,
  -56.7608,
  -56.8305,
  -56.8988,
  -56.9661,
  -57.0322,
  -57.0977,
  -57.1625,
  -57.2269,
  -57.2896,
  -57.3526,
  -57.4152,
  -57.478,
  -57.5417,
  -57.6069,
  -57.6738,
  -57.7422,
  -57.8117,
  -57.8815,
  -57.9513,
  -58.0205,
  -58.0888,
  -58.156,
  -58.2226,
  -58.2892,
  -58.3564,
  -58.4246,
  -58.4933,
  -58.5642,
  -58.6354,
  -58.7066,
  -58.7771,
  -58.8464,
  -58.9139,
  -58.9796,
  -59.0434,
  -59.1055,
  -59.1661,
  -59.2253,
  -59.2836,
  -59.3408,
  -59.3978,
  -59.4558,
  -59.5158,
  -59.5779,
  -59.643,
  -59.71,
  -59.7807,
  -59.8536,
  -59.9282,
  -60.0034,
  -60.0776,
  -60.1496,
  -60.2186,
  -60.2845,
  -60.3477,
  -60.4098,
  -60.4723,
  -60.5359,
  -60.6013,
  -60.6679,
  -60.7347,
  -60.801,
  -60.8658,
  -60.9287,
  -60.9891,
  -61.0458,
  -61.1005,
  -61.1525,
  -61.2022,
  -61.2507,
  -61.2993,
  -61.349,
  -61.4001,
  -61.4525,
  -61.5063,
  -61.5611,
  -61.6166,
  -61.6728,
  -61.729,
  -61.7851,
  -61.8406,
  -61.8955,
  -61.9492,
  -62.002,
  -62.0533,
  -62.1038,
  -62.153,
  -62.2007,
  -62.2495,
  -62.2982,
  -62.3468,
  -62.395,
  -62.442,
  -62.4879,
  -62.5322,
  -62.5747,
  -62.6151,
  -62.6535,
  -62.6897,
  -62.7235,
  -62.7553,
  -62.7854,
  -62.8138,
  -62.8409,
  -62.8674,
  -62.8938,
  -62.9205,
  -62.9482,
  -62.977,
  -63.0063,
  -63.0359,
  -63.0659,
  -63.0949,
  -63.1253,
  -63.1559,
  -63.1855,
  -63.2134,
  -63.2388,
  -63.2611,
  -63.2796,
  -63.2951,
  -63.3074,
  -63.3169,
  -63.3238,
  -63.328,
  -63.3296,
  -63.3284,
  -63.3242,
  -63.3175,
  -63.3081,
  -63.2966,
  -63.2832,
  -63.2683,
  -63.252,
  -63.2347,
  -63.2157,
  -63.1952,
  -63.173,
  -63.149,
  -63.1225,
  -63.0955,
  -63.0671,
  -63.0377,
  -63.0073,
  -62.9756,
  -62.9427,
  -62.9083,
  -62.8726,
  -62.8357,
  -62.7975,
  -62.7584,
  -62.7184,
  -62.6776,
  -62.6357,
  -62.5927,
  -62.5484,
  -62.503,
  -62.4562,
  -62.4083,
  -62.3593,
  -62.3095,
  -62.2588,
  -62.2072,
  -62.1548,
  -62.1014,
  -62.0477,
  -61.9936,
  -61.9389,
  -61.8835,
  -61.8265,
  -61.7664,
  -61.705,
  -61.6416,
  -61.5758,
  -61.5078,
  -61.4378,
  -61.3653,
  -61.2904,
  -61.2139,
  -61.1355,
  -61.0551,
  -60.9734,
  -60.8905,
  -60.807,
  -60.723,
  -60.6387,
  -60.5542,
  -60.4694,
  -60.384,
  -60.2982,
  -60.2117,
  -60.1248,
  -60.0375,
  -59.9499,
  -59.8621,
  -59.7737,
  -59.6851,
  -59.5965,
  -59.5084,
  -59.4213,
  -59.3357,
  -59.2516,
  -59.1685,
  -59.0861,
  -59.0044,
  -58.9233,
  -58.8433,
  -58.7645,
  -58.6868,
  -58.6094,
  -58.5345,
  -58.4616,
  -58.3909,
  -58.3226,
  -58.2567,
  -58.1929,
  -58.1311,
  -58.0711,
  -58.0133,
  -57.9577,
  -57.9044,
  -57.8535,
  -57.8048,
  -57.7587,
  -57.7149,
  -57.6732,
  -57.6326,
  -57.5934,
  -57.5557,
  -57.5191,
  -57.4838,
  -57.4496,
  -57.4163,
  -57.3838,
  -57.352,
  -47.5876,
  -47.4663,
  -47.3714,
  -47.3073,
  -47.2732,
  -47.2699,
  -47.2921,
  -47.3373,
  -47.4013,
  -47.4831,
  -47.5822,
  -47.7004,
  -47.8405,
  -48.0065,
  -48.2033,
  -48.434,
  -48.6981,
  -48.9925,
  -49.3114,
  -49.6448,
  -49.9852,
  -50.3223,
  -50.6495,
  -50.9621,
  -51.2589,
  -51.5395,
  -51.8056,
  -52.0596,
  -52.3029,
  -52.5368,
  -52.7622,
  -52.9795,
  -53.1884,
  -53.3887,
  -53.58,
  -53.7611,
  -53.934,
  -54.098,
  -54.2541,
  -54.4027,
  -54.5451,
  -54.6824,
  -54.8155,
  -54.9449,
  -55.0714,
  -55.195,
  -55.3156,
  -55.4325,
  -55.5454,
  -55.6538,
  -55.7576,
  -55.8558,
  -55.9508,
  -56.0421,
  -56.1299,
  -56.2148,
  -56.2976,
  -56.3792,
  -56.4603,
  -56.5408,
  -56.6206,
  -56.6998,
  -56.7777,
  -56.8543,
  -56.9291,
  -57.0021,
  -57.0736,
  -57.1425,
  -57.2111,
  -57.2783,
  -57.3448,
  -57.4104,
  -57.4752,
  -57.5396,
  -57.6036,
  -57.6674,
  -57.7309,
  -57.795,
  -57.8603,
  -57.9273,
  -57.996,
  -58.0666,
  -58.1381,
  -58.2102,
  -58.2822,
  -58.3524,
  -58.4228,
  -58.4921,
  -58.5607,
  -58.6292,
  -58.6984,
  -58.7688,
  -58.8405,
  -58.9134,
  -58.9868,
  -59.0602,
  -59.1331,
  -59.2048,
  -59.2749,
  -59.3434,
  -59.4098,
  -59.4749,
  -59.5382,
  -59.6001,
  -59.6597,
  -59.7191,
  -59.7781,
  -59.8377,
  -59.8984,
  -59.9613,
  -60.0269,
  -60.0949,
  -60.1652,
  -60.2372,
  -60.3104,
  -60.3836,
  -60.4556,
  -60.5252,
  -60.5918,
  -60.6553,
  -60.717,
  -60.7783,
  -60.8402,
  -60.9037,
  -60.9687,
  -61.0366,
  -61.1055,
  -61.1742,
  -61.2418,
  -61.3077,
  -61.3708,
  -61.4314,
  -61.4883,
  -61.5418,
  -61.5928,
  -61.6425,
  -61.6919,
  -61.742,
  -61.7933,
  -61.8461,
  -61.9002,
  -61.9554,
  -62.0116,
  -62.0681,
  -62.1245,
  -62.1795,
  -62.2347,
  -62.2889,
  -62.3423,
  -62.3946,
  -62.4458,
  -62.4958,
  -62.5443,
  -62.5919,
  -62.6391,
  -62.6863,
  -62.733,
  -62.7791,
  -62.8243,
  -62.868,
  -62.9103,
  -62.9508,
  -62.9891,
  -63.025,
  -63.0584,
  -63.0893,
  -63.1175,
  -63.1438,
  -63.168,
  -63.1894,
  -63.2104,
  -63.2314,
  -63.2527,
  -63.2752,
  -63.2989,
  -63.324,
  -63.35,
  -63.3768,
  -63.4046,
  -63.4331,
  -63.4618,
  -63.4902,
  -63.5172,
  -63.5418,
  -63.5635,
  -63.5814,
  -63.5961,
  -63.6072,
  -63.6148,
  -63.6196,
  -63.6213,
  -63.6201,
  -63.616,
  -63.6091,
  -63.5996,
  -63.5868,
  -63.5728,
  -63.5571,
  -63.54,
  -63.5215,
  -63.502,
  -63.4809,
  -63.4583,
  -63.4342,
  -63.4085,
  -63.3813,
  -63.3527,
  -63.323,
  -63.2925,
  -63.2612,
  -63.2291,
  -63.196,
  -63.1618,
  -63.1266,
  -63.0901,
  -63.052,
  -63.0132,
  -62.9733,
  -62.9322,
  -62.8902,
  -62.8468,
  -62.8021,
  -62.7561,
  -62.7089,
  -62.6598,
  -62.6108,
  -62.5612,
  -62.5107,
  -62.459,
  -62.4064,
  -62.353,
  -62.2996,
  -62.2458,
  -62.1911,
  -62.1352,
  -62.0779,
  -62.0185,
  -61.9569,
  -61.8934,
  -61.8279,
  -61.7607,
  -61.6917,
  -61.6207,
  -61.5478,
  -61.4729,
  -61.3959,
  -61.3172,
  -61.2372,
  -61.1561,
  -61.0743,
  -60.9918,
  -60.9086,
  -60.8247,
  -60.7401,
  -60.6549,
  -60.5691,
  -60.4826,
  -60.3956,
  -60.3082,
  -60.2208,
  -60.1322,
  -60.0446,
  -59.9567,
  -59.8687,
  -59.7809,
  -59.694,
  -59.6086,
  -59.5245,
  -59.4414,
  -59.3593,
  -59.2781,
  -59.1978,
  -59.1186,
  -59.0406,
  -58.9637,
  -58.8879,
  -58.8133,
  -58.7402,
  -58.6691,
  -58.6001,
  -58.5334,
  -58.4689,
  -58.4067,
  -58.3466,
  -58.2887,
  -58.2329,
  -58.179,
  -58.1273,
  -58.0777,
  -58.0307,
  -57.9862,
  -57.9436,
  -57.9025,
  -57.8624,
  -57.8237,
  -57.7864,
  -57.7505,
  -57.7155,
  -57.6818,
  -57.649,
  -57.6166,
  -47.675,
  -47.5651,
  -47.4824,
  -47.4302,
  -47.4083,
  -47.4147,
  -47.4453,
  -47.4954,
  -47.5622,
  -47.6437,
  -47.7405,
  -47.8547,
  -47.9891,
  -48.1487,
  -48.3358,
  -48.5568,
  -48.8116,
  -49.0963,
  -49.4059,
  -49.7328,
  -50.0676,
  -50.4009,
  -50.7264,
  -51.0397,
  -51.339,
  -51.6244,
  -51.8977,
  -52.1607,
  -52.4147,
  -52.6595,
  -52.8971,
  -53.1264,
  -53.3466,
  -53.5571,
  -53.7573,
  -53.9469,
  -54.126,
  -54.2957,
  -54.4564,
  -54.6096,
  -54.7564,
  -54.8984,
  -55.0366,
  -55.1717,
  -55.3043,
  -55.4334,
  -55.5607,
  -55.6847,
  -55.8048,
  -55.9203,
  -56.031,
  -56.1369,
  -56.2384,
  -56.3353,
  -56.4281,
  -56.5173,
  -56.6036,
  -56.688,
  -56.7712,
  -56.8535,
  -56.9347,
  -57.0138,
  -57.0926,
  -57.1699,
  -57.2455,
  -57.3191,
  -57.3907,
  -57.4606,
  -57.5292,
  -57.5964,
  -57.6625,
  -57.7279,
  -57.7927,
  -57.8572,
  -57.9217,
  -57.9858,
  -58.0504,
  -58.1156,
  -58.1825,
  -58.2502,
  -58.3207,
  -58.3932,
  -58.4668,
  -58.5409,
  -58.6148,
  -58.688,
  -58.7604,
  -58.8319,
  -58.9026,
  -58.9732,
  -59.0443,
  -59.1168,
  -59.1907,
  -59.2656,
  -59.3411,
  -59.4165,
  -59.4917,
  -59.5648,
  -59.6375,
  -59.7084,
  -59.7776,
  -59.8452,
  -59.9113,
  -59.9757,
  -60.0387,
  -60.1001,
  -60.161,
  -60.2219,
  -60.2837,
  -60.3472,
  -60.4129,
  -60.4811,
  -60.5511,
  -60.6226,
  -60.6945,
  -60.7659,
  -60.8352,
  -60.9028,
  -60.9672,
  -61.029,
  -61.0895,
  -61.1498,
  -61.2112,
  -61.275,
  -61.3414,
  -61.4101,
  -61.4804,
  -61.5511,
  -61.6209,
  -61.6891,
  -61.7548,
  -61.8176,
  -61.8769,
  -61.9326,
  -61.9853,
  -62.0361,
  -62.086,
  -62.1355,
  -62.187,
  -62.2397,
  -62.2939,
  -62.3493,
  -62.4055,
  -62.4619,
  -62.5181,
  -62.5735,
  -62.6279,
  -62.6814,
  -62.7341,
  -62.786,
  -62.8367,
  -62.8858,
  -62.9334,
  -62.9798,
  -63.0253,
  -63.0705,
  -63.1148,
  -63.1585,
  -63.201,
  -63.2424,
  -63.2815,
  -63.3197,
  -63.356,
  -63.3896,
  -63.4206,
  -63.4487,
  -63.474,
  -63.4967,
  -63.517,
  -63.5349,
  -63.5511,
  -63.5671,
  -63.583,
  -63.6003,
  -63.6191,
  -63.6396,
  -63.6616,
  -63.6849,
  -63.7099,
  -63.736,
  -63.7623,
  -63.7883,
  -63.8133,
  -63.8364,
  -63.8567,
  -63.8723,
  -63.8855,
  -63.895,
  -63.9011,
  -63.9036,
  -63.9029,
  -63.8991,
  -63.8924,
  -63.883,
  -63.8713,
  -63.8573,
  -63.8412,
  -63.8233,
  -63.804,
  -63.7835,
  -63.7618,
  -63.7384,
  -63.7136,
  -63.6876,
  -63.6601,
  -63.6313,
  -63.6014,
  -63.5706,
  -63.539,
  -63.5069,
  -63.4744,
  -63.4413,
  -63.4074,
  -63.3716,
  -63.3355,
  -63.298,
  -63.2593,
  -63.2195,
  -63.1785,
  -63.1362,
  -63.0926,
  -63.0477,
  -63.0014,
  -62.9539,
  -62.9057,
  -62.8566,
  -62.807,
  -62.7562,
  -62.7045,
  -62.6519,
  -62.5989,
  -62.5453,
  -62.4912,
  -62.4361,
  -62.3796,
  -62.3217,
  -62.2616,
  -62.1998,
  -62.136,
  -62.0706,
  -62.0037,
  -61.9353,
  -61.8652,
  -61.7933,
  -61.7195,
  -61.6438,
  -61.5655,
  -61.487,
  -61.4077,
  -61.3276,
  -61.2466,
  -61.1646,
  -61.0817,
  -60.9977,
  -60.9128,
  -60.8272,
  -60.741,
  -60.6542,
  -60.567,
  -60.4799,
  -60.3928,
  -60.3059,
  -60.2189,
  -60.1318,
  -60.0449,
  -59.9586,
  -59.8733,
  -59.7894,
  -59.7064,
  -59.6245,
  -59.5436,
  -59.4639,
  -59.3855,
  -59.3087,
  -59.2328,
  -59.1579,
  -59.0838,
  -59.011,
  -58.9398,
  -58.8705,
  -58.8035,
  -58.7387,
  -58.6763,
  -58.6163,
  -58.5584,
  -58.5022,
  -58.4476,
  -58.3951,
  -58.3437,
  -58.2957,
  -58.2504,
  -58.2072,
  -58.1653,
  -58.1244,
  -58.0846,
  -58.0464,
  -58.0094,
  -57.974,
  -57.9397,
  -57.9062,
  -57.8734,
  -47.7757,
  -47.6788,
  -47.6096,
  -47.5704,
  -47.5605,
  -47.5768,
  -47.615,
  -47.6704,
  -47.7388,
  -47.821,
  -47.9165,
  -48.028,
  -48.1586,
  -48.3127,
  -48.4942,
  -48.7065,
  -48.9507,
  -49.2243,
  -49.5236,
  -49.8406,
  -50.167,
  -50.4944,
  -50.8158,
  -51.1266,
  -51.4269,
  -51.7161,
  -51.9955,
  -52.2669,
  -52.5312,
  -52.7888,
  -53.0388,
  -53.2804,
  -53.5122,
  -53.7331,
  -53.9422,
  -54.1393,
  -54.3248,
  -54.4996,
  -54.6647,
  -54.8206,
  -54.9714,
  -55.1174,
  -55.2602,
  -55.4004,
  -55.5388,
  -55.6752,
  -55.8093,
  -55.9405,
  -56.0683,
  -56.1915,
  -56.3099,
  -56.4231,
  -56.5314,
  -56.6343,
  -56.7323,
  -56.8246,
  -56.9143,
  -57.0012,
  -57.0864,
  -57.1702,
  -57.2528,
  -57.334,
  -57.4135,
  -57.4914,
  -57.5674,
  -57.6413,
  -57.713,
  -57.7827,
  -57.8509,
  -57.9178,
  -57.9836,
  -58.0489,
  -58.1128,
  -58.1775,
  -58.2423,
  -58.3072,
  -58.3727,
  -58.4392,
  -58.5071,
  -58.5771,
  -58.6495,
  -58.7236,
  -58.7988,
  -58.8745,
  -58.9501,
  -59.0252,
  -59.0995,
  -59.173,
  -59.2458,
  -59.3186,
  -59.3908,
  -59.4653,
  -59.5409,
  -59.6179,
  -59.6954,
  -59.773,
  -59.8504,
  -59.9267,
  -60.0018,
  -60.0753,
  -60.1472,
  -60.2175,
  -60.286,
  -60.3528,
  -60.4178,
  -60.4813,
  -60.544,
  -60.6061,
  -60.6688,
  -60.732,
  -60.7981,
  -60.8665,
  -60.9365,
  -61.0073,
  -61.0783,
  -61.1486,
  -61.2172,
  -61.2831,
  -61.3463,
  -61.4073,
  -61.4669,
  -61.5266,
  -61.5876,
  -61.6512,
  -61.7175,
  -61.7867,
  -61.8577,
  -61.9295,
  -62.0007,
  -62.0705,
  -62.1372,
  -62.202,
  -62.2632,
  -62.3208,
  -62.3754,
  -62.4275,
  -62.4782,
  -62.5288,
  -62.5799,
  -62.6324,
  -62.6863,
  -62.7416,
  -62.7977,
  -62.8538,
  -62.9092,
  -62.9636,
  -63.0168,
  -63.0694,
  -63.1213,
  -63.1725,
  -63.2225,
  -63.271,
  -63.3166,
  -63.3617,
  -63.4052,
  -63.4479,
  -63.4895,
  -63.5302,
  -63.5699,
  -63.6087,
  -63.6462,
  -63.6823,
  -63.7164,
  -63.748,
  -63.7769,
  -63.8029,
  -63.8258,
  -63.8455,
  -63.8619,
  -63.8758,
  -63.8882,
  -63.8992,
  -63.9103,
  -63.9228,
  -63.9366,
  -63.9521,
  -63.9683,
  -63.9883,
  -64.0097,
  -64.0323,
  -64.0554,
  -64.0785,
  -64.1007,
  -64.1212,
  -64.1389,
  -64.1535,
  -64.1647,
  -64.1722,
  -64.1761,
  -64.1762,
  -64.1732,
  -64.167,
  -64.1578,
  -64.1462,
  -64.1326,
  -64.1168,
  -64.0989,
  -64.0792,
  -64.058,
  -64.0353,
  -64.0112,
  -63.9857,
  -63.9589,
  -63.9299,
  -63.9008,
  -63.8706,
  -63.8394,
  -63.8074,
  -63.775,
  -63.7423,
  -63.7093,
  -63.6761,
  -63.6424,
  -63.608,
  -63.5723,
  -63.5352,
  -63.4967,
  -63.4569,
  -63.4159,
  -63.3738,
  -63.3303,
  -63.2853,
  -63.2389,
  -63.1913,
  -63.1429,
  -63.0938,
  -63.0441,
  -62.9933,
  -62.9416,
  -62.8891,
  -62.8361,
  -62.7827,
  -62.7283,
  -62.6725,
  -62.6146,
  -62.5561,
  -62.4955,
  -62.4328,
  -62.3684,
  -62.3026,
  -62.2356,
  -62.1673,
  -62.0975,
  -62.0262,
  -61.9531,
  -61.8783,
  -61.802,
  -61.7247,
  -61.6469,
  -61.5686,
  -61.4893,
  -61.4087,
  -61.3269,
  -61.2438,
  -61.1597,
  -61.0747,
  -60.989,
  -60.9027,
  -60.816,
  -60.7294,
  -60.6428,
  -60.5564,
  -60.4703,
  -60.3843,
  -60.2985,
  -60.2131,
  -60.1285,
  -60.0448,
  -59.962,
  -59.8802,
  -59.7995,
  -59.7203,
  -59.6419,
  -59.5659,
  -59.491,
  -59.4168,
  -59.3435,
  -59.2711,
  -59.2001,
  -59.1308,
  -59.0637,
  -58.9992,
  -58.9373,
  -58.8776,
  -58.8199,
  -58.7635,
  -58.7081,
  -58.6547,
  -58.6035,
  -58.5548,
  -58.5087,
  -58.4646,
  -58.4219,
  -58.3803,
  -58.3397,
  -58.3006,
  -58.2629,
  -58.2266,
  -58.1915,
  -58.1572,
  -58.1237,
  -47.8878,
  -47.8057,
  -47.751,
  -47.7245,
  -47.7265,
  -47.7525,
  -47.7978,
  -47.8582,
  -47.9304,
  -48.0137,
  -48.1091,
  -48.2191,
  -48.3475,
  -48.4979,
  -48.6743,
  -48.879,
  -49.1143,
  -49.3776,
  -49.6641,
  -49.9699,
  -50.2861,
  -50.6051,
  -50.9205,
  -51.2293,
  -51.5293,
  -51.8211,
  -52.1057,
  -52.3847,
  -52.6585,
  -52.9269,
  -53.1885,
  -53.4415,
  -53.6842,
  -53.914,
  -54.1317,
  -54.3363,
  -54.5281,
  -54.7082,
  -54.8777,
  -55.0384,
  -55.1926,
  -55.3421,
  -55.4888,
  -55.6335,
  -55.7771,
  -55.9194,
  -56.06,
  -56.1985,
  -56.3337,
  -56.464,
  -56.5903,
  -56.7114,
  -56.827,
  -56.9363,
  -57.0396,
  -57.1372,
  -57.2304,
  -57.3199,
  -57.4069,
  -57.4921,
  -57.5757,
  -57.6577,
  -57.7378,
  -57.816,
  -57.8922,
  -57.9664,
  -58.0372,
  -58.1067,
  -58.1746,
  -58.2412,
  -58.3072,
  -58.3724,
  -58.4375,
  -58.5025,
  -58.5677,
  -58.6331,
  -58.6992,
  -58.7664,
  -58.8354,
  -58.9064,
  -58.9798,
  -59.0552,
  -59.1318,
  -59.209,
  -59.285,
  -59.3616,
  -59.4375,
  -59.5127,
  -59.5876,
  -59.6623,
  -59.7375,
  -59.8138,
  -59.8914,
  -59.9702,
  -60.0498,
  -60.1295,
  -60.2089,
  -60.2876,
  -60.3651,
  -60.4411,
  -60.5156,
  -60.5883,
  -60.6583,
  -60.7274,
  -60.7942,
  -60.8596,
  -60.9238,
  -60.9874,
  -61.0512,
  -61.1161,
  -61.1827,
  -61.2511,
  -61.3212,
  -61.3919,
  -61.4623,
  -61.5319,
  -61.5996,
  -61.6649,
  -61.7274,
  -61.7879,
  -61.8471,
  -61.9064,
  -61.9663,
  -62.0295,
  -62.0955,
  -62.1644,
  -62.2353,
  -62.3072,
  -62.3789,
  -62.4495,
  -62.518,
  -62.5841,
  -62.647,
  -62.7063,
  -62.7621,
  -62.8152,
  -62.8665,
  -62.9172,
  -62.9681,
  -63.0203,
  -63.0738,
  -63.1286,
  -63.1843,
  -63.2386,
  -63.2929,
  -63.346,
  -63.398,
  -63.4494,
  -63.5004,
  -63.5507,
  -63.6,
  -63.6476,
  -63.6933,
  -63.7368,
  -63.7785,
  -63.8187,
  -63.8575,
  -63.8953,
  -63.9321,
  -63.9681,
  -64.003,
  -64.0365,
  -64.0683,
  -64.0979,
  -64.1247,
  -64.1485,
  -64.1691,
  -64.1851,
  -64.1987,
  -64.2092,
  -64.2174,
  -64.2244,
  -64.2312,
  -64.2389,
  -64.2475,
  -64.258,
  -64.2711,
  -64.2864,
  -64.304,
  -64.3229,
  -64.3417,
  -64.361,
  -64.3795,
  -64.3965,
  -64.4111,
  -64.4229,
  -64.4314,
  -64.4364,
  -64.4377,
  -64.4356,
  -64.4301,
  -64.4216,
  -64.4092,
  -64.3958,
  -64.3804,
  -64.3629,
  -64.3433,
  -64.3221,
  -64.299,
  -64.2744,
  -64.2484,
  -64.221,
  -64.1924,
  -64.1626,
  -64.132,
  -64.1003,
  -64.0681,
  -64.0351,
  -64.0018,
  -63.9683,
  -63.9349,
  -63.9013,
  -63.8674,
  -63.8329,
  -63.7974,
  -63.7605,
  -63.7221,
  -63.6825,
  -63.6418,
  -63.5999,
  -63.5566,
  -63.5119,
  -63.4646,
  -63.417,
  -63.3686,
  -63.3194,
  -63.2694,
  -63.2186,
  -63.167,
  -63.1147,
  -63.0617,
  -63.0082,
  -62.954,
  -62.898,
  -62.8407,
  -62.7814,
  -62.7202,
  -62.6572,
  -62.5923,
  -62.5261,
  -62.4585,
  -62.3899,
  -62.32,
  -62.2485,
  -62.1755,
  -62.1011,
  -62.0257,
  -61.9494,
  -61.8729,
  -61.796,
  -61.7182,
  -61.6393,
  -61.5588,
  -61.4769,
  -61.3938,
  -61.3098,
  -61.2249,
  -61.1384,
  -61.0525,
  -60.9667,
  -60.8808,
  -60.7952,
  -60.7101,
  -60.6252,
  -60.5404,
  -60.4558,
  -60.3719,
  -60.2886,
  -60.206,
  -60.1243,
  -60.0439,
  -59.9651,
  -59.8882,
  -59.8129,
  -59.7388,
  -59.6654,
  -59.5927,
  -59.5207,
  -59.4501,
  -59.3813,
  -59.3147,
  -59.2506,
  -59.1891,
  -59.1298,
  -59.0723,
  -59.0159,
  -58.9605,
  -58.9065,
  -58.8546,
  -58.8053,
  -58.7585,
  -58.7139,
  -58.6706,
  -58.6284,
  -58.5872,
  -58.5473,
  -58.5087,
  -58.4714,
  -58.4352,
  -58.4002,
  -58.3658,
  -48.0115,
  -47.9454,
  -47.9062,
  -47.8942,
  -47.9072,
  -47.9423,
  -47.9941,
  -48.0587,
  -48.1338,
  -48.219,
  -48.3154,
  -48.4254,
  -48.5533,
  -48.7012,
  -48.8744,
  -49.074,
  -49.3014,
  -49.5552,
  -49.8316,
  -50.1255,
  -50.4305,
  -50.7401,
  -51.0484,
  -51.3529,
  -51.6514,
  -51.9441,
  -52.2324,
  -52.5174,
  -52.7983,
  -53.0761,
  -53.3479,
  -53.6111,
  -53.8634,
  -54.1031,
  -54.329,
  -54.5407,
  -54.7387,
  -54.9239,
  -55.0979,
  -55.2625,
  -55.4198,
  -55.5724,
  -55.7224,
  -55.8702,
  -56.0183,
  -56.1659,
  -56.3127,
  -56.458,
  -56.6005,
  -56.7396,
  -56.874,
  -57.003,
  -57.1255,
  -57.2412,
  -57.3498,
  -57.452,
  -57.5484,
  -57.6405,
  -57.7294,
  -57.8158,
  -57.8994,
  -57.9821,
  -58.0628,
  -58.1414,
  -58.2177,
  -58.2916,
  -58.3636,
  -58.4333,
  -58.5011,
  -58.5677,
  -58.6338,
  -58.6995,
  -58.7646,
  -58.83,
  -58.8957,
  -58.9616,
  -59.0284,
  -59.0953,
  -59.1648,
  -59.2364,
  -59.3103,
  -59.3866,
  -59.4641,
  -59.5422,
  -59.6205,
  -59.6983,
  -59.7753,
  -59.852,
  -59.9285,
  -60.0051,
  -60.0823,
  -60.1603,
  -60.2395,
  -60.3201,
  -60.4015,
  -60.4823,
  -60.5638,
  -60.6445,
  -60.7243,
  -60.803,
  -60.8799,
  -60.9549,
  -61.0281,
  -61.0995,
  -61.1684,
  -61.2358,
  -61.3012,
  -61.3664,
  -61.4314,
  -61.4971,
  -61.5641,
  -61.6327,
  -61.7027,
  -61.7734,
  -61.844,
  -61.9123,
  -61.9798,
  -62.0449,
  -62.1076,
  -62.1682,
  -62.2277,
  -62.2872,
  -62.3477,
  -62.4104,
  -62.4757,
  -62.5437,
  -62.6138,
  -62.685,
  -62.7563,
  -62.8267,
  -62.8953,
  -62.9619,
  -63.0255,
  -63.0857,
  -63.1425,
  -63.1962,
  -63.2469,
  -63.2975,
  -63.3478,
  -63.3993,
  -63.4525,
  -63.5071,
  -63.562,
  -63.6163,
  -63.6694,
  -63.7209,
  -63.7715,
  -63.8216,
  -63.8714,
  -63.9209,
  -63.9693,
  -64.0162,
  -64.0608,
  -64.103,
  -64.1427,
  -64.1805,
  -64.2166,
  -64.2515,
  -64.2845,
  -64.3175,
  -64.3495,
  -64.3802,
  -64.4095,
  -64.4368,
  -64.4618,
  -64.4837,
  -64.5021,
  -64.5167,
  -64.5275,
  -64.5351,
  -64.54,
  -64.5434,
  -64.5462,
  -64.5493,
  -64.5532,
  -64.5591,
  -64.5674,
  -64.5787,
  -64.5915,
  -64.606,
  -64.6206,
  -64.6354,
  -64.6494,
  -64.6608,
  -64.6714,
  -64.6796,
  -64.6849,
  -64.6869,
  -64.6854,
  -64.6805,
  -64.6725,
  -64.6617,
  -64.6484,
  -64.6331,
  -64.6163,
  -64.5974,
  -64.5763,
  -64.5533,
  -64.5288,
  -64.5024,
  -64.4743,
  -64.4451,
  -64.4148,
  -64.3835,
  -64.3515,
  -64.3187,
  -64.2854,
  -64.2516,
  -64.2176,
  -64.1834,
  -64.1492,
  -64.114,
  -64.0795,
  -64.0446,
  -64.0088,
  -63.9717,
  -63.9335,
  -63.894,
  -63.8535,
  -63.8118,
  -63.7688,
  -63.7242,
  -63.6782,
  -63.631,
  -63.5828,
  -63.5337,
  -63.4837,
  -63.433,
  -63.3818,
  -63.33,
  -63.2777,
  -63.2242,
  -63.17,
  -63.1141,
  -63.0563,
  -62.9967,
  -62.9351,
  -62.8715,
  -62.8063,
  -62.7396,
  -62.6716,
  -62.6025,
  -62.5319,
  -62.459,
  -62.3858,
  -62.3116,
  -62.2365,
  -62.161,
  -62.0853,
  -62.0095,
  -61.9331,
  -61.8557,
  -61.7767,
  -61.6962,
  -61.6143,
  -61.5313,
  -61.4476,
  -61.3632,
  -61.2784,
  -61.1934,
  -61.1082,
  -61.0234,
  -60.9392,
  -60.8553,
  -60.7716,
  -60.6881,
  -60.6048,
  -60.522,
  -60.4394,
  -60.358,
  -60.2775,
  -60.1991,
  -60.1226,
  -60.0479,
  -59.9743,
  -59.9012,
  -59.8289,
  -59.7574,
  -59.6873,
  -59.6191,
  -59.5531,
  -59.4897,
  -59.4287,
  -59.3698,
  -59.3115,
  -59.2553,
  -59.2001,
  -59.146,
  -59.0941,
  -59.0445,
  -58.9973,
  -58.9523,
  -58.9084,
  -58.8662,
  -58.8249,
  -58.7846,
  -58.7453,
  -58.7068,
  -58.6697,
  -58.6335,
  -58.5981,
  -48.1504,
  -48.1007,
  -48.0765,
  -48.0774,
  -48.101,
  -48.1437,
  -48.2012,
  -48.2688,
  -48.3467,
  -48.4341,
  -48.5324,
  -48.6446,
  -48.7738,
  -48.9231,
  -49.0951,
  -49.2915,
  -49.5134,
  -49.7593,
  -50.026,
  -50.3092,
  -50.6034,
  -50.9034,
  -51.2032,
  -51.5022,
  -51.7981,
  -52.091,
  -52.3817,
  -52.6708,
  -52.9583,
  -53.2428,
  -53.522,
  -53.793,
  -54.0531,
  -54.3004,
  -54.5335,
  -54.752,
  -54.956,
  -55.1466,
  -55.3242,
  -55.4927,
  -55.6535,
  -55.8091,
  -55.962,
  -56.1139,
  -56.2658,
  -56.4179,
  -56.5698,
  -56.7211,
  -56.8705,
  -57.0169,
  -57.1589,
  -57.2951,
  -57.4244,
  -57.5461,
  -57.6591,
  -57.7656,
  -57.8656,
  -57.9604,
  -58.0512,
  -58.1389,
  -58.2242,
  -58.3074,
  -58.3884,
  -58.4674,
  -58.5437,
  -58.6177,
  -58.6897,
  -58.7598,
  -58.8282,
  -58.8954,
  -58.9618,
  -59.0269,
  -59.0927,
  -59.1585,
  -59.2245,
  -59.291,
  -59.3581,
  -59.4264,
  -59.4962,
  -59.5682,
  -59.6423,
  -59.7187,
  -59.7967,
  -59.8755,
  -59.9544,
  -60.0328,
  -60.1109,
  -60.1885,
  -60.2663,
  -60.3435,
  -60.4223,
  -60.502,
  -60.5829,
  -60.665,
  -60.7482,
  -60.8316,
  -60.915,
  -60.9978,
  -61.0795,
  -61.1602,
  -61.2394,
  -61.3168,
  -61.3922,
  -61.4655,
  -61.5366,
  -61.6056,
  -61.673,
  -61.7394,
  -61.8047,
  -61.8714,
  -61.9391,
  -62.008,
  -62.0782,
  -62.1489,
  -62.2195,
  -62.2893,
  -62.3573,
  -62.4231,
  -62.4866,
  -62.5481,
  -62.6083,
  -62.6682,
  -62.7285,
  -62.7903,
  -62.8545,
  -62.9212,
  -62.9899,
  -63.0599,
  -63.129,
  -63.1985,
  -63.2665,
  -63.3326,
  -63.3961,
  -63.4565,
  -63.5136,
  -63.5677,
  -63.6195,
  -63.6701,
  -63.7202,
  -63.7712,
  -63.8235,
  -63.877,
  -63.9308,
  -63.9839,
  -64.0355,
  -64.0855,
  -64.1347,
  -64.1834,
  -64.2323,
  -64.2808,
  -64.3274,
  -64.3733,
  -64.417,
  -64.4578,
  -64.4958,
  -64.5314,
  -64.565,
  -64.5972,
  -64.6282,
  -64.6581,
  -64.6871,
  -64.715,
  -64.7415,
  -64.7663,
  -64.7889,
  -64.8086,
  -64.8246,
  -64.8369,
  -64.8452,
  -64.8501,
  -64.8521,
  -64.8525,
  -64.8519,
  -64.8509,
  -64.8498,
  -64.8513,
  -64.8552,
  -64.8616,
  -64.87,
  -64.8795,
  -64.8894,
  -64.8992,
  -64.9082,
  -64.9161,
  -64.9223,
  -64.9265,
  -64.9281,
  -64.9265,
  -64.9216,
  -64.9136,
  -64.9026,
  -64.8892,
  -64.8738,
  -64.8568,
  -64.8381,
  -64.8178,
  -64.7955,
  -64.7712,
  -64.745,
  -64.7169,
  -64.6864,
  -64.6558,
  -64.6241,
  -64.5916,
  -64.5584,
  -64.5246,
  -64.4902,
  -64.4556,
  -64.4208,
  -64.3858,
  -64.3507,
  -64.3155,
  -64.2801,
  -64.2443,
  -64.208,
  -64.1708,
  -64.1326,
  -64.0933,
  -64.053,
  -64.0116,
  -63.9689,
  -63.9247,
  -63.879,
  -63.8321,
  -63.7842,
  -63.7353,
  -63.6855,
  -63.6351,
  -63.5841,
  -63.5328,
  -63.4807,
  -63.4267,
  -63.3722,
  -63.3161,
  -63.2582,
  -63.1985,
  -63.1371,
  -63.0739,
  -63.0087,
  -62.9419,
  -62.8737,
  -62.8039,
  -62.7329,
  -62.6605,
  -62.587,
  -62.5124,
  -62.4373,
  -62.3618,
  -62.2865,
  -62.2113,
  -62.1359,
  -62.0597,
  -61.9821,
  -61.9029,
  -61.8222,
  -61.7405,
  -61.6579,
  -61.5746,
  -61.491,
  -61.4069,
  -61.3229,
  -61.2393,
  -61.1561,
  -61.0735,
  -60.991,
  -60.9085,
  -60.8258,
  -60.7433,
  -60.6599,
  -60.5782,
  -60.4978,
  -60.4194,
  -60.3432,
  -60.2687,
  -60.1954,
  -60.1228,
  -60.0509,
  -59.9798,
  -59.9104,
  -59.8427,
  -59.7772,
  -59.714,
  -59.6532,
  -59.5943,
  -59.5371,
  -59.4809,
  -59.4258,
  -59.372,
  -59.3203,
  -59.2708,
  -59.2237,
  -59.1785,
  -59.1348,
  -59.0926,
  -59.0512,
  -59.0108,
  -58.9712,
  -58.9323,
  -58.8944,
  -58.8574,
  -58.8214,
  -48.3071,
  -48.2736,
  -48.2631,
  -48.2759,
  -48.3085,
  -48.3571,
  -48.4189,
  -48.4906,
  -48.5708,
  -48.6606,
  -48.7617,
  -48.8767,
  -49.0088,
  -49.1604,
  -49.3337,
  -49.5294,
  -49.7483,
  -49.9877,
  -50.2469,
  -50.5208,
  -50.8053,
  -51.0961,
  -51.3896,
  -51.6828,
  -51.9755,
  -52.2669,
  -52.5582,
  -52.8492,
  -53.1397,
  -53.4282,
  -53.7121,
  -53.9884,
  -54.2532,
  -54.5065,
  -54.7459,
  -54.9703,
  -55.1799,
  -55.3759,
  -55.5593,
  -55.7322,
  -55.8964,
  -56.0551,
  -56.2107,
  -56.3653,
  -56.5201,
  -56.6757,
  -56.832,
  -56.9882,
  -57.1425,
  -57.2951,
  -57.4436,
  -57.5863,
  -57.7216,
  -57.8486,
  -57.9671,
  -58.0777,
  -58.1812,
  -58.2786,
  -58.3715,
  -58.4607,
  -58.547,
  -58.6307,
  -58.7121,
  -58.7913,
  -58.8679,
  -58.9413,
  -59.0134,
  -59.0841,
  -59.1532,
  -59.2215,
  -59.2888,
  -59.3556,
  -59.4221,
  -59.4883,
  -59.5546,
  -59.6214,
  -59.6888,
  -59.7574,
  -59.8273,
  -59.8992,
  -59.9733,
  -60.0495,
  -60.1264,
  -60.2054,
  -60.2847,
  -60.3636,
  -60.442,
  -60.5203,
  -60.5991,
  -60.6785,
  -60.7588,
  -60.8401,
  -60.9225,
  -61.0061,
  -61.0905,
  -61.1755,
  -61.2603,
  -61.3446,
  -61.4281,
  -61.5107,
  -61.5918,
  -61.6701,
  -61.7475,
  -61.823,
  -61.8962,
  -61.9674,
  -62.0366,
  -62.1048,
  -62.1725,
  -62.2402,
  -62.3085,
  -62.3775,
  -62.4477,
  -62.5185,
  -62.5893,
  -62.6595,
  -62.7285,
  -62.7956,
  -62.8606,
  -62.9237,
  -62.9839,
  -63.0442,
  -63.1042,
  -63.1651,
  -63.2278,
  -63.2927,
  -63.3596,
  -63.4278,
  -63.4965,
  -63.5644,
  -63.6314,
  -63.6965,
  -63.7591,
  -63.8189,
  -63.8758,
  -63.93,
  -63.9819,
  -64.0323,
  -64.0822,
  -64.1325,
  -64.1839,
  -64.2361,
  -64.2876,
  -64.3392,
  -64.3891,
  -64.4377,
  -64.4855,
  -64.5331,
  -64.5808,
  -64.6283,
  -64.6751,
  -64.7202,
  -64.7628,
  -64.8024,
  -64.8388,
  -64.8725,
  -64.9038,
  -64.9334,
  -64.9616,
  -64.9885,
  -65.0144,
  -65.0392,
  -65.0627,
  -65.0849,
  -65.1049,
  -65.1208,
  -65.1342,
  -65.1439,
  -65.1497,
  -65.1518,
  -65.1514,
  -65.1491,
  -65.1457,
  -65.1418,
  -65.138,
  -65.1356,
  -65.1353,
  -65.1371,
  -65.1407,
  -65.1452,
  -65.15,
  -65.1545,
  -65.1584,
  -65.1613,
  -65.1629,
  -65.163,
  -65.1603,
  -65.1549,
  -65.1463,
  -65.1347,
  -65.1195,
  -65.1033,
  -65.0855,
  -65.0664,
  -65.0459,
  -65.0239,
  -65.0001,
  -64.9743,
  -64.9466,
  -64.917,
  -64.8861,
  -64.8542,
  -64.8214,
  -64.7878,
  -64.7534,
  -64.7187,
  -64.6836,
  -64.6482,
  -64.6127,
  -64.5769,
  -64.5408,
  -64.5044,
  -64.4679,
  -64.4312,
  -64.3941,
  -64.3566,
  -64.3184,
  -64.2792,
  -64.2389,
  -64.1965,
  -64.1541,
  -64.1099,
  -64.065,
  -64.0186,
  -63.9713,
  -63.9228,
  -63.8734,
  -63.8231,
  -63.7725,
  -63.7214,
  -63.6695,
  -63.6164,
  -63.5616,
  -63.5054,
  -63.4477,
  -63.3885,
  -63.3277,
  -63.2653,
  -63.2009,
  -63.1346,
  -63.0665,
  -62.9964,
  -62.9248,
  -62.8517,
  -62.7774,
  -62.7024,
  -62.6267,
  -62.5508,
  -62.4754,
  -62.4002,
  -62.3253,
  -62.2498,
  -62.1734,
  -62.0955,
  -62.0152,
  -61.9348,
  -61.8533,
  -61.7712,
  -61.6885,
  -61.6056,
  -61.5227,
  -61.4404,
  -61.3586,
  -61.2773,
  -61.1957,
  -61.1141,
  -61.0321,
  -60.9498,
  -60.8675,
  -60.7856,
  -60.7052,
  -60.6268,
  -60.5506,
  -60.4762,
  -60.4029,
  -60.3304,
  -60.2588,
  -60.1882,
  -60.1192,
  -60.0521,
  -59.9872,
  -59.9242,
  -59.8629,
  -59.8035,
  -59.7457,
  -59.6895,
  -59.6348,
  -59.5817,
  -59.5305,
  -59.4816,
  -59.4347,
  -59.3899,
  -59.3467,
  -59.3048,
  -59.2639,
  -59.2239,
  -59.1847,
  -59.1458,
  -59.1077,
  -59.0693,
  -59.0332,
  -48.4826,
  -48.4648,
  -48.4681,
  -48.491,
  -48.5309,
  -48.5844,
  -48.6489,
  -48.7229,
  -48.8053,
  -48.8977,
  -49.0021,
  -49.12,
  -49.2561,
  -49.4119,
  -49.5881,
  -49.7851,
  -50.0033,
  -50.2406,
  -50.4945,
  -50.7616,
  -51.0383,
  -51.3215,
  -51.6082,
  -51.8962,
  -52.1847,
  -52.4737,
  -52.7625,
  -53.053,
  -53.3437,
  -53.633,
  -53.9184,
  -54.1973,
  -54.4667,
  -54.7243,
  -54.9689,
  -55.1989,
  -55.4144,
  -55.6159,
  -55.8045,
  -55.9819,
  -56.1497,
  -56.3112,
  -56.4681,
  -56.6247,
  -56.7817,
  -56.9396,
  -57.0989,
  -57.2589,
  -57.4185,
  -57.5761,
  -57.7296,
  -57.8775,
  -58.0179,
  -58.1493,
  -58.2719,
  -58.386,
  -58.4925,
  -58.5926,
  -58.6874,
  -58.777,
  -58.8643,
  -58.9488,
  -59.0307,
  -59.1102,
  -59.1873,
  -59.2621,
  -59.335,
  -59.4063,
  -59.4764,
  -59.5456,
  -59.6141,
  -59.682,
  -59.7493,
  -59.8163,
  -59.883,
  -59.9503,
  -60.017,
  -60.0858,
  -60.1559,
  -60.2274,
  -60.3011,
  -60.377,
  -60.4545,
  -60.5334,
  -60.6126,
  -60.6914,
  -60.7699,
  -60.8487,
  -60.9279,
  -61.008,
  -61.0893,
  -61.1718,
  -61.2554,
  -61.3401,
  -61.4245,
  -61.5105,
  -61.5969,
  -61.6828,
  -61.7678,
  -61.8518,
  -61.9344,
  -62.0154,
  -62.0946,
  -62.1721,
  -62.2474,
  -62.3208,
  -62.3922,
  -62.4625,
  -62.5318,
  -62.6008,
  -62.6698,
  -62.7392,
  -62.8093,
  -62.879,
  -62.9501,
  -63.0209,
  -63.0908,
  -63.1592,
  -63.2258,
  -63.2902,
  -63.3527,
  -63.4135,
  -63.4733,
  -63.5333,
  -63.5944,
  -63.6574,
  -63.722,
  -63.7881,
  -63.8547,
  -63.921,
  -63.9862,
  -64.0495,
  -64.1108,
  -64.1697,
  -64.2251,
  -64.2792,
  -64.3312,
  -64.3816,
  -64.4314,
  -64.4813,
  -64.5314,
  -64.5824,
  -64.6328,
  -64.6828,
  -64.7312,
  -64.7782,
  -64.8247,
  -64.871,
  -64.9176,
  -64.9642,
  -65.01,
  -65.0541,
  -65.0956,
  -65.1339,
  -65.169,
  -65.2011,
  -65.2296,
  -65.257,
  -65.2826,
  -65.3069,
  -65.3297,
  -65.3514,
  -65.3719,
  -65.3911,
  -65.408,
  -65.4221,
  -65.4328,
  -65.4396,
  -65.4427,
  -65.4427,
  -65.44,
  -65.4352,
  -65.4293,
  -65.4225,
  -65.4156,
  -65.4094,
  -65.4048,
  -65.4021,
  -65.4007,
  -65.4005,
  -65.4003,
  -65.3989,
  -65.3978,
  -65.3958,
  -65.3928,
  -65.388,
  -65.3812,
  -65.3714,
  -65.3586,
  -65.3432,
  -65.3256,
  -65.3061,
  -65.2854,
  -65.2637,
  -65.241,
  -65.2169,
  -65.1913,
  -65.164,
  -65.1348,
  -65.104,
  -65.072,
  -65.039,
  -65.0052,
  -64.9707,
  -64.9356,
  -64.9001,
  -64.8644,
  -64.8283,
  -64.7911,
  -64.7544,
  -64.7173,
  -64.6799,
  -64.6424,
  -64.6048,
  -64.5671,
  -64.5293,
  -64.4909,
  -64.4516,
  -64.4113,
  -64.3698,
  -64.3272,
  -64.2836,
  -64.2389,
  -64.1933,
  -64.1464,
  -64.0982,
  -64.0487,
  -63.9986,
  -63.948,
  -63.8968,
  -63.8453,
  -63.7923,
  -63.7378,
  -63.6819,
  -63.6248,
  -63.5666,
  -63.5068,
  -63.4454,
  -63.3818,
  -63.3159,
  -63.2469,
  -63.1766,
  -63.1044,
  -63.0307,
  -62.9557,
  -62.8798,
  -62.8034,
  -62.727,
  -62.6511,
  -62.5758,
  -62.501,
  -62.4262,
  -62.3505,
  -62.2736,
  -62.1953,
  -62.1157,
  -62.0351,
  -61.9537,
  -61.8719,
  -61.79,
  -61.7085,
  -61.6276,
  -61.5472,
  -61.4671,
  -61.3869,
  -61.3062,
  -61.2246,
  -61.1425,
  -61.0601,
  -60.9782,
  -60.8977,
  -60.8192,
  -60.7425,
  -60.6678,
  -60.5944,
  -60.522,
  -60.4506,
  -60.3804,
  -60.3121,
  -60.2456,
  -60.1808,
  -60.1167,
  -60.0548,
  -59.9946,
  -59.9363,
  -59.8796,
  -59.8249,
  -59.7722,
  -59.7217,
  -59.6734,
  -59.6273,
  -59.5833,
  -59.5411,
  -59.5001,
  -59.4602,
  -59.4211,
  -59.3823,
  -59.3438,
  -59.3061,
  -59.2692,
  -59.2334,
  -48.6791,
  -48.6757,
  -48.6902,
  -48.7214,
  -48.7667,
  -48.8233,
  -48.8888,
  -48.9641,
  -49.0484,
  -49.1434,
  -49.2513,
  -49.3748,
  -49.5161,
  -49.6769,
  -49.8576,
  -50.0579,
  -50.2773,
  -50.5139,
  -50.7648,
  -51.0275,
  -51.2987,
  -51.5747,
  -51.8557,
  -52.1386,
  -52.4227,
  -52.7081,
  -52.9949,
  -53.2828,
  -53.571,
  -53.8584,
  -54.1427,
  -54.4218,
  -54.693,
  -54.9536,
  -55.2022,
  -55.4376,
  -55.6579,
  -55.865,
  -56.0588,
  -56.2408,
  -56.4126,
  -56.5768,
  -56.7366,
  -56.8947,
  -57.0528,
  -57.2122,
  -57.3733,
  -57.5356,
  -57.698,
  -57.8589,
  -58.0162,
  -58.1676,
  -58.3115,
  -58.4454,
  -58.571,
  -58.6879,
  -58.7969,
  -58.8992,
  -58.9961,
  -59.0882,
  -59.1765,
  -59.2617,
  -59.3441,
  -59.4242,
  -59.5019,
  -59.5775,
  -59.6514,
  -59.7235,
  -59.7947,
  -59.8649,
  -59.9335,
  -60.0026,
  -60.071,
  -60.1389,
  -60.2066,
  -60.2743,
  -60.3424,
  -60.4114,
  -60.4816,
  -60.553,
  -60.6263,
  -60.7016,
  -60.7787,
  -60.8569,
  -60.9357,
  -61.0145,
  -61.0929,
  -61.1705,
  -61.2497,
  -61.33,
  -61.4118,
  -61.4949,
  -61.5792,
  -61.6647,
  -61.7511,
  -61.8384,
  -61.9257,
  -62.013,
  -62.0994,
  -62.1847,
  -62.2685,
  -62.3508,
  -62.4316,
  -62.5109,
  -62.5885,
  -62.6641,
  -62.737,
  -62.8094,
  -62.8806,
  -62.9511,
  -63.021,
  -63.091,
  -63.1613,
  -63.232,
  -63.3031,
  -63.3741,
  -63.4446,
  -63.514,
  -63.5817,
  -63.6474,
  -63.7108,
  -63.7721,
  -63.8318,
  -63.891,
  -63.9507,
  -64.0116,
  -64.073,
  -64.1365,
  -64.2005,
  -64.2644,
  -64.3276,
  -64.3891,
  -64.4487,
  -64.5065,
  -64.5622,
  -64.6161,
  -64.6683,
  -64.7188,
  -64.7684,
  -64.8175,
  -64.867,
  -64.9162,
  -64.9651,
  -65.013,
  -65.0597,
  -65.1055,
  -65.1507,
  -65.1957,
  -65.2402,
  -65.2856,
  -65.3302,
  -65.3731,
  -65.4133,
  -65.4504,
  -65.4844,
  -65.5151,
  -65.5433,
  -65.5689,
  -65.5925,
  -65.6143,
  -65.6344,
  -65.6532,
  -65.6706,
  -65.6866,
  -65.7006,
  -65.7116,
  -65.7192,
  -65.7231,
  -65.7237,
  -65.7209,
  -65.7151,
  -65.7082,
  -65.6995,
  -65.6903,
  -65.6803,
  -65.6704,
  -65.6618,
  -65.6546,
  -65.6485,
  -65.6435,
  -65.6387,
  -65.6336,
  -65.6278,
  -65.6211,
  -65.6134,
  -65.6039,
  -65.5922,
  -65.5777,
  -65.5604,
  -65.5409,
  -65.5194,
  -65.4964,
  -65.4725,
  -65.4478,
  -65.4223,
  -65.3958,
  -65.3681,
  -65.3379,
  -65.3072,
  -65.2753,
  -65.2422,
  -65.2084,
  -65.1738,
  -65.1386,
  -65.1029,
  -65.0669,
  -65.0307,
  -64.9942,
  -64.9574,
  -64.9203,
  -64.8825,
  -64.8443,
  -64.806,
  -64.7677,
  -64.7296,
  -64.6912,
  -64.6526,
  -64.613,
  -64.5724,
  -64.5309,
  -64.4881,
  -64.4446,
  -64.4002,
  -64.3547,
  -64.3082,
  -64.2602,
  -64.2098,
  -64.1599,
  -64.1093,
  -64.0585,
  -64.0071,
  -63.9545,
  -63.9006,
  -63.8452,
  -63.789,
  -63.7315,
  -63.6727,
  -63.612,
  -63.549,
  -63.4834,
  -63.4152,
  -63.3449,
  -63.2723,
  -63.1981,
  -63.1225,
  -63.0459,
  -62.9688,
  -62.8918,
  -62.8153,
  -62.7398,
  -62.6651,
  -62.5906,
  -62.5157,
  -62.4396,
  -62.3621,
  -62.2832,
  -62.203,
  -62.122,
  -62.0407,
  -61.9597,
  -61.879,
  -61.7992,
  -61.72,
  -61.6411,
  -61.5618,
  -61.4809,
  -61.3999,
  -61.3178,
  -61.2354,
  -61.1535,
  -61.0727,
  -60.9937,
  -60.9166,
  -60.8413,
  -60.7674,
  -60.6949,
  -60.6236,
  -60.554,
  -60.4862,
  -60.4202,
  -60.3554,
  -60.292,
  -60.2297,
  -60.1686,
  -60.1095,
  -60.0526,
  -59.9979,
  -59.9457,
  -59.896,
  -59.8486,
  -59.8034,
  -59.7605,
  -59.7193,
  -59.6797,
  -59.6411,
  -59.603,
  -59.5654,
  -59.5278,
  -59.4909,
  -59.4547,
  -59.4196,
  -48.8937,
  -48.9021,
  -48.9263,
  -48.9636,
  -49.0125,
  -49.0711,
  -49.1385,
  -49.2148,
  -49.3006,
  -49.3983,
  -49.5103,
  -49.6389,
  -49.7865,
  -49.9533,
  -50.1395,
  -50.3441,
  -50.5648,
  -50.8021,
  -51.0518,
  -51.3117,
  -51.5791,
  -51.8516,
  -52.1278,
  -52.406,
  -52.6855,
  -52.9665,
  -53.249,
  -53.5329,
  -53.8168,
  -54.1005,
  -54.3821,
  -54.6587,
  -54.93,
  -55.1928,
  -55.4449,
  -55.685,
  -55.9118,
  -56.1247,
  -56.3238,
  -56.5104,
  -56.6859,
  -56.853,
  -57.0145,
  -57.1735,
  -57.3322,
  -57.4921,
  -57.6539,
  -57.8163,
  -57.9801,
  -58.1427,
  -58.3018,
  -58.4551,
  -58.6009,
  -58.7379,
  -58.8654,
  -58.9843,
  -59.0953,
  -59.1995,
  -59.2978,
  -59.3913,
  -59.4808,
  -59.5669,
  -59.65,
  -59.7296,
  -59.808,
  -59.8843,
  -59.9591,
  -60.0326,
  -60.1048,
  -60.1762,
  -60.247,
  -60.3173,
  -60.387,
  -60.456,
  -60.5245,
  -60.5929,
  -60.6617,
  -60.731,
  -60.8012,
  -60.8727,
  -60.9457,
  -61.0195,
  -61.096,
  -61.1736,
  -61.2519,
  -61.3302,
  -61.4084,
  -61.4866,
  -61.5657,
  -61.6459,
  -61.7274,
  -61.8105,
  -61.8952,
  -61.9812,
  -62.0684,
  -62.1563,
  -62.2448,
  -62.3331,
  -62.4207,
  -62.5062,
  -62.5913,
  -62.6751,
  -62.7573,
  -62.8384,
  -62.918,
  -62.9959,
  -63.0723,
  -63.147,
  -63.22,
  -63.2923,
  -63.3635,
  -63.4342,
  -63.5048,
  -63.5754,
  -63.6461,
  -63.7169,
  -63.7874,
  -63.8572,
  -63.9256,
  -63.9908,
  -64.0549,
  -64.1165,
  -64.1761,
  -64.2347,
  -64.2932,
  -64.3523,
  -64.4123,
  -64.473,
  -64.5342,
  -64.5955,
  -64.6561,
  -64.7157,
  -64.7738,
  -64.8305,
  -64.8855,
  -64.939,
  -64.991,
  -65.0416,
  -65.091,
  -65.1393,
  -65.1866,
  -65.2342,
  -65.2811,
  -65.3274,
  -65.3728,
  -65.4174,
  -65.4615,
  -65.5055,
  -65.5496,
  -65.5935,
  -65.6366,
  -65.6781,
  -65.7173,
  -65.7534,
  -65.7863,
  -65.8162,
  -65.8433,
  -65.8677,
  -65.8896,
  -65.9092,
  -65.927,
  -65.943,
  -65.9567,
  -65.9696,
  -65.9804,
  -65.9882,
  -65.9929,
  -65.994,
  -65.9917,
  -65.9863,
  -65.9786,
  -65.9692,
  -65.9583,
  -65.9456,
  -65.9327,
  -65.9194,
  -65.9068,
  -65.8954,
  -65.8851,
  -65.8758,
  -65.8667,
  -65.8573,
  -65.8473,
  -65.8361,
  -65.8236,
  -65.809,
  -65.7922,
  -65.7718,
  -65.75,
  -65.7259,
  -65.7002,
  -65.6734,
  -65.6461,
  -65.6181,
  -65.5895,
  -65.5604,
  -65.5303,
  -65.4992,
  -65.4667,
  -65.4333,
  -65.3989,
  -65.364,
  -65.3286,
  -65.2927,
  -65.2565,
  -65.2202,
  -65.184,
  -65.1475,
  -65.1106,
  -65.0732,
  -65.0353,
  -64.9969,
  -64.9583,
  -64.9194,
  -64.8808,
  -64.841,
  -64.8019,
  -64.762,
  -64.7213,
  -64.6795,
  -64.6365,
  -64.5928,
  -64.5482,
  -64.5027,
  -64.456,
  -64.408,
  -64.359,
  -64.3094,
  -64.2592,
  -64.2089,
  -64.1577,
  -64.1053,
  -64.0519,
  -63.9973,
  -63.9415,
  -63.8847,
  -63.8264,
  -63.7662,
  -63.7034,
  -63.638,
  -63.5698,
  -63.4993,
  -63.4267,
  -63.3521,
  -63.276,
  -63.1988,
  -63.1211,
  -63.0434,
  -62.9666,
  -62.8898,
  -62.8151,
  -62.7409,
  -62.6665,
  -62.591,
  -62.5141,
  -62.4355,
  -62.3556,
  -62.2749,
  -62.1938,
  -62.1131,
  -62.0332,
  -61.9543,
  -61.8762,
  -61.798,
  -61.7193,
  -61.6397,
  -61.5589,
  -61.477,
  -61.3945,
  -61.3123,
  -61.2311,
  -61.1515,
  -61.0736,
  -60.9975,
  -60.923,
  -60.8502,
  -60.7789,
  -60.7095,
  -60.6421,
  -60.5764,
  -60.5118,
  -60.4481,
  -60.3853,
  -60.324,
  -60.2646,
  -60.2076,
  -60.1533,
  -60.1015,
  -60.0526,
  -60.0061,
  -59.9623,
  -59.9207,
  -59.881,
  -59.8426,
  -59.8043,
  -59.7674,
  -59.731,
  -59.6949,
  -59.6592,
  -59.6238,
  -59.5902,
  -49.1211,
  -49.1417,
  -49.174,
  -49.2164,
  -49.2676,
  -49.3271,
  -49.3949,
  -49.4717,
  -49.5593,
  -49.6599,
  -49.7753,
  -49.9096,
  -50.0632,
  -50.2363,
  -50.4287,
  -50.6383,
  -50.8632,
  -51.1019,
  -51.3515,
  -51.6097,
  -51.8745,
  -52.1434,
  -52.4152,
  -52.6891,
  -52.9642,
  -53.2395,
  -53.5172,
  -53.7959,
  -54.0751,
  -54.3541,
  -54.6321,
  -54.9074,
  -55.178,
  -55.4421,
  -55.6972,
  -55.9415,
  -56.1736,
  -56.3919,
  -56.5963,
  -56.7874,
  -56.9666,
  -57.1354,
  -57.2986,
  -57.4583,
  -57.6172,
  -57.777,
  -57.9386,
  -58.1017,
  -58.2654,
  -58.4279,
  -58.587,
  -58.7408,
  -58.8871,
  -59.0246,
  -59.1533,
  -59.2731,
  -59.3853,
  -59.49,
  -59.5898,
  -59.6844,
  -59.7747,
  -59.8615,
  -59.9454,
  -60.0267,
  -60.1057,
  -60.1828,
  -60.2585,
  -60.3332,
  -60.4069,
  -60.4795,
  -60.5514,
  -60.6227,
  -60.6935,
  -60.7638,
  -60.8322,
  -60.9015,
  -60.9709,
  -61.0406,
  -61.1112,
  -61.1827,
  -61.2558,
  -61.3303,
  -61.4064,
  -61.4835,
  -61.5611,
  -61.6389,
  -61.7168,
  -61.7948,
  -61.8732,
  -61.9527,
  -62.0338,
  -62.1166,
  -62.2012,
  -62.2865,
  -62.3742,
  -62.4629,
  -62.5523,
  -62.6416,
  -62.7303,
  -62.818,
  -62.9042,
  -62.989,
  -63.0727,
  -63.1552,
  -63.2369,
  -63.3173,
  -63.3959,
  -63.4727,
  -63.5481,
  -63.6221,
  -63.6947,
  -63.7663,
  -63.8362,
  -63.9065,
  -63.9767,
  -64.0468,
  -64.1168,
  -64.1862,
  -64.2545,
  -64.321,
  -64.3852,
  -64.4471,
  -64.5069,
  -64.565,
  -64.6225,
  -64.68,
  -64.7374,
  -64.7953,
  -64.8533,
  -64.9116,
  -64.9698,
  -65.0273,
  -65.0831,
  -65.1386,
  -65.1929,
  -65.246,
  -65.2976,
  -65.3478,
  -65.3968,
  -65.4445,
  -65.4913,
  -65.5373,
  -65.5827,
  -65.6274,
  -65.6716,
  -65.7152,
  -65.7583,
  -65.8014,
  -65.844,
  -65.8861,
  -65.9276,
  -65.9675,
  -66.0056,
  -66.0399,
  -66.0723,
  -66.1017,
  -66.1281,
  -66.1517,
  -66.1724,
  -66.1906,
  -66.2063,
  -66.2201,
  -66.2319,
  -66.2417,
  -66.2494,
  -66.2543,
  -66.2557,
  -66.2536,
  -66.2481,
  -66.2397,
  -66.2288,
  -66.2161,
  -66.2021,
  -66.1867,
  -66.1701,
  -66.1536,
  -66.1377,
  -66.1217,
  -66.1077,
  -66.0947,
  -66.0818,
  -66.0685,
  -66.0546,
  -66.0391,
  -66.0219,
  -66.0023,
  -65.9803,
  -65.9559,
  -65.9291,
  -65.9004,
  -65.8705,
  -65.8397,
  -65.8086,
  -65.7772,
  -65.7454,
  -65.7129,
  -65.68,
  -65.6465,
  -65.612,
  -65.5768,
  -65.5411,
  -65.5048,
  -65.4683,
  -65.4319,
  -65.3943,
  -65.358,
  -65.3218,
  -65.2858,
  -65.2492,
  -65.2122,
  -65.1745,
  -65.1363,
  -65.0976,
  -65.0588,
  -65.02,
  -64.9809,
  -64.9414,
  -64.9012,
  -64.8601,
  -64.8177,
  -64.7743,
  -64.7299,
  -64.6849,
  -64.639,
  -64.5921,
  -64.5443,
  -64.4956,
  -64.4464,
  -64.3968,
  -64.3467,
  -64.2958,
  -64.2438,
  -64.1909,
  -64.1366,
  -64.0811,
  -64.0245,
  -63.9653,
  -63.9051,
  -63.8424,
  -63.777,
  -63.7088,
  -63.6383,
  -63.5656,
  -63.4909,
  -63.4143,
  -63.3364,
  -63.258,
  -63.1798,
  -63.1023,
  -63.0263,
  -62.9517,
  -62.8777,
  -62.8037,
  -62.7287,
  -62.652,
  -62.5737,
  -62.4938,
  -62.4131,
  -62.3324,
  -62.2521,
  -62.1727,
  -62.0943,
  -62.0166,
  -61.939,
  -61.8608,
  -61.7813,
  -61.7004,
  -61.6184,
  -61.5357,
  -61.453,
  -61.3712,
  -61.2906,
  -61.2119,
  -61.135,
  -61.0589,
  -60.9856,
  -60.9151,
  -60.8447,
  -60.7773,
  -60.7114,
  -60.6469,
  -60.5831,
  -60.5204,
  -60.4591,
  -60.3999,
  -60.3432,
  -60.2894,
  -60.2385,
  -60.1906,
  -60.1455,
  -60.103,
  -60.0628,
  -60.0244,
  -59.9875,
  -59.9516,
  -59.9159,
  -59.8806,
  -59.8459,
  -59.8118,
  -59.7782,
  -59.7458,
  -49.3569,
  -49.3875,
  -49.4263,
  -49.4728,
  -49.5259,
  -49.5849,
  -49.653,
  -49.731,
  -49.8207,
  -49.9249,
  -50.0462,
  -50.1863,
  -50.3465,
  -50.5263,
  -50.7244,
  -50.9386,
  -51.1667,
  -51.4067,
  -51.6563,
  -51.913,
  -52.1741,
  -52.4397,
  -52.7078,
  -52.9776,
  -53.2484,
  -53.5202,
  -53.7932,
  -54.0671,
  -54.3415,
  -54.6163,
  -54.8905,
  -55.1634,
  -55.4333,
  -55.6983,
  -55.9558,
  -56.203,
  -56.4396,
  -56.6629,
  -56.8721,
  -57.0676,
  -57.2503,
  -57.4226,
  -57.5875,
  -57.7481,
  -57.9071,
  -58.0662,
  -58.2268,
  -58.3886,
  -58.5508,
  -58.7118,
  -58.8696,
  -59.0209,
  -59.1663,
  -59.3034,
  -59.432,
  -59.5524,
  -59.6653,
  -59.7717,
  -59.8724,
  -59.9679,
  -60.059,
  -60.1465,
  -60.2309,
  -60.3127,
  -60.3923,
  -60.4702,
  -60.5468,
  -60.6223,
  -60.6962,
  -60.7702,
  -60.8431,
  -60.9155,
  -60.9873,
  -61.0587,
  -61.1295,
  -61.1996,
  -61.2696,
  -61.3398,
  -61.4107,
  -61.4827,
  -61.5559,
  -61.6305,
  -61.7064,
  -61.7831,
  -61.8604,
  -61.9378,
  -62.0143,
  -62.0918,
  -62.1696,
  -62.2484,
  -62.3286,
  -62.4107,
  -62.4952,
  -62.5817,
  -62.6699,
  -62.7594,
  -62.8495,
  -62.9396,
  -63.029,
  -63.1175,
  -63.2047,
  -63.2906,
  -63.3757,
  -63.4598,
  -63.5435,
  -63.6246,
  -63.7054,
  -63.7845,
  -63.8616,
  -63.9376,
  -64.0119,
  -64.0845,
  -64.1556,
  -64.2256,
  -64.295,
  -64.3641,
  -64.433,
  -64.5017,
  -64.5692,
  -64.6352,
  -64.6993,
  -64.7614,
  -64.8211,
  -64.8789,
  -64.9357,
  -64.9904,
  -65.0459,
  -65.101,
  -65.1561,
  -65.2116,
  -65.2674,
  -65.3232,
  -65.3782,
  -65.4327,
  -65.4862,
  -65.5384,
  -65.5893,
  -65.6389,
  -65.6871,
  -65.734,
  -65.7796,
  -65.8241,
  -65.868,
  -65.9114,
  -65.9547,
  -65.9967,
  -66.0391,
  -66.0809,
  -66.1218,
  -66.1621,
  -66.2015,
  -66.2396,
  -66.2767,
  -66.3115,
  -66.3438,
  -66.373,
  -66.3993,
  -66.4225,
  -66.4425,
  -66.4597,
  -66.4739,
  -66.4855,
  -66.4946,
  -66.5016,
  -66.5061,
  -66.5076,
  -66.5059,
  -66.5005,
  -66.4908,
  -66.4791,
  -66.4649,
  -66.4486,
  -66.431,
  -66.412,
  -66.3925,
  -66.3729,
  -66.3535,
  -66.3353,
  -66.318,
  -66.3014,
  -66.2851,
  -66.2683,
  -66.2504,
  -66.2307,
  -66.2088,
  -66.1844,
  -66.1575,
  -66.128,
  -66.0964,
  -66.0631,
  -66.0288,
  -65.9938,
  -65.9588,
  -65.9236,
  -65.8875,
  -65.8518,
  -65.8157,
  -65.7792,
  -65.7424,
  -65.7051,
  -65.6673,
  -65.6299,
  -65.5927,
  -65.5555,
  -65.5187,
  -65.4824,
  -65.4468,
  -65.4111,
  -65.3752,
  -65.3389,
  -65.302,
  -65.2645,
  -65.2263,
  -65.1876,
  -65.1486,
  -65.1093,
  -65.0693,
  -65.0286,
  -64.987,
  -64.9443,
  -64.9005,
  -64.8556,
  -64.8098,
  -64.7632,
  -64.715,
  -64.6672,
  -64.6189,
  -64.5701,
  -64.521,
  -64.4713,
  -64.4207,
  -64.3689,
  -64.3158,
  -64.2616,
  -64.2059,
  -64.1491,
  -64.0907,
  -64.0301,
  -63.967,
  -63.9014,
  -63.8332,
  -63.7628,
  -63.6902,
  -63.6153,
  -63.5384,
  -63.46,
  -63.3807,
  -63.3017,
  -63.2237,
  -63.1475,
  -63.073,
  -62.9991,
  -62.9252,
  -62.8503,
  -62.7738,
  -62.6956,
  -62.6159,
  -62.5354,
  -62.4548,
  -62.3737,
  -62.2948,
  -62.2169,
  -62.1395,
  -62.0621,
  -61.984,
  -61.9044,
  -61.8233,
  -61.741,
  -61.6578,
  -61.5746,
  -61.492,
  -61.4104,
  -61.3305,
  -61.2525,
  -61.1765,
  -61.1027,
  -61.0309,
  -60.9612,
  -60.8934,
  -60.8273,
  -60.7625,
  -60.699,
  -60.6364,
  -60.5757,
  -60.5174,
  -60.4616,
  -60.4089,
  -60.3593,
  -60.3126,
  -60.2687,
  -60.2276,
  -60.1887,
  -60.1518,
  -60.1162,
  -60.0817,
  -60.0477,
  -60.0141,
  -59.9809,
  -59.948,
  -59.9159,
  -59.8849,
  -49.5916,
  -49.6306,
  -49.6754,
  -49.7254,
  -49.7807,
  -49.8419,
  -49.9112,
  -49.9911,
  -50.084,
  -50.1927,
  -50.3196,
  -50.4662,
  -50.6327,
  -50.8186,
  -51.0218,
  -51.2389,
  -51.4692,
  -51.7098,
  -51.9586,
  -52.2134,
  -52.4726,
  -52.7346,
  -52.9988,
  -53.2649,
  -53.5317,
  -53.7995,
  -54.0686,
  -54.3386,
  -54.6093,
  -54.8804,
  -55.1507,
  -55.4217,
  -55.6912,
  -55.9571,
  -56.2169,
  -56.4683,
  -56.7087,
  -56.9362,
  -57.1495,
  -57.3487,
  -57.5345,
  -57.7094,
  -57.8761,
  -58.0375,
  -58.1965,
  -58.355,
  -58.5132,
  -58.673,
  -58.8327,
  -58.9909,
  -59.1459,
  -59.2958,
  -59.439,
  -59.5747,
  -59.7024,
  -59.8224,
  -59.9353,
  -60.0423,
  -60.1435,
  -60.2394,
  -60.331,
  -60.4188,
  -60.5025,
  -60.5847,
  -60.6649,
  -60.7434,
  -60.8209,
  -60.8974,
  -60.9732,
  -61.0482,
  -61.1224,
  -61.1959,
  -61.2684,
  -61.3409,
  -61.4126,
  -61.4838,
  -61.5544,
  -61.6253,
  -61.6967,
  -61.7682,
  -61.8417,
  -61.9167,
  -61.9926,
  -62.0695,
  -62.1465,
  -62.2238,
  -62.3009,
  -62.3779,
  -62.4552,
  -62.5331,
  -62.6127,
  -62.6941,
  -62.778,
  -62.8646,
  -62.9532,
  -63.0434,
  -63.1341,
  -63.2247,
  -63.3137,
  -63.4028,
  -63.4908,
  -63.5778,
  -63.6642,
  -63.7499,
  -63.8348,
  -63.9188,
  -64.0013,
  -64.082,
  -64.1614,
  -64.2391,
  -64.3149,
  -64.3885,
  -64.4598,
  -64.5293,
  -64.5977,
  -64.6656,
  -64.7321,
  -64.7992,
  -64.8654,
  -64.9306,
  -64.9942,
  -65.0561,
  -65.1159,
  -65.1737,
  -65.2298,
  -65.2844,
  -65.338,
  -65.391,
  -65.4439,
  -65.4971,
  -65.5506,
  -65.6047,
  -65.6584,
  -65.7119,
  -65.7643,
  -65.8155,
  -65.8654,
  -65.9129,
  -65.9598,
  -66.0054,
  -66.0496,
  -66.0929,
  -66.1358,
  -66.1784,
  -66.2212,
  -66.264,
  -66.3058,
  -66.3462,
  -66.3853,
  -66.4235,
  -66.461,
  -66.4977,
  -66.5336,
  -66.5678,
  -66.5999,
  -66.6292,
  -66.6554,
  -66.6784,
  -66.6981,
  -66.7144,
  -66.7264,
  -66.7362,
  -66.743,
  -66.7473,
  -66.7487,
  -66.7472,
  -66.7423,
  -66.7339,
  -66.7216,
  -66.7066,
  -66.6892,
  -66.6695,
  -66.6482,
  -66.6257,
  -66.603,
  -66.58,
  -66.5576,
  -66.536,
  -66.5154,
  -66.4957,
  -66.476,
  -66.4558,
  -66.434,
  -66.4101,
  -66.3837,
  -66.3535,
  -66.3217,
  -66.2876,
  -66.2513,
  -66.2135,
  -66.1748,
  -66.1356,
  -66.0966,
  -66.0577,
  -66.0188,
  -65.9799,
  -65.9406,
  -65.901,
  -65.8614,
  -65.8215,
  -65.7818,
  -65.7427,
  -65.7041,
  -65.6662,
  -65.6291,
  -65.5928,
  -65.5575,
  -65.5227,
  -65.4879,
  -65.4527,
  -65.4168,
  -65.3801,
  -65.3426,
  -65.3031,
  -65.2638,
  -65.2239,
  -65.1834,
  -65.1424,
  -65.1007,
  -65.0579,
  -65.0139,
  -64.9685,
  -64.9217,
  -64.8742,
  -64.8265,
  -64.7785,
  -64.7303,
  -64.6821,
  -64.6335,
  -64.5841,
  -64.5334,
  -64.4814,
  -64.428,
  -64.3732,
  -64.3171,
  -64.2596,
  -64.2004,
  -64.1392,
  -64.0756,
  -64.0097,
  -63.9417,
  -63.8713,
  -63.7988,
  -63.7238,
  -63.6464,
  -63.5674,
  -63.4864,
  -63.4067,
  -63.3282,
  -63.2516,
  -63.1767,
  -63.1027,
  -63.0288,
  -62.9538,
  -62.8772,
  -62.799,
  -62.7196,
  -62.6394,
  -62.5593,
  -62.4799,
  -62.4015,
  -62.324,
  -62.2467,
  -62.1692,
  -62.0909,
  -62.011,
  -61.9295,
  -61.8466,
  -61.7629,
  -61.679,
  -61.5955,
  -61.5129,
  -61.4317,
  -61.3524,
  -61.2754,
  -61.2007,
  -61.1285,
  -61.0581,
  -60.9896,
  -60.923,
  -60.8582,
  -60.7947,
  -60.7329,
  -60.6734,
  -60.6162,
  -60.5621,
  -60.5109,
  -60.4619,
  -60.4168,
  -60.374,
  -60.3338,
  -60.2961,
  -60.2604,
  -60.2262,
  -60.1934,
  -60.1609,
  -60.1291,
  -60.0976,
  -60.0665,
  -60.0362,
  -60.0065,
  -49.8195,
  -49.8666,
  -49.9172,
  -49.9711,
  -50.0294,
  -50.0934,
  -50.1653,
  -50.2484,
  -50.3457,
  -50.4587,
  -50.5919,
  -50.7448,
  -50.9174,
  -51.1086,
  -51.3159,
  -51.5364,
  -51.7678,
  -52.008,
  -52.2548,
  -52.5066,
  -52.7622,
  -53.0206,
  -53.281,
  -53.5431,
  -53.8053,
  -54.0704,
  -54.3366,
  -54.6039,
  -54.872,
  -55.1409,
  -55.4108,
  -55.6809,
  -55.9503,
  -56.2172,
  -56.4792,
  -56.7332,
  -56.9766,
  -57.2072,
  -57.4235,
  -57.6255,
  -57.813,
  -57.9899,
  -58.1582,
  -58.3209,
  -58.4801,
  -58.6381,
  -58.7957,
  -58.9532,
  -59.1098,
  -59.2644,
  -59.4155,
  -59.5618,
  -59.7019,
  -59.835,
  -59.961,
  -60.08,
  -60.1918,
  -60.2984,
  -60.3998,
  -60.496,
  -60.5879,
  -60.676,
  -60.7608,
  -60.8433,
  -60.9238,
  -61.0028,
  -61.0809,
  -61.1584,
  -61.2352,
  -61.3113,
  -61.3867,
  -61.4609,
  -61.5345,
  -61.6068,
  -61.6793,
  -61.7512,
  -61.8227,
  -61.8943,
  -61.9664,
  -62.0393,
  -62.1134,
  -62.1889,
  -62.2653,
  -62.3424,
  -62.4195,
  -62.4964,
  -62.5733,
  -62.65,
  -62.7269,
  -62.8047,
  -62.8837,
  -62.9638,
  -63.0475,
  -63.134,
  -63.2226,
  -63.313,
  -63.404,
  -63.4948,
  -63.585,
  -63.6746,
  -63.7632,
  -63.851,
  -63.9384,
  -64.0252,
  -64.1114,
  -64.1965,
  -64.2805,
  -64.3632,
  -64.4444,
  -64.523,
  -64.6001,
  -64.6745,
  -64.746,
  -64.815,
  -64.8825,
  -64.949,
  -65.015,
  -65.0802,
  -65.145,
  -65.209,
  -65.2718,
  -65.3331,
  -65.3923,
  -65.4501,
  -65.5057,
  -65.5593,
  -65.6116,
  -65.6629,
  -65.714,
  -65.7654,
  -65.8163,
  -65.8687,
  -65.9213,
  -65.9736,
  -66.0252,
  -66.0756,
  -66.1245,
  -66.1718,
  -66.2178,
  -66.2622,
  -66.3056,
  -66.3478,
  -66.3896,
  -66.4319,
  -66.4741,
  -66.5161,
  -66.557,
  -66.5962,
  -66.6341,
  -66.6708,
  -66.7066,
  -66.7407,
  -66.7753,
  -66.8088,
  -66.8403,
  -66.8694,
  -66.8957,
  -66.9187,
  -66.938,
  -66.9537,
  -66.9655,
  -66.9735,
  -66.9781,
  -66.9797,
  -66.9782,
  -66.9736,
  -66.9657,
  -66.9541,
  -66.9389,
  -66.9208,
  -66.9002,
  -66.8773,
  -66.8524,
  -66.827,
  -66.8011,
  -66.7745,
  -66.7491,
  -66.7244,
  -66.7006,
  -66.6775,
  -66.6544,
  -66.6304,
  -66.6046,
  -66.5765,
  -66.5456,
  -66.5121,
  -66.4758,
  -66.4372,
  -66.3966,
  -66.3546,
  -66.3115,
  -66.2682,
  -66.225,
  -66.1825,
  -66.14,
  -66.0975,
  -66.0549,
  -66.012,
  -65.9693,
  -65.9267,
  -65.8846,
  -65.8437,
  -65.8028,
  -65.7641,
  -65.7266,
  -65.6903,
  -65.6552,
  -65.6209,
  -65.5868,
  -65.5525,
  -65.5176,
  -65.4816,
  -65.4444,
  -65.406,
  -65.3665,
  -65.3262,
  -65.2852,
  -65.2441,
  -65.2026,
  -65.1597,
  -65.1153,
  -65.0691,
  -65.0215,
  -64.9734,
  -64.925,
  -64.8766,
  -64.8286,
  -64.7807,
  -64.7321,
  -64.6826,
  -64.6316,
  -64.5791,
  -64.5249,
  -64.4685,
  -64.4116,
  -64.3532,
  -64.2932,
  -64.2311,
  -64.1674,
  -64.1015,
  -64.0335,
  -63.9633,
  -63.8908,
  -63.8156,
  -63.738,
  -63.6584,
  -63.5776,
  -63.4969,
  -63.4177,
  -63.3403,
  -63.2646,
  -63.1898,
  -63.1153,
  -63.0401,
  -62.9635,
  -62.8856,
  -62.8066,
  -62.7269,
  -62.6474,
  -62.5685,
  -62.4905,
  -62.4131,
  -62.3361,
  -62.2583,
  -62.1797,
  -62.0994,
  -62.0174,
  -61.9341,
  -61.8498,
  -61.7651,
  -61.6807,
  -61.596,
  -61.5135,
  -61.4332,
  -61.3551,
  -61.2795,
  -61.2061,
  -61.1349,
  -61.0657,
  -60.9984,
  -60.9334,
  -60.8703,
  -60.8095,
  -60.7512,
  -60.6957,
  -60.6433,
  -60.594,
  -60.5478,
  -60.5037,
  -60.4623,
  -60.4233,
  -60.3867,
  -60.3523,
  -60.3198,
  -60.2887,
  -60.2584,
  -60.2285,
  -60.1988,
  -60.1695,
  -60.1408,
  -60.1127,
  -50.0334,
  -50.0878,
  -50.1447,
  -50.2038,
  -50.2653,
  -50.3335,
  -50.4101,
  -50.4983,
  -50.6014,
  -50.7218,
  -50.8615,
  -51.0208,
  -51.199,
  -51.3946,
  -51.6046,
  -51.8266,
  -52.0577,
  -52.2958,
  -52.5397,
  -52.7865,
  -53.038,
  -53.292,
  -53.5485,
  -53.8068,
  -54.0678,
  -54.3301,
  -54.5945,
  -54.8605,
  -55.1277,
  -55.3962,
  -55.6658,
  -55.9362,
  -56.2065,
  -56.4747,
  -56.7373,
  -56.9933,
  -57.2387,
  -57.4711,
  -57.6892,
  -57.8928,
  -58.0832,
  -58.2619,
  -58.4318,
  -58.5954,
  -58.7551,
  -58.9127,
  -59.0688,
  -59.2238,
  -59.3771,
  -59.5276,
  -59.6735,
  -59.8155,
  -59.9516,
  -60.0816,
  -60.2053,
  -60.3229,
  -60.4346,
  -60.5408,
  -60.642,
  -60.7381,
  -60.8301,
  -60.9182,
  -61.0031,
  -61.0855,
  -61.1661,
  -61.2455,
  -61.3242,
  -61.4014,
  -61.4792,
  -61.5563,
  -61.6328,
  -61.7083,
  -61.7828,
  -61.8565,
  -61.9297,
  -62.0026,
  -62.0749,
  -62.1473,
  -62.2201,
  -62.2938,
  -62.3686,
  -62.4446,
  -62.5215,
  -62.5989,
  -62.6761,
  -62.7522,
  -62.8289,
  -62.9055,
  -62.9823,
  -63.0601,
  -63.139,
  -63.2199,
  -63.3035,
  -63.3898,
  -63.4783,
  -63.5685,
  -63.6594,
  -63.7503,
  -63.8404,
  -63.93,
  -64.0191,
  -64.1075,
  -64.1945,
  -64.2823,
  -64.3693,
  -64.4555,
  -64.5408,
  -64.6249,
  -64.7079,
  -64.7889,
  -64.8675,
  -64.9425,
  -65.0145,
  -65.0832,
  -65.1499,
  -65.2152,
  -65.2796,
  -65.343,
  -65.4059,
  -65.4683,
  -65.5298,
  -65.5902,
  -65.6485,
  -65.7057,
  -65.7604,
  -65.8134,
  -65.8648,
  -65.9149,
  -65.9647,
  -66.0146,
  -66.0652,
  -66.1165,
  -66.1683,
  -66.2196,
  -66.2703,
  -66.3197,
  -66.3677,
  -66.4143,
  -66.4594,
  -66.5033,
  -66.5459,
  -66.5878,
  -66.6294,
  -66.6699,
  -66.7113,
  -66.7524,
  -66.7924,
  -66.8307,
  -66.8672,
  -66.9023,
  -66.9367,
  -66.9705,
  -67.0039,
  -67.0364,
  -67.0673,
  -67.096,
  -67.122,
  -67.1446,
  -67.1635,
  -67.1783,
  -67.189,
  -67.1954,
  -67.1981,
  -67.197,
  -67.1923,
  -67.1848,
  -67.1742,
  -67.159,
  -67.1411,
  -67.1203,
  -67.097,
  -67.0714,
  -67.0438,
  -67.0154,
  -66.9869,
  -66.9586,
  -66.9304,
  -66.9028,
  -66.8757,
  -66.8491,
  -66.8222,
  -66.7943,
  -66.7645,
  -66.7322,
  -66.6971,
  -66.6592,
  -66.6187,
  -66.5758,
  -66.531,
  -66.4847,
  -66.4376,
  -66.3902,
  -66.3422,
  -66.2957,
  -66.2495,
  -66.2034,
  -66.1573,
  -66.1111,
  -66.065,
  -66.0195,
  -65.9752,
  -65.9323,
  -65.8913,
  -65.8519,
  -65.8142,
  -65.7779,
  -65.7427,
  -65.7086,
  -65.6746,
  -65.6406,
  -65.6062,
  -65.5704,
  -65.5335,
  -65.4948,
  -65.4549,
  -65.4143,
  -65.3733,
  -65.332,
  -65.2903,
  -65.2471,
  -65.2023,
  -65.1546,
  -65.1066,
  -65.0574,
  -65.0082,
  -64.9596,
  -64.9113,
  -64.8631,
  -64.8143,
  -64.7644,
  -64.7129,
  -64.6597,
  -64.6048,
  -64.5485,
  -64.4908,
  -64.4315,
  -64.3708,
  -64.3084,
  -64.2443,
  -64.1784,
  -64.1108,
  -64.0409,
  -63.9684,
  -63.8929,
  -63.815,
  -63.7347,
  -63.6532,
  -63.5715,
  -63.4911,
  -63.4123,
  -63.3352,
  -63.2593,
  -63.184,
  -63.1081,
  -63.0314,
  -62.9539,
  -62.8744,
  -62.7954,
  -62.7166,
  -62.6382,
  -62.5608,
  -62.4836,
  -62.4062,
  -62.3282,
  -62.2491,
  -62.1686,
  -62.0861,
  -62.0022,
  -61.9173,
  -61.8318,
  -61.7465,
  -61.6617,
  -61.5783,
  -61.4967,
  -61.4174,
  -61.3405,
  -61.2662,
  -61.194,
  -61.124,
  -61.0563,
  -60.9912,
  -60.9285,
  -60.8687,
  -60.8119,
  -60.7583,
  -60.7078,
  -60.6604,
  -60.6158,
  -60.5733,
  -60.5329,
  -60.4949,
  -60.4592,
  -60.4262,
  -60.3955,
  -60.3665,
  -60.3383,
  -60.3104,
  -60.2827,
  -60.2553,
  -60.2282,
  -60.2019,
  -50.2265,
  -50.2886,
  -50.3524,
  -50.4182,
  -50.4872,
  -50.5616,
  -50.6445,
  -50.7396,
  -50.8497,
  -50.9772,
  -51.1235,
  -51.2887,
  -51.4717,
  -51.6698,
  -51.8819,
  -52.1041,
  -52.3337,
  -52.5689,
  -52.8088,
  -53.0521,
  -53.2989,
  -53.5485,
  -53.801,
  -54.0564,
  -54.3148,
  -54.5758,
  -54.8393,
  -55.1048,
  -55.3726,
  -55.641,
  -55.9117,
  -56.1834,
  -56.4551,
  -56.7248,
  -56.9898,
  -57.2468,
  -57.493,
  -57.726,
  -57.9445,
  -58.149,
  -58.3402,
  -58.5201,
  -58.6912,
  -58.8559,
  -59.015,
  -59.1722,
  -59.3271,
  -59.4798,
  -59.6297,
  -59.7763,
  -59.9186,
  -60.0559,
  -60.1879,
  -60.3143,
  -60.4352,
  -60.551,
  -60.6615,
  -60.7668,
  -60.8674,
  -60.9634,
  -61.0551,
  -61.1421,
  -61.2268,
  -61.3091,
  -61.3896,
  -61.4692,
  -61.5482,
  -61.6272,
  -61.7058,
  -61.784,
  -61.8614,
  -61.9378,
  -62.0133,
  -62.0879,
  -62.162,
  -62.2356,
  -62.3088,
  -62.381,
  -62.4548,
  -62.5293,
  -62.6048,
  -62.6814,
  -62.7587,
  -62.8366,
  -62.9143,
  -62.9915,
  -63.0683,
  -63.145,
  -63.222,
  -63.2997,
  -63.3789,
  -63.46,
  -63.5435,
  -63.6295,
  -63.7175,
  -63.8061,
  -63.8964,
  -63.9869,
  -64.0772,
  -64.1668,
  -64.2559,
  -64.3448,
  -64.4332,
  -64.5212,
  -64.6088,
  -64.6959,
  -64.7824,
  -64.8681,
  -64.9523,
  -65.0347,
  -65.1143,
  -65.1902,
  -65.2625,
  -65.3314,
  -65.3978,
  -65.4612,
  -65.5241,
  -65.586,
  -65.6471,
  -65.7076,
  -65.7679,
  -65.8272,
  -65.8855,
  -65.9419,
  -65.9963,
  -66.0485,
  -66.0992,
  -66.1489,
  -66.1979,
  -66.247,
  -66.2967,
  -66.3469,
  -66.3978,
  -66.4484,
  -66.498,
  -66.5466,
  -66.5925,
  -66.6384,
  -66.6831,
  -66.7269,
  -66.7697,
  -66.8116,
  -66.8533,
  -66.8944,
  -66.9353,
  -66.9753,
  -67.0141,
  -67.0512,
  -67.0867,
  -67.1209,
  -67.1541,
  -67.1863,
  -67.2181,
  -67.2491,
  -67.2788,
  -67.3065,
  -67.3315,
  -67.3536,
  -67.3709,
  -67.3851,
  -67.3946,
  -67.3993,
  -67.4001,
  -67.3969,
  -67.3898,
  -67.3796,
  -67.3664,
  -67.3499,
  -67.3297,
  -67.3064,
  -67.2807,
  -67.2528,
  -67.2232,
  -67.1929,
  -67.1623,
  -67.1318,
  -67.1012,
  -67.0707,
  -67.0404,
  -67.0101,
  -66.9792,
  -66.9471,
  -66.9132,
  -66.8753,
  -66.8359,
  -66.7939,
  -66.7493,
  -66.7027,
  -66.6541,
  -66.6036,
  -66.5522,
  -66.5007,
  -66.4499,
  -66.3997,
  -66.3498,
  -66.3001,
  -66.2503,
  -66.2003,
  -66.151,
  -66.1024,
  -66.0556,
  -66.0108,
  -65.9684,
  -65.9283,
  -65.8903,
  -65.8539,
  -65.8187,
  -65.7844,
  -65.7503,
  -65.7159,
  -65.681,
  -65.6441,
  -65.6068,
  -65.5678,
  -65.5279,
  -65.4871,
  -65.4459,
  -65.4044,
  -65.3622,
  -65.3186,
  -65.2731,
  -65.2256,
  -65.1766,
  -65.1268,
  -65.0773,
  -65.0281,
  -64.9791,
  -64.9303,
  -64.8811,
  -64.8306,
  -64.7784,
  -64.7244,
  -64.6688,
  -64.6119,
  -64.5536,
  -64.4937,
  -64.4324,
  -64.3696,
  -64.3055,
  -64.24,
  -64.1726,
  -64.1028,
  -64.0304,
  -63.9538,
  -63.8755,
  -63.7946,
  -63.7122,
  -63.6297,
  -63.5477,
  -63.4671,
  -63.3881,
  -63.3106,
  -63.2341,
  -63.1575,
  -63.0807,
  -63.0031,
  -62.9249,
  -62.8465,
  -62.7683,
  -62.6906,
  -62.6133,
  -62.536,
  -62.4586,
  -62.3803,
  -62.3008,
  -62.2199,
  -62.1371,
  -62.0529,
  -61.9674,
  -61.8813,
  -61.7951,
  -61.7094,
  -61.6249,
  -61.5421,
  -61.4615,
  -61.3833,
  -61.3078,
  -61.2347,
  -61.1641,
  -61.0964,
  -61.0316,
  -60.9697,
  -60.911,
  -60.8555,
  -60.8026,
  -60.754,
  -60.7084,
  -60.6653,
  -60.6242,
  -60.5849,
  -60.5478,
  -60.5135,
  -60.4821,
  -60.4532,
  -60.4263,
  -60.4003,
  -60.3745,
  -60.3486,
  -60.3231,
  -60.2979,
  -60.2735,
  -50.3972,
  -50.4678,
  -50.5395,
  -50.6131,
  -50.69,
  -50.7726,
  -50.8639,
  -50.9672,
  -51.0843,
  -51.2193,
  -51.3722,
  -51.5428,
  -51.7299,
  -51.9316,
  -52.1444,
  -52.3658,
  -52.5932,
  -52.825,
  -53.0607,
  -53.2997,
  -53.5419,
  -53.7876,
  -54.0367,
  -54.2884,
  -54.5452,
  -54.8053,
  -55.0687,
  -55.3351,
  -55.6042,
  -55.8755,
  -56.1483,
  -56.4219,
  -56.6952,
  -56.966,
  -57.2315,
  -57.4887,
  -57.7344,
  -57.9668,
  -58.1848,
  -58.3879,
  -58.5793,
  -58.7599,
  -58.9317,
  -59.0969,
  -59.2573,
  -59.4143,
  -59.5681,
  -59.7187,
  -59.8657,
  -60.0084,
  -60.1465,
  -60.2794,
  -60.4072,
  -60.5301,
  -60.6482,
  -60.7608,
  -60.8698,
  -60.9742,
  -61.0742,
  -61.1699,
  -61.2612,
  -61.3488,
  -61.4331,
  -61.515,
  -61.5953,
  -61.6749,
  -61.7541,
  -61.8333,
  -61.9126,
  -61.9916,
  -62.0701,
  -62.1467,
  -62.2233,
  -62.2988,
  -62.3738,
  -62.4482,
  -62.5221,
  -62.5961,
  -62.6708,
  -62.7463,
  -62.8228,
  -62.9,
  -62.9778,
  -63.056,
  -63.1339,
  -63.2114,
  -63.2886,
  -63.3655,
  -63.4428,
  -63.5202,
  -63.5999,
  -63.6814,
  -63.7649,
  -63.8505,
  -63.9379,
  -64.0265,
  -64.116,
  -64.2057,
  -64.2956,
  -64.385,
  -64.4743,
  -64.5628,
  -64.6515,
  -64.7395,
  -64.8275,
  -64.9152,
  -65.0028,
  -65.0895,
  -65.174,
  -65.2573,
  -65.3378,
  -65.4146,
  -65.4874,
  -65.5567,
  -65.6233,
  -65.6874,
  -65.7496,
  -65.8102,
  -65.8699,
  -65.9292,
  -65.9882,
  -66.0465,
  -66.1037,
  -66.1593,
  -66.213,
  -66.2647,
  -66.3149,
  -66.3641,
  -66.4116,
  -66.46,
  -66.5088,
  -66.5584,
  -66.6084,
  -66.6579,
  -66.7068,
  -66.7547,
  -66.8016,
  -66.8472,
  -66.892,
  -66.9362,
  -66.9793,
  -67.0217,
  -67.0632,
  -67.104,
  -67.1441,
  -67.1831,
  -67.2205,
  -67.2564,
  -67.2907,
  -67.324,
  -67.355,
  -67.3858,
  -67.4159,
  -67.4451,
  -67.473,
  -67.4993,
  -67.5229,
  -67.5438,
  -67.5609,
  -67.5744,
  -67.583,
  -67.5867,
  -67.586,
  -67.5809,
  -67.5721,
  -67.5598,
  -67.5443,
  -67.5255,
  -67.5031,
  -67.4777,
  -67.4497,
  -67.4197,
  -67.3883,
  -67.3562,
  -67.323,
  -67.291,
  -67.2585,
  -67.2257,
  -67.1925,
  -67.159,
  -67.1244,
  -67.0884,
  -67.0503,
  -67.0091,
  -66.9653,
  -66.9191,
  -66.8707,
  -66.8203,
  -66.7676,
  -66.7134,
  -66.6583,
  -66.6028,
  -66.5478,
  -66.4935,
  -66.4397,
  -66.3859,
  -66.3325,
  -66.2791,
  -66.2264,
  -66.1751,
  -66.1246,
  -66.0777,
  -66.0338,
  -65.9923,
  -65.9532,
  -65.9159,
  -65.8803,
  -65.8455,
  -65.8105,
  -65.7757,
  -65.7403,
  -65.7037,
  -65.666,
  -65.6269,
  -65.5867,
  -65.5457,
  -65.5043,
  -65.4623,
  -65.4195,
  -65.3751,
  -65.3286,
  -65.2803,
  -65.2306,
  -65.1802,
  -65.1299,
  -65.0799,
  -65.0304,
  -64.9809,
  -64.9308,
  -64.8795,
  -64.8266,
  -64.7711,
  -64.715,
  -64.6574,
  -64.5987,
  -64.5386,
  -64.477,
  -64.4143,
  -64.3503,
  -64.2851,
  -64.2181,
  -64.1486,
  -64.0762,
  -64.0005,
  -63.9218,
  -63.8402,
  -63.7569,
  -63.6728,
  -63.5892,
  -63.5068,
  -63.4259,
  -63.3468,
  -63.2688,
  -63.1916,
  -63.1143,
  -63.0364,
  -62.9583,
  -62.8799,
  -62.8016,
  -62.7238,
  -62.6463,
  -62.5688,
  -62.4908,
  -62.412,
  -62.3325,
  -62.2514,
  -62.1688,
  -62.0847,
  -61.9981,
  -61.9116,
  -61.8249,
  -61.7383,
  -61.6527,
  -61.5686,
  -61.4865,
  -61.4069,
  -61.3301,
  -61.2563,
  -61.1855,
  -61.1182,
  -61.0542,
  -60.9934,
  -60.936,
  -60.882,
  -60.8315,
  -60.7844,
  -60.7404,
  -60.6988,
  -60.6589,
  -60.621,
  -60.5854,
  -60.5525,
  -60.5225,
  -60.4955,
  -60.4704,
  -60.4461,
  -60.4223,
  -60.3987,
  -60.3753,
  -60.3524,
  -60.3299,
  -50.5419,
  -50.6218,
  -50.7022,
  -50.7838,
  -50.87,
  -50.9622,
  -51.0633,
  -51.176,
  -51.3028,
  -51.4455,
  -51.6047,
  -51.78,
  -51.9705,
  -52.1739,
  -52.3871,
  -52.6073,
  -52.8322,
  -53.0606,
  -53.2916,
  -53.5266,
  -53.7649,
  -54.0072,
  -54.2537,
  -54.5044,
  -54.7601,
  -55.0202,
  -55.2842,
  -55.552,
  -55.8233,
  -56.0971,
  -56.3725,
  -56.6483,
  -56.923,
  -57.1934,
  -57.4585,
  -57.7145,
  -57.9586,
  -58.1892,
  -58.4056,
  -58.6084,
  -58.7992,
  -58.9796,
  -59.1517,
  -59.3173,
  -59.4779,
  -59.6345,
  -59.7874,
  -59.9363,
  -60.0807,
  -60.2193,
  -60.3535,
  -60.4826,
  -60.6067,
  -60.7263,
  -60.8417,
  -60.9533,
  -61.0608,
  -61.1642,
  -61.2634,
  -61.3584,
  -61.4492,
  -61.5362,
  -61.62,
  -61.7014,
  -61.7813,
  -61.8594,
  -61.9385,
  -62.0179,
  -62.0976,
  -62.1773,
  -62.2568,
  -62.3356,
  -62.4131,
  -62.4896,
  -62.5653,
  -62.6404,
  -62.7154,
  -62.7904,
  -62.8662,
  -62.9427,
  -63.0203,
  -63.0982,
  -63.1755,
  -63.2539,
  -63.3321,
  -63.41,
  -63.4877,
  -63.5654,
  -63.6435,
  -63.7227,
  -63.8029,
  -63.8852,
  -63.9687,
  -64.0539,
  -64.1404,
  -64.2279,
  -64.316,
  -64.4046,
  -64.4936,
  -64.5826,
  -64.6714,
  -64.7589,
  -64.8474,
  -64.9357,
  -65.0239,
  -65.1124,
  -65.2007,
  -65.2882,
  -65.3743,
  -65.4582,
  -65.5393,
  -65.6169,
  -65.6904,
  -65.7605,
  -65.8275,
  -65.8919,
  -65.954,
  -66.0141,
  -66.0733,
  -66.1316,
  -66.1892,
  -66.2453,
  -66.3015,
  -66.3563,
  -66.4095,
  -66.4607,
  -66.5105,
  -66.5591,
  -66.607,
  -66.6549,
  -66.7029,
  -66.7518,
  -66.801,
  -66.85,
  -66.8985,
  -66.946,
  -66.993,
  -67.0389,
  -67.0841,
  -67.1289,
  -67.1725,
  -67.2153,
  -67.256,
  -67.2965,
  -67.3358,
  -67.3736,
  -67.4098,
  -67.4444,
  -67.4776,
  -67.5097,
  -67.5403,
  -67.5699,
  -67.5985,
  -67.6259,
  -67.6519,
  -67.6763,
  -67.6986,
  -67.7179,
  -67.7337,
  -67.7456,
  -67.7533,
  -67.756,
  -67.7541,
  -67.748,
  -67.7378,
  -67.7228,
  -67.7054,
  -67.6845,
  -67.6601,
  -67.6327,
  -67.6025,
  -67.5711,
  -67.5383,
  -67.505,
  -67.4716,
  -67.438,
  -67.4041,
  -67.369,
  -67.3332,
  -67.2966,
  -67.2585,
  -67.2189,
  -67.1772,
  -67.1322,
  -67.0846,
  -67.0348,
  -66.9827,
  -66.9283,
  -66.8718,
  -66.8135,
  -66.7535,
  -66.6943,
  -66.6355,
  -66.5771,
  -66.5191,
  -66.4612,
  -66.4039,
  -66.3471,
  -66.2914,
  -66.2372,
  -66.1852,
  -66.1362,
  -66.09,
  -66.0467,
  -66.0059,
  -65.9672,
  -65.93,
  -65.8938,
  -65.8577,
  -65.8217,
  -65.7853,
  -65.7482,
  -65.7102,
  -65.6709,
  -65.6306,
  -65.5893,
  -65.5475,
  -65.5047,
  -65.4608,
  -65.4143,
  -65.3668,
  -65.3178,
  -65.2672,
  -65.2163,
  -65.1653,
  -65.1147,
  -65.0641,
  -65.0136,
  -64.9626,
  -64.9104,
  -64.8568,
  -64.8018,
  -64.7453,
  -64.6875,
  -64.6285,
  -64.5682,
  -64.5068,
  -64.4441,
  -64.3804,
  -64.3155,
  -64.2488,
  -64.1796,
  -64.1071,
  -64.0314,
  -63.952,
  -63.8697,
  -63.7854,
  -63.7001,
  -63.6149,
  -63.5305,
  -63.4477,
  -63.367,
  -63.2878,
  -63.2087,
  -63.1305,
  -63.052,
  -62.9733,
  -62.8946,
  -62.816,
  -62.7375,
  -62.6592,
  -62.581,
  -62.5023,
  -62.4231,
  -62.3433,
  -62.2624,
  -62.1802,
  -62.0965,
  -62.0112,
  -61.9246,
  -61.8375,
  -61.7504,
  -61.6639,
  -61.5785,
  -61.495,
  -61.414,
  -61.3362,
  -61.2619,
  -61.1912,
  -61.1247,
  -61.062,
  -61.0029,
  -60.9472,
  -60.8948,
  -60.8458,
  -60.8001,
  -60.7573,
  -60.7169,
  -60.6785,
  -60.6419,
  -60.6076,
  -60.5762,
  -60.5478,
  -60.5224,
  -60.4986,
  -60.4763,
  -60.4547,
  -60.4334,
  -60.4108,
  -60.3903,
  -60.3705,
  -50.6576,
  -50.7476,
  -50.8379,
  -50.9301,
  -51.0264,
  -51.1292,
  -51.2406,
  -51.3632,
  -51.499,
  -51.6493,
  -51.8146,
  -51.9945,
  -52.1864,
  -52.3909,
  -52.604,
  -52.823,
  -53.0457,
  -53.2713,
  -53.5003,
  -53.7325,
  -53.9683,
  -54.2084,
  -54.4532,
  -54.703,
  -54.9583,
  -55.2191,
  -55.4845,
  -55.7534,
  -56.0273,
  -56.3038,
  -56.5816,
  -56.8592,
  -57.1348,
  -57.4059,
  -57.6695,
  -57.9232,
  -58.1645,
  -58.3921,
  -58.6059,
  -58.8068,
  -58.9963,
  -59.176,
  -59.3468,
  -59.5124,
  -59.673,
  -59.8292,
  -59.9813,
  -60.1287,
  -60.2711,
  -60.4079,
  -60.5391,
  -60.6651,
  -60.7863,
  -60.9031,
  -61.0163,
  -61.126,
  -61.2322,
  -61.3347,
  -61.4331,
  -61.5263,
  -61.6163,
  -61.7026,
  -61.7855,
  -61.8662,
  -61.9456,
  -62.0241,
  -62.1029,
  -62.1822,
  -62.2623,
  -62.3424,
  -62.4224,
  -62.502,
  -62.5804,
  -62.6578,
  -62.7342,
  -62.8101,
  -62.8852,
  -62.9615,
  -63.0385,
  -63.1164,
  -63.1947,
  -63.2734,
  -63.3522,
  -63.431,
  -63.5097,
  -63.5883,
  -63.6669,
  -63.7456,
  -63.8248,
  -63.905,
  -63.9866,
  -64.0692,
  -64.1531,
  -64.2378,
  -64.3222,
  -64.4083,
  -64.4949,
  -64.582,
  -64.6698,
  -64.7579,
  -64.8463,
  -64.9347,
  -65.023,
  -65.1116,
  -65.2004,
  -65.2893,
  -65.3778,
  -65.4656,
  -65.5519,
  -65.6359,
  -65.7174,
  -65.7956,
  -65.87,
  -65.9402,
  -66.0079,
  -66.0729,
  -66.1354,
  -66.1958,
  -66.2547,
  -66.3122,
  -66.369,
  -66.4249,
  -66.4802,
  -66.5345,
  -66.5872,
  -66.6381,
  -66.6875,
  -66.7357,
  -66.7831,
  -66.8304,
  -66.878,
  -66.926,
  -66.9748,
  -67.0237,
  -67.0714,
  -67.1194,
  -67.1669,
  -67.2134,
  -67.2594,
  -67.3048,
  -67.3494,
  -67.3924,
  -67.4341,
  -67.4743,
  -67.5127,
  -67.5492,
  -67.5842,
  -67.6176,
  -67.65,
  -67.6809,
  -67.7105,
  -67.7386,
  -67.7657,
  -67.7915,
  -67.8156,
  -67.8382,
  -67.8575,
  -67.8748,
  -67.8889,
  -67.8992,
  -67.9054,
  -67.907,
  -67.9039,
  -67.8968,
  -67.8854,
  -67.8701,
  -67.8509,
  -67.8281,
  -67.8017,
  -67.7723,
  -67.7409,
  -67.708,
  -67.6743,
  -67.6403,
  -67.606,
  -67.571,
  -67.5353,
  -67.4982,
  -67.46,
  -67.4207,
  -67.3798,
  -67.3358,
  -67.2905,
  -67.2424,
  -67.1915,
  -67.1385,
  -67.0831,
  -67.0251,
  -66.9651,
  -66.9031,
  -66.8403,
  -66.7772,
  -66.7143,
  -66.6519,
  -66.59,
  -66.5286,
  -66.4677,
  -66.4076,
  -66.3488,
  -66.2916,
  -66.2369,
  -66.185,
  -66.1363,
  -66.0906,
  -66.0475,
  -66.0066,
  -65.9674,
  -65.9291,
  -65.8903,
  -65.8528,
  -65.8152,
  -65.7774,
  -65.7387,
  -65.6991,
  -65.6585,
  -65.6169,
  -65.5743,
  -65.5306,
  -65.4857,
  -65.4388,
  -65.3902,
  -65.3399,
  -65.2888,
  -65.2374,
  -65.186,
  -65.1346,
  -65.083,
  -65.0312,
  -64.9791,
  -64.9259,
  -64.8716,
  -64.8159,
  -64.7591,
  -64.7012,
  -64.6421,
  -64.5818,
  -64.5204,
  -64.458,
  -64.3946,
  -64.33,
  -64.2625,
  -64.1934,
  -64.1208,
  -64.0446,
  -63.9648,
  -63.8817,
  -63.7965,
  -63.7098,
  -63.6231,
  -63.5374,
  -63.4532,
  -63.371,
  -63.2905,
  -63.2111,
  -63.132,
  -63.0527,
  -62.973,
  -62.8933,
  -62.8139,
  -62.7344,
  -62.6549,
  -62.5754,
  -62.4957,
  -62.416,
  -62.336,
  -62.2554,
  -62.1736,
  -62.0903,
  -62.0054,
  -61.919,
  -61.8318,
  -61.7444,
  -61.6571,
  -61.571,
  -61.4865,
  -61.4046,
  -61.3261,
  -61.2516,
  -61.1817,
  -61.1164,
  -61.0544,
  -60.9972,
  -60.9435,
  -60.893,
  -60.8456,
  -60.8015,
  -60.76,
  -60.721,
  -60.6837,
  -60.6486,
  -60.6156,
  -60.5854,
  -60.5582,
  -60.5337,
  -60.5115,
  -60.4908,
  -60.4709,
  -60.4518,
  -60.433,
  -60.4147,
  -60.3975,
  -50.7458,
  -50.846,
  -50.9466,
  -51.0489,
  -51.1551,
  -51.2684,
  -51.3903,
  -51.5219,
  -51.6668,
  -51.8247,
  -51.9958,
  -52.1798,
  -52.3751,
  -52.5803,
  -52.793,
  -53.0111,
  -53.2322,
  -53.4562,
  -53.6834,
  -53.914,
  -54.1487,
  -54.3883,
  -54.6319,
  -54.8823,
  -55.1385,
  -55.4008,
  -55.6683,
  -55.9404,
  -56.2168,
  -56.4955,
  -56.7753,
  -57.0542,
  -57.3299,
  -57.5996,
  -57.8606,
  -58.1108,
  -58.3482,
  -58.5711,
  -58.7818,
  -58.9802,
  -59.1678,
  -59.3461,
  -59.5171,
  -59.6822,
  -59.8423,
  -59.9982,
  -60.1495,
  -60.2959,
  -60.4365,
  -60.5713,
  -60.7002,
  -60.8239,
  -60.9428,
  -61.0567,
  -61.168,
  -61.2764,
  -61.3815,
  -61.4831,
  -61.5807,
  -61.6743,
  -61.7635,
  -61.8489,
  -61.9308,
  -62.0106,
  -62.0892,
  -62.1675,
  -62.2462,
  -62.3253,
  -62.405,
  -62.4852,
  -62.5645,
  -62.6444,
  -62.7233,
  -62.8012,
  -62.8781,
  -62.955,
  -63.0323,
  -63.11,
  -63.1884,
  -63.2675,
  -63.3469,
  -63.4264,
  -63.5059,
  -63.5854,
  -63.6649,
  -63.7443,
  -63.8241,
  -63.9042,
  -63.9841,
  -64.0657,
  -64.1485,
  -64.232,
  -64.3162,
  -64.4005,
  -64.4848,
  -64.5693,
  -64.6543,
  -64.7398,
  -64.826,
  -64.9132,
  -65.001,
  -65.0893,
  -65.1778,
  -65.2666,
  -65.3559,
  -65.4451,
  -65.5327,
  -65.6202,
  -65.7062,
  -65.7902,
  -65.8717,
  -65.9504,
  -66.0256,
  -66.0978,
  -66.1665,
  -66.2323,
  -66.2957,
  -66.3565,
  -66.4153,
  -66.4725,
  -66.5288,
  -66.5842,
  -66.6388,
  -66.6927,
  -66.7454,
  -66.7963,
  -66.8449,
  -66.8931,
  -66.9405,
  -66.9872,
  -67.0344,
  -67.0824,
  -67.131,
  -67.1802,
  -67.2295,
  -67.2786,
  -67.3267,
  -67.3742,
  -67.4206,
  -67.4669,
  -67.5121,
  -67.5553,
  -67.5968,
  -67.6363,
  -67.6737,
  -67.7093,
  -67.7431,
  -67.7755,
  -67.8061,
  -67.8363,
  -67.8654,
  -67.8926,
  -67.9182,
  -67.942,
  -67.964,
  -67.9844,
  -68.0025,
  -68.0177,
  -68.0297,
  -68.0381,
  -68.0426,
  -68.0429,
  -68.0386,
  -68.0301,
  -68.0173,
  -68.0009,
  -67.9802,
  -67.9555,
  -67.9273,
  -67.8963,
  -67.8636,
  -67.8299,
  -67.7947,
  -67.76,
  -67.7246,
  -67.6885,
  -67.651,
  -67.6119,
  -67.5717,
  -67.5297,
  -67.4863,
  -67.4408,
  -67.3926,
  -67.3416,
  -67.2881,
  -67.2322,
  -67.1737,
  -67.1123,
  -67.0489,
  -66.9833,
  -66.9168,
  -66.85,
  -66.7831,
  -66.7166,
  -66.651,
  -66.5862,
  -66.5223,
  -66.4596,
  -66.397,
  -66.3371,
  -66.2794,
  -66.2244,
  -66.1724,
  -66.1235,
  -66.0771,
  -66.0333,
  -65.9911,
  -65.9506,
  -65.9111,
  -65.872,
  -65.8332,
  -65.7943,
  -65.7549,
  -65.7146,
  -65.6733,
  -65.6307,
  -65.5871,
  -65.5423,
  -65.496,
  -65.4478,
  -65.398,
  -65.3469,
  -65.2951,
  -65.243,
  -65.191,
  -65.1389,
  -65.0864,
  -65.0335,
  -64.9791,
  -64.9248,
  -64.8697,
  -64.8134,
  -64.756,
  -64.6978,
  -64.6386,
  -64.5785,
  -64.5173,
  -64.4551,
  -64.3919,
  -64.3274,
  -64.2609,
  -64.1917,
  -64.1188,
  -64.0421,
  -63.9614,
  -63.8776,
  -63.7915,
  -63.7038,
  -63.6161,
  -63.5292,
  -63.444,
  -63.3608,
  -63.2789,
  -63.1981,
  -63.1176,
  -63.0371,
  -62.9565,
  -62.8758,
  -62.7949,
  -62.7141,
  -62.6331,
  -62.5522,
  -62.4713,
  -62.3909,
  -62.3104,
  -62.2288,
  -62.1474,
  -62.0644,
  -61.9798,
  -61.8938,
  -61.8068,
  -61.7193,
  -61.6321,
  -61.5457,
  -61.4609,
  -61.3789,
  -61.3005,
  -61.2266,
  -61.1577,
  -61.0939,
  -61.0348,
  -60.9798,
  -60.9282,
  -60.8797,
  -60.8342,
  -60.7917,
  -60.752,
  -60.7147,
  -60.679,
  -60.6452,
  -60.6137,
  -60.5845,
  -60.5579,
  -60.5339,
  -60.5125,
  -60.4929,
  -60.4748,
  -60.4577,
  -60.4414,
  -60.4257,
  -60.411,
  -50.8043,
  -50.9151,
  -51.0246,
  -51.1371,
  -51.2534,
  -51.3763,
  -51.5085,
  -51.6508,
  -51.8045,
  -51.9695,
  -52.1462,
  -52.3338,
  -52.5314,
  -52.7374,
  -52.9502,
  -53.1678,
  -53.3885,
  -53.6109,
  -53.8377,
  -54.0683,
  -54.3035,
  -54.544,
  -54.7902,
  -55.0425,
  -55.3009,
  -55.5657,
  -55.836,
  -56.1107,
  -56.3893,
  -56.67,
  -56.951,
  -57.2291,
  -57.5038,
  -57.7711,
  -58.0285,
  -58.2743,
  -58.5072,
  -58.7267,
  -58.9336,
  -59.129,
  -59.3142,
  -59.4907,
  -59.6604,
  -59.8246,
  -59.9842,
  -60.1395,
  -60.2902,
  -60.4345,
  -60.5739,
  -60.707,
  -60.8344,
  -60.9562,
  -61.0736,
  -61.1871,
  -61.2974,
  -61.4047,
  -61.5092,
  -61.6102,
  -61.7073,
  -61.7998,
  -61.8881,
  -61.9726,
  -62.0539,
  -62.133,
  -62.2101,
  -62.288,
  -62.3662,
  -62.4451,
  -62.5245,
  -62.6044,
  -62.6843,
  -62.764,
  -62.8432,
  -62.9212,
  -62.9986,
  -63.0762,
  -63.1545,
  -63.2336,
  -63.3138,
  -63.3943,
  -63.4751,
  -63.5547,
  -63.635,
  -63.7152,
  -63.7957,
  -63.8764,
  -63.9575,
  -64.0396,
  -64.1223,
  -64.2057,
  -64.2899,
  -64.3745,
  -64.4592,
  -64.5434,
  -64.627,
  -64.7102,
  -64.7936,
  -64.8776,
  -64.9624,
  -65.0474,
  -65.1345,
  -65.2225,
  -65.3115,
  -65.4006,
  -65.4901,
  -65.5792,
  -65.6679,
  -65.7552,
  -65.8405,
  -65.924,
  -66.0055,
  -66.0841,
  -66.1603,
  -66.233,
  -66.3027,
  -66.3694,
  -66.4335,
  -66.4953,
  -66.5543,
  -66.6104,
  -66.6665,
  -66.722,
  -66.7772,
  -66.8312,
  -66.8845,
  -66.936,
  -66.9859,
  -67.0349,
  -67.0825,
  -67.1297,
  -67.1773,
  -67.2253,
  -67.2744,
  -67.324,
  -67.3736,
  -67.4232,
  -67.4721,
  -67.5206,
  -67.5678,
  -67.614,
  -67.6585,
  -67.7017,
  -67.743,
  -67.7816,
  -67.8178,
  -67.8521,
  -67.8849,
  -67.9168,
  -67.9474,
  -67.977,
  -68.0051,
  -68.0315,
  -68.0561,
  -68.0786,
  -68.0989,
  -68.1171,
  -68.1329,
  -68.1462,
  -68.1558,
  -68.1621,
  -68.1645,
  -68.1631,
  -68.1577,
  -68.1469,
  -68.1328,
  -68.1147,
  -68.0925,
  -68.0667,
  -68.0364,
  -68.0037,
  -67.9696,
  -67.9351,
  -67.9006,
  -67.8651,
  -67.8287,
  -67.7913,
  -67.7523,
  -67.7121,
  -67.6699,
  -67.6263,
  -67.5804,
  -67.5325,
  -67.4822,
  -67.429,
  -67.3731,
  -67.3145,
  -67.2531,
  -67.1889,
  -67.1212,
  -67.0524,
  -66.9823,
  -66.9118,
  -66.8413,
  -66.7712,
  -66.702,
  -66.634,
  -66.5674,
  -66.5022,
  -66.438,
  -66.3757,
  -66.3152,
  -66.2569,
  -66.2015,
  -66.1487,
  -66.0983,
  -66.0504,
  -66.0049,
  -65.9615,
  -65.9198,
  -65.8789,
  -65.8388,
  -65.7989,
  -65.7586,
  -65.7174,
  -65.6747,
  -65.6309,
  -65.5859,
  -65.5384,
  -65.4904,
  -65.4407,
  -65.3898,
  -65.338,
  -65.2858,
  -65.2333,
  -65.1806,
  -65.1276,
  -65.074,
  -65.02,
  -64.9654,
  -64.9099,
  -64.8537,
  -64.7965,
  -64.7388,
  -64.68,
  -64.6207,
  -64.5605,
  -64.4995,
  -64.4377,
  -64.3746,
  -64.3101,
  -64.2433,
  -64.1736,
  -64.1003,
  -64.0229,
  -63.9414,
  -63.8567,
  -63.7698,
  -63.6815,
  -63.5928,
  -63.5051,
  -63.4189,
  -63.3334,
  -63.2504,
  -63.168,
  -63.086,
  -63.0041,
  -62.9222,
  -62.8404,
  -62.7583,
  -62.676,
  -62.5934,
  -62.5112,
  -62.4294,
  -62.348,
  -62.2669,
  -62.1859,
  -62.1043,
  -62.0214,
  -61.937,
  -61.8511,
  -61.7644,
  -61.6775,
  -61.591,
  -61.5052,
  -61.4213,
  -61.3401,
  -61.2627,
  -61.1901,
  -61.1227,
  -61.0606,
  -61.0037,
  -60.951,
  -60.9017,
  -60.8555,
  -60.8122,
  -60.7719,
  -60.7341,
  -60.699,
  -60.665,
  -60.6329,
  -60.6025,
  -60.5737,
  -60.5474,
  -60.5235,
  -60.5011,
  -60.482,
  -60.4651,
  -60.4497,
  -60.4356,
  -60.4222,
  -60.4097,
  -50.832,
  -50.9526,
  -51.0734,
  -51.1955,
  -51.3217,
  -51.454,
  -51.595,
  -51.7463,
  -51.908,
  -52.0799,
  -52.2616,
  -52.4518,
  -52.6517,
  -52.8591,
  -53.0723,
  -53.2901,
  -53.5113,
  -53.7353,
  -53.9631,
  -54.1953,
  -54.4326,
  -54.6758,
  -54.9251,
  -55.1807,
  -55.4428,
  -55.711,
  -55.9834,
  -56.2609,
  -56.5417,
  -56.8238,
  -57.1053,
  -57.3836,
  -57.6562,
  -57.9202,
  -58.1733,
  -58.4142,
  -58.6419,
  -58.8568,
  -59.0597,
  -59.2515,
  -59.4338,
  -59.6072,
  -59.7754,
  -59.9385,
  -60.097,
  -60.2516,
  -60.4017,
  -60.5461,
  -60.6843,
  -60.8163,
  -60.9423,
  -61.0631,
  -61.1794,
  -61.2921,
  -61.4019,
  -61.5089,
  -61.6127,
  -61.7135,
  -61.8087,
  -61.9007,
  -61.9883,
  -62.0719,
  -62.1527,
  -62.2314,
  -62.309,
  -62.3864,
  -62.4644,
  -62.5429,
  -62.6219,
  -62.7013,
  -62.7805,
  -62.8596,
  -62.9382,
  -63.0161,
  -63.0936,
  -63.1707,
  -63.2501,
  -63.3308,
  -63.4127,
  -63.4951,
  -63.5773,
  -63.6593,
  -63.7408,
  -63.822,
  -63.9036,
  -63.9857,
  -64.0688,
  -64.153,
  -64.2378,
  -64.3234,
  -64.4092,
  -64.495,
  -64.5806,
  -64.6639,
  -64.7474,
  -64.8297,
  -64.9121,
  -64.9949,
  -65.0784,
  -65.1633,
  -65.2495,
  -65.3373,
  -65.4265,
  -65.516,
  -65.6056,
  -65.6948,
  -65.7832,
  -65.87,
  -65.9549,
  -66.0378,
  -66.1187,
  -66.1974,
  -66.2723,
  -66.3455,
  -66.4159,
  -66.4839,
  -66.5487,
  -66.6115,
  -66.6712,
  -66.729,
  -66.7854,
  -66.8413,
  -66.8972,
  -66.9521,
  -67.0056,
  -67.0579,
  -67.1089,
  -67.1589,
  -67.2076,
  -67.256,
  -67.3044,
  -67.3533,
  -67.4018,
  -67.4516,
  -67.5018,
  -67.5517,
  -67.6014,
  -67.6504,
  -67.698,
  -67.7447,
  -67.7898,
  -67.8328,
  -67.8735,
  -67.9113,
  -67.9468,
  -67.9805,
  -68.0129,
  -68.0445,
  -68.0744,
  -68.103,
  -68.13,
  -68.1555,
  -68.1789,
  -68.1997,
  -68.2183,
  -68.2335,
  -68.2471,
  -68.258,
  -68.2654,
  -68.2696,
  -68.2701,
  -68.2671,
  -68.2604,
  -68.2493,
  -68.2339,
  -68.2143,
  -68.1905,
  -68.1628,
  -68.1311,
  -68.0969,
  -68.0616,
  -68.0259,
  -67.9902,
  -67.9536,
  -67.9162,
  -67.8777,
  -67.8377,
  -67.7964,
  -67.7533,
  -67.7073,
  -67.6598,
  -67.6102,
  -67.5579,
  -67.5024,
  -67.4446,
  -67.3835,
  -67.3197,
  -67.2528,
  -67.1834,
  -67.1116,
  -67.0385,
  -66.9649,
  -66.8912,
  -66.8178,
  -66.7456,
  -66.675,
  -66.606,
  -66.5386,
  -66.4723,
  -66.4074,
  -66.3441,
  -66.2827,
  -66.2234,
  -66.1661,
  -66.1114,
  -66.0593,
  -66.009,
  -65.9621,
  -65.9172,
  -65.874,
  -65.832,
  -65.7905,
  -65.7489,
  -65.7063,
  -65.6624,
  -65.6167,
  -65.5698,
  -65.5213,
  -65.4713,
  -65.42,
  -65.368,
  -65.3156,
  -65.2631,
  -65.2103,
  -65.1572,
  -65.1033,
  -65.0488,
  -64.9935,
  -64.9374,
  -64.8808,
  -64.8237,
  -64.7659,
  -64.7074,
  -64.6481,
  -64.5883,
  -64.528,
  -64.4669,
  -64.4052,
  -64.3411,
  -64.2761,
  -64.2089,
  -64.1383,
  -64.0643,
  -63.9859,
  -63.9037,
  -63.8182,
  -63.7304,
  -63.6412,
  -63.5517,
  -63.4632,
  -63.376,
  -63.2904,
  -63.2059,
  -63.1217,
  -63.0382,
  -62.9547,
  -62.8714,
  -62.7883,
  -62.705,
  -62.6215,
  -62.538,
  -62.4547,
  -62.3719,
  -62.2896,
  -62.2078,
  -62.126,
  -62.0439,
  -61.9608,
  -61.8764,
  -61.791,
  -61.705,
  -61.6191,
  -61.5339,
  -61.4497,
  -61.3674,
  -61.288,
  -61.2124,
  -61.1407,
  -61.0753,
  -61.0155,
  -60.9608,
  -60.9106,
  -60.864,
  -60.8205,
  -60.7799,
  -60.7418,
  -60.7064,
  -60.6733,
  -60.6414,
  -60.611,
  -60.5818,
  -60.5538,
  -60.5275,
  -60.5031,
  -60.4812,
  -60.4621,
  -60.4457,
  -60.4316,
  -60.419,
  -60.4076,
  -60.397,
  -50.8303,
  -50.9606,
  -51.0908,
  -51.2224,
  -51.3574,
  -51.4977,
  -51.6471,
  -51.8062,
  -51.9747,
  -52.1529,
  -52.3395,
  -52.534,
  -52.7363,
  -52.9452,
  -53.1596,
  -53.3784,
  -53.6012,
  -53.8273,
  -54.0574,
  -54.2928,
  -54.5326,
  -54.7798,
  -55.0336,
  -55.2937,
  -55.5602,
  -55.8325,
  -56.1095,
  -56.39,
  -56.6728,
  -56.9559,
  -57.2372,
  -57.5139,
  -57.7836,
  -58.0436,
  -58.2921,
  -58.5278,
  -58.7494,
  -58.9595,
  -59.1579,
  -59.3461,
  -59.5256,
  -59.6977,
  -59.864,
  -60.0257,
  -60.1833,
  -60.3368,
  -60.4858,
  -60.629,
  -60.7663,
  -60.8973,
  -61.0225,
  -61.1425,
  -61.2572,
  -61.3696,
  -61.4793,
  -61.5863,
  -61.6901,
  -61.7903,
  -61.8863,
  -61.9776,
  -62.0648,
  -62.1481,
  -62.2284,
  -62.3069,
  -62.3844,
  -62.4615,
  -62.5392,
  -62.6172,
  -62.6957,
  -62.7733,
  -62.8517,
  -62.9298,
  -63.0073,
  -63.0848,
  -63.1623,
  -63.2409,
  -63.3213,
  -63.4034,
  -63.4868,
  -63.571,
  -63.6552,
  -63.7385,
  -63.8212,
  -63.9041,
  -63.9875,
  -64.0717,
  -64.1559,
  -64.242,
  -64.3292,
  -64.4169,
  -64.505,
  -64.5925,
  -64.6789,
  -64.764,
  -64.8476,
  -64.9301,
  -65.0118,
  -65.0937,
  -65.1764,
  -65.2605,
  -65.3461,
  -65.4334,
  -65.5219,
  -65.6115,
  -65.7015,
  -65.7898,
  -65.8778,
  -65.9641,
  -66.0484,
  -66.1307,
  -66.2112,
  -66.2893,
  -66.3651,
  -66.4385,
  -66.5098,
  -66.5784,
  -66.6444,
  -66.7076,
  -66.7684,
  -66.827,
  -66.8845,
  -66.9412,
  -66.997,
  -67.0528,
  -67.1077,
  -67.1603,
  -67.2126,
  -67.2635,
  -67.314,
  -67.3638,
  -67.4136,
  -67.4636,
  -67.5138,
  -67.5641,
  -67.6145,
  -67.665,
  -67.715,
  -67.7642,
  -67.8125,
  -67.8595,
  -67.9048,
  -67.9477,
  -67.9878,
  -68.0255,
  -68.0609,
  -68.0949,
  -68.1261,
  -68.1565,
  -68.1859,
  -68.2136,
  -68.2397,
  -68.2637,
  -68.2852,
  -68.3044,
  -68.3209,
  -68.3352,
  -68.3463,
  -68.3546,
  -68.3598,
  -68.3617,
  -68.3605,
  -68.3558,
  -68.3472,
  -68.3348,
  -68.3182,
  -68.2977,
  -68.2726,
  -68.2432,
  -68.2105,
  -68.1752,
  -68.1378,
  -68.1009,
  -68.0636,
  -68.0257,
  -67.9871,
  -67.9474,
  -67.9066,
  -67.8644,
  -67.8205,
  -67.7747,
  -67.7266,
  -67.6758,
  -67.6218,
  -67.5648,
  -67.5049,
  -67.4416,
  -67.3749,
  -67.3056,
  -67.2335,
  -67.1593,
  -67.0839,
  -67.0078,
  -66.9314,
  -66.8559,
  -66.7816,
  -66.7091,
  -66.6373,
  -66.568,
  -66.5,
  -66.4328,
  -66.3667,
  -66.3018,
  -66.2383,
  -66.177,
  -66.1178,
  -66.061,
  -66.0072,
  -65.9561,
  -65.9074,
  -65.8608,
  -65.8159,
  -65.772,
  -65.7281,
  -65.6834,
  -65.6374,
  -65.5898,
  -65.5406,
  -65.4897,
  -65.4379,
  -65.3851,
  -65.332,
  -65.279,
  -65.226,
  -65.173,
  -65.1196,
  -65.0653,
  -65.009,
  -64.9526,
  -64.8956,
  -64.8376,
  -64.7793,
  -64.7207,
  -64.6614,
  -64.6018,
  -64.5415,
  -64.4809,
  -64.4195,
  -64.3572,
  -64.2936,
  -64.228,
  -64.1595,
  -64.0879,
  -64.0125,
  -63.9331,
  -63.8498,
  -63.7634,
  -63.6747,
  -63.5847,
  -63.4943,
  -63.4048,
  -63.3165,
  -63.2294,
  -63.143,
  -63.0573,
  -62.9719,
  -62.887,
  -62.8025,
  -62.7178,
  -62.6337,
  -62.5494,
  -62.4653,
  -62.3814,
  -62.2969,
  -62.214,
  -62.1313,
  -62.0488,
  -61.966,
  -61.8825,
  -61.7984,
  -61.7135,
  -61.6287,
  -61.5444,
  -61.4609,
  -61.3789,
  -61.299,
  -61.2221,
  -61.1491,
  -61.0808,
  -61.0179,
  -60.9605,
  -60.9085,
  -60.8611,
  -60.8173,
  -60.7767,
  -60.739,
  -60.7039,
  -60.6711,
  -60.6403,
  -60.6106,
  -60.582,
  -60.5539,
  -60.5265,
  -60.5001,
  -60.4753,
  -60.4531,
  -60.4336,
  -60.4174,
  -60.4039,
  -60.3924,
  -60.3824,
  -60.3734,
  -50.7973,
  -50.9365,
  -51.0756,
  -51.2159,
  -51.3594,
  -51.5088,
  -51.6658,
  -51.8316,
  -52.0065,
  -52.1899,
  -52.3811,
  -52.5791,
  -52.7839,
  -52.9945,
  -53.2107,
  -53.4306,
  -53.6558,
  -53.885,
  -54.1191,
  -54.3588,
  -54.6044,
  -54.8567,
  -55.1158,
  -55.3812,
  -55.6526,
  -55.9293,
  -56.2101,
  -56.4938,
  -56.7784,
  -57.0623,
  -57.3419,
  -57.6167,
  -57.8832,
  -58.139,
  -58.3827,
  -58.6132,
  -58.8308,
  -59.0362,
  -59.2302,
  -59.4148,
  -59.5914,
  -59.7613,
  -59.9259,
  -60.0861,
  -60.2424,
  -60.3946,
  -60.541,
  -60.6831,
  -60.8192,
  -60.9495,
  -61.0738,
  -61.1934,
  -61.3089,
  -61.4212,
  -61.531,
  -61.6382,
  -61.742,
  -61.8421,
  -61.9378,
  -62.029,
  -62.116,
  -62.1992,
  -62.2787,
  -62.3573,
  -62.4348,
  -62.5119,
  -62.5892,
  -62.6668,
  -62.7446,
  -62.8221,
  -62.8995,
  -62.9762,
  -63.0529,
  -63.1298,
  -63.2072,
  -63.2862,
  -63.3673,
  -63.4507,
  -63.5358,
  -63.6218,
  -63.7068,
  -63.7919,
  -63.8766,
  -63.9614,
  -64.0466,
  -64.1329,
  -64.2202,
  -64.3089,
  -64.3986,
  -64.4888,
  -64.5791,
  -64.6684,
  -64.7561,
  -64.8424,
  -64.927,
  -65.0099,
  -65.0918,
  -65.1733,
  -65.2545,
  -65.3377,
  -65.4227,
  -65.5094,
  -65.5976,
  -65.6869,
  -65.7765,
  -65.8656,
  -65.9535,
  -66.0392,
  -66.1229,
  -66.2044,
  -66.2845,
  -66.3622,
  -66.4379,
  -66.5117,
  -66.5837,
  -66.6533,
  -66.7201,
  -66.7841,
  -66.8446,
  -66.904,
  -66.9621,
  -67.0195,
  -67.0765,
  -67.1333,
  -67.1892,
  -67.2441,
  -67.2978,
  -67.3503,
  -67.4027,
  -67.4542,
  -67.5054,
  -67.5565,
  -67.6074,
  -67.6588,
  -67.7101,
  -67.7611,
  -67.8114,
  -67.8612,
  -67.9102,
  -67.9565,
  -68.002,
  -68.0449,
  -68.0852,
  -68.1232,
  -68.1592,
  -68.1932,
  -68.2253,
  -68.2555,
  -68.2842,
  -68.3108,
  -68.3354,
  -68.3575,
  -68.3771,
  -68.3943,
  -68.4087,
  -68.4204,
  -68.4292,
  -68.4349,
  -68.4379,
  -68.4377,
  -68.4344,
  -68.4264,
  -68.416,
  -68.4024,
  -68.3846,
  -68.3628,
  -68.3367,
  -68.3066,
  -68.2732,
  -68.2374,
  -68.2003,
  -68.1625,
  -68.124,
  -68.085,
  -68.0451,
  -68.0043,
  -67.9623,
  -67.9189,
  -67.8744,
  -67.8281,
  -67.7793,
  -67.7276,
  -67.6726,
  -67.6145,
  -67.553,
  -67.4879,
  -67.4178,
  -67.3459,
  -67.2715,
  -67.1951,
  -67.1177,
  -67.0396,
  -66.9614,
  -66.8842,
  -66.8086,
  -66.735,
  -66.6631,
  -66.5926,
  -66.5232,
  -66.4541,
  -66.3852,
  -66.3168,
  -66.2497,
  -66.1842,
  -66.1206,
  -66.0592,
  -66.0003,
  -65.944,
  -65.8907,
  -65.84,
  -65.7913,
  -65.7436,
  -65.6962,
  -65.6484,
  -65.5994,
  -65.5477,
  -65.4957,
  -65.4425,
  -65.389,
  -65.3349,
  -65.2809,
  -65.2271,
  -65.1738,
  -65.1205,
  -65.0667,
  -65.012,
  -64.9563,
  -64.8991,
  -64.8411,
  -64.7823,
  -64.723,
  -64.6634,
  -64.6034,
  -64.5434,
  -64.4826,
  -64.4213,
  -64.3592,
  -64.2961,
  -64.2314,
  -64.1645,
  -64.0946,
  -64.0211,
  -63.9439,
  -63.8629,
  -63.7785,
  -63.6909,
  -63.6011,
  -63.51,
  -63.4174,
  -63.3266,
  -63.2368,
  -63.148,
  -63.0599,
  -62.9726,
  -62.8857,
  -62.7993,
  -62.7134,
  -62.6281,
  -62.5432,
  -62.4587,
  -62.3745,
  -62.2903,
  -62.2065,
  -62.1232,
  -62.0402,
  -61.9572,
  -61.8738,
  -61.7903,
  -61.7065,
  -61.6227,
  -61.5393,
  -61.4567,
  -61.3755,
  -61.2961,
  -61.219,
  -61.145,
  -61.0749,
  -61.0096,
  -60.9494,
  -60.8948,
  -60.8456,
  -60.8011,
  -60.7604,
  -60.7231,
  -60.6885,
  -60.6565,
  -60.6267,
  -60.5984,
  -60.5712,
  -60.5443,
  -60.5166,
  -60.4899,
  -60.4637,
  -60.4387,
  -60.4159,
  -60.3965,
  -60.3803,
  -60.3671,
  -60.3561,
  -60.347,
  -60.3394,
  -50.7348,
  -50.8826,
  -51.0296,
  -51.1777,
  -51.3292,
  -51.486,
  -51.6501,
  -51.8222,
  -52.0028,
  -52.1911,
  -52.3858,
  -52.5872,
  -52.7946,
  -53.0075,
  -53.2261,
  -53.4496,
  -53.6779,
  -53.9112,
  -54.1501,
  -54.3948,
  -54.646,
  -54.9042,
  -55.1692,
  -55.4403,
  -55.7171,
  -55.9974,
  -56.2822,
  -56.569,
  -56.8557,
  -57.1401,
  -57.4199,
  -57.6927,
  -57.9559,
  -58.2077,
  -58.447,
  -58.6726,
  -58.8853,
  -59.086,
  -59.276,
  -59.4571,
  -59.6298,
  -59.7975,
  -59.9602,
  -60.1189,
  -60.2736,
  -60.4243,
  -60.5702,
  -60.7109,
  -60.8459,
  -60.975,
  -61.0989,
  -61.2181,
  -61.3336,
  -61.4461,
  -61.556,
  -61.6633,
  -61.7662,
  -61.8664,
  -61.9619,
  -62.0529,
  -62.1399,
  -62.2235,
  -62.3043,
  -62.3832,
  -62.461,
  -62.5386,
  -62.616,
  -62.6933,
  -62.7705,
  -62.847,
  -62.9231,
  -62.9988,
  -63.0745,
  -63.1499,
  -63.2272,
  -63.3067,
  -63.3887,
  -63.4731,
  -63.5596,
  -63.6472,
  -63.735,
  -63.8221,
  -63.9089,
  -63.9955,
  -64.0828,
  -64.1715,
  -64.2617,
  -64.3527,
  -64.4449,
  -64.5375,
  -64.6299,
  -64.7204,
  -64.8102,
  -64.8981,
  -64.9839,
  -65.068,
  -65.1506,
  -65.2322,
  -65.314,
  -65.3967,
  -65.4809,
  -65.5671,
  -65.6547,
  -65.7436,
  -65.8326,
  -65.9211,
  -66.0084,
  -66.0938,
  -66.1768,
  -66.258,
  -66.3375,
  -66.4144,
  -66.4903,
  -66.5647,
  -66.6374,
  -66.7076,
  -66.7752,
  -66.8399,
  -66.902,
  -66.9621,
  -67.021,
  -67.0791,
  -67.1368,
  -67.1941,
  -67.2506,
  -67.3067,
  -67.3621,
  -67.4164,
  -67.4703,
  -67.5237,
  -67.5767,
  -67.6286,
  -67.6811,
  -67.7333,
  -67.7856,
  -67.8374,
  -67.8884,
  -67.9386,
  -67.9882,
  -68.0359,
  -68.0817,
  -68.1254,
  -68.1665,
  -68.2053,
  -68.2418,
  -68.2762,
  -68.3088,
  -68.3389,
  -68.3668,
  -68.3921,
  -68.415,
  -68.4351,
  -68.4526,
  -68.4667,
  -68.4788,
  -68.4883,
  -68.4947,
  -68.4981,
  -68.4987,
  -68.4962,
  -68.4906,
  -68.4817,
  -68.4693,
  -68.4537,
  -68.4345,
  -68.4116,
  -68.3849,
  -68.3542,
  -68.3204,
  -68.2841,
  -68.2468,
  -68.2087,
  -68.1698,
  -68.1298,
  -68.0889,
  -68.0472,
  -68.0044,
  -67.9593,
  -67.9138,
  -67.8666,
  -67.8169,
  -67.7646,
  -67.7091,
  -67.6502,
  -67.5874,
  -67.5209,
  -67.4508,
  -67.3773,
  -67.301,
  -67.2225,
  -67.143,
  -67.0632,
  -66.9838,
  -66.9057,
  -66.8293,
  -66.7548,
  -66.6823,
  -66.6109,
  -66.5402,
  -66.4692,
  -66.3983,
  -66.3275,
  -66.2569,
  -66.1874,
  -66.1182,
  -66.052,
  -65.9882,
  -65.9269,
  -65.8683,
  -65.8122,
  -65.7582,
  -65.7057,
  -65.6537,
  -65.601,
  -65.5478,
  -65.4935,
  -65.4383,
  -65.3825,
  -65.3268,
  -65.2712,
  -65.2165,
  -65.1623,
  -65.1084,
  -65.0547,
  -65.0004,
  -64.9453,
  -64.8889,
  -64.8312,
  -64.7724,
  -64.7129,
  -64.653,
  -64.5927,
  -64.532,
  -64.4712,
  -64.41,
  -64.3471,
  -64.2842,
  -64.2198,
  -64.1537,
  -64.0849,
  -64.0129,
  -63.9373,
  -63.8579,
  -63.7747,
  -63.688,
  -63.5989,
  -63.5078,
  -63.4151,
  -63.3221,
  -63.2297,
  -63.1382,
  -63.0477,
  -62.9578,
  -62.8688,
  -62.7803,
  -62.6928,
  -62.6063,
  -62.5206,
  -62.4358,
  -62.3514,
  -62.2675,
  -62.1838,
  -62.1003,
  -62.0169,
  -61.9337,
  -61.8506,
  -61.7675,
  -61.6842,
  -61.6011,
  -61.5185,
  -61.4369,
  -61.3565,
  -61.2777,
  -61.2011,
  -61.126,
  -61.0553,
  -60.9884,
  -60.926,
  -60.8688,
  -60.8171,
  -60.7707,
  -60.7291,
  -60.6915,
  -60.6573,
  -60.6261,
  -60.5975,
  -60.5709,
  -60.5455,
  -60.5208,
  -60.496,
  -60.4707,
  -60.445,
  -60.4192,
  -60.3943,
  -60.3715,
  -60.3519,
  -60.3357,
  -60.3226,
  -60.3119,
  -60.3032,
  -60.2964,
  -50.6422,
  -50.7981,
  -50.9526,
  -51.1081,
  -51.2658,
  -51.4295,
  -51.6001,
  -51.7783,
  -51.9641,
  -52.1572,
  -52.3567,
  -52.5621,
  -52.7724,
  -52.9881,
  -53.2095,
  -53.4362,
  -53.6684,
  -53.9061,
  -54.15,
  -54.3995,
  -54.6566,
  -54.9209,
  -55.192,
  -55.4689,
  -55.7512,
  -56.0375,
  -56.3266,
  -56.6164,
  -56.9051,
  -57.1904,
  -57.4695,
  -57.7403,
  -58.0006,
  -58.2488,
  -58.4838,
  -58.7042,
  -58.9125,
  -59.1088,
  -59.2949,
  -59.4726,
  -59.6436,
  -59.8092,
  -59.9701,
  -60.1274,
  -60.2805,
  -60.4295,
  -60.5737,
  -60.7128,
  -60.8464,
  -60.9746,
  -61.0978,
  -61.2158,
  -61.3312,
  -61.4438,
  -61.5537,
  -61.661,
  -61.765,
  -61.8648,
  -61.9603,
  -62.0512,
  -62.1383,
  -62.2223,
  -62.3037,
  -62.3834,
  -62.4621,
  -62.5403,
  -62.6182,
  -62.6943,
  -62.7711,
  -62.8469,
  -62.9222,
  -62.9971,
  -63.0723,
  -63.1483,
  -63.2258,
  -63.3056,
  -63.3886,
  -63.4741,
  -63.5618,
  -63.6506,
  -63.74,
  -63.8293,
  -63.9179,
  -64.0069,
  -64.0967,
  -64.1869,
  -64.2796,
  -64.3734,
  -64.4681,
  -64.5631,
  -64.6579,
  -64.7518,
  -64.8436,
  -64.9332,
  -65.0204,
  -65.106,
  -65.1897,
  -65.272,
  -65.3538,
  -65.4364,
  -65.5202,
  -65.6055,
  -65.6919,
  -65.7798,
  -65.867,
  -65.9547,
  -66.0413,
  -66.1263,
  -66.2094,
  -66.2906,
  -66.3706,
  -66.4491,
  -66.5259,
  -66.6009,
  -66.6739,
  -66.7447,
  -66.8127,
  -66.8775,
  -66.9399,
  -67.0003,
  -67.0595,
  -67.1182,
  -67.1758,
  -67.2324,
  -67.2896,
  -67.3466,
  -67.4034,
  -67.4595,
  -67.5154,
  -67.5709,
  -67.6262,
  -67.6811,
  -67.7352,
  -67.7886,
  -67.8415,
  -67.8943,
  -67.9462,
  -67.9972,
  -68.0469,
  -68.0953,
  -68.1423,
  -68.1873,
  -68.2293,
  -68.2689,
  -68.3063,
  -68.3405,
  -68.3735,
  -68.4033,
  -68.4304,
  -68.4544,
  -68.4757,
  -68.4944,
  -68.5099,
  -68.5227,
  -68.5328,
  -68.5399,
  -68.5443,
  -68.5453,
  -68.5437,
  -68.5392,
  -68.5314,
  -68.5206,
  -68.5063,
  -68.4886,
  -68.4678,
  -68.4439,
  -68.4163,
  -68.3849,
  -68.3498,
  -68.3134,
  -68.2761,
  -68.2381,
  -68.1988,
  -68.1584,
  -68.117,
  -68.0748,
  -68.0316,
  -67.9866,
  -67.9403,
  -67.8922,
  -67.8418,
  -67.7889,
  -67.7325,
  -67.673,
  -67.6098,
  -67.5429,
  -67.4723,
  -67.3978,
  -67.3205,
  -67.2409,
  -67.1599,
  -67.0788,
  -66.9983,
  -66.9194,
  -66.8413,
  -66.7664,
  -66.6933,
  -66.6209,
  -66.549,
  -66.4771,
  -66.4047,
  -66.3319,
  -66.2587,
  -66.1857,
  -66.1133,
  -66.0422,
  -65.9733,
  -65.9068,
  -65.8425,
  -65.7807,
  -65.7208,
  -65.6621,
  -65.604,
  -65.5458,
  -65.4869,
  -65.4278,
  -65.3684,
  -65.3098,
  -65.2516,
  -65.1944,
  -65.1384,
  -65.0833,
  -65.0286,
  -64.9742,
  -64.9183,
  -64.8626,
  -64.8058,
  -64.7475,
  -64.688,
  -64.6278,
  -64.5672,
  -64.5064,
  -64.4452,
  -64.3838,
  -64.322,
  -64.2594,
  -64.1955,
  -64.1296,
  -64.0614,
  -63.9903,
  -63.9158,
  -63.8374,
  -63.755,
  -63.6692,
  -63.5802,
  -63.4887,
  -63.3955,
  -63.3011,
  -63.2065,
  -63.1122,
  -63.0188,
  -62.9265,
  -62.835,
  -62.7443,
  -62.6548,
  -62.5666,
  -62.4799,
  -62.3945,
  -62.3102,
  -62.2257,
  -62.1429,
  -62.0602,
  -61.9774,
  -61.8947,
  -61.812,
  -61.7293,
  -61.6468,
  -61.5644,
  -61.4825,
  -61.4014,
  -61.3217,
  -61.2435,
  -61.1673,
  -61.0934,
  -61.0224,
  -60.9548,
  -60.8911,
  -60.8321,
  -60.7779,
  -60.7289,
  -60.6853,
  -60.6466,
  -60.6119,
  -60.5808,
  -60.5529,
  -60.5277,
  -60.5045,
  -60.4823,
  -60.4603,
  -60.4378,
  -60.4144,
  -60.39,
  -60.3648,
  -60.3404,
  -60.3179,
  -60.2983,
  -60.2821,
  -60.2688,
  -60.2583,
  -60.25,
  -60.244,
  -50.5204,
  -50.6833,
  -50.8451,
  -51.0073,
  -51.1724,
  -51.3429,
  -51.5196,
  -51.7036,
  -51.8947,
  -52.0924,
  -52.296,
  -52.5051,
  -52.7191,
  -52.9381,
  -53.1616,
  -53.3919,
  -53.6282,
  -53.8709,
  -54.12,
  -54.3763,
  -54.6393,
  -54.9097,
  -55.1867,
  -55.4696,
  -55.7574,
  -56.0489,
  -56.3423,
  -56.6353,
  -56.9261,
  -57.2112,
  -57.4898,
  -57.759,
  -58.0171,
  -58.2621,
  -58.4935,
  -58.7112,
  -58.9156,
  -59.1081,
  -59.2907,
  -59.4653,
  -59.6335,
  -59.7969,
  -59.9562,
  -60.1118,
  -60.2634,
  -60.4096,
  -60.5523,
  -60.6898,
  -60.822,
  -60.9491,
  -61.0713,
  -61.1897,
  -61.3047,
  -61.417,
  -61.5267,
  -61.6337,
  -61.7374,
  -61.8369,
  -61.9321,
  -62.0231,
  -62.1102,
  -62.1937,
  -62.276,
  -62.357,
  -62.4369,
  -62.5159,
  -62.5942,
  -62.6717,
  -62.7482,
  -62.8238,
  -62.8988,
  -62.9733,
  -63.0484,
  -63.1246,
  -63.2027,
  -63.2835,
  -63.3671,
  -63.4535,
  -63.5422,
  -63.6313,
  -63.7222,
  -63.8132,
  -63.9042,
  -63.9956,
  -64.0879,
  -64.1818,
  -64.2772,
  -64.3737,
  -64.4711,
  -64.5689,
  -64.6661,
  -64.7619,
  -64.8558,
  -64.9476,
  -65.0367,
  -65.1235,
  -65.2085,
  -65.2909,
  -65.3732,
  -65.4553,
  -65.5383,
  -65.6226,
  -65.7082,
  -65.7948,
  -65.8818,
  -65.9689,
  -66.0549,
  -66.14,
  -66.2234,
  -66.3055,
  -66.3862,
  -66.4654,
  -66.5431,
  -66.6188,
  -66.6923,
  -66.763,
  -66.8296,
  -66.8943,
  -66.9564,
  -67.0169,
  -67.076,
  -67.1342,
  -67.192,
  -67.2498,
  -67.3076,
  -67.3654,
  -67.4236,
  -67.4818,
  -67.5398,
  -67.598,
  -67.6556,
  -67.7124,
  -67.7681,
  -67.8229,
  -67.8771,
  -67.9304,
  -67.983,
  -68.0339,
  -68.0849,
  -68.1348,
  -68.1827,
  -68.2285,
  -68.2716,
  -68.3126,
  -68.3514,
  -68.3872,
  -68.4201,
  -68.4496,
  -68.4758,
  -68.4989,
  -68.5189,
  -68.536,
  -68.5499,
  -68.5608,
  -68.569,
  -68.5739,
  -68.5761,
  -68.5751,
  -68.5715,
  -68.5649,
  -68.5542,
  -68.5413,
  -68.5251,
  -68.5058,
  -68.4834,
  -68.4581,
  -68.4295,
  -68.3977,
  -68.3635,
  -68.3274,
  -68.2898,
  -68.2517,
  -68.2125,
  -68.1723,
  -68.1312,
  -68.0888,
  -68.045,
  -67.9995,
  -67.9524,
  -67.9036,
  -67.8526,
  -67.799,
  -67.7423,
  -67.6824,
  -67.6181,
  -67.5509,
  -67.4801,
  -67.4058,
  -67.3284,
  -67.2485,
  -67.1671,
  -67.0855,
  -67.0044,
  -66.9248,
  -66.8471,
  -66.7715,
  -66.6975,
  -66.6241,
  -66.5514,
  -66.4786,
  -66.4052,
  -66.3311,
  -66.2559,
  -66.1802,
  -66.1044,
  -66.0292,
  -65.9552,
  -65.8829,
  -65.8127,
  -65.7447,
  -65.6782,
  -65.6128,
  -65.5469,
  -65.4818,
  -65.4165,
  -65.3515,
  -65.2875,
  -65.225,
  -65.1639,
  -65.1047,
  -65.0468,
  -64.9901,
  -64.934,
  -64.8782,
  -64.8223,
  -64.7659,
  -64.7083,
  -64.6494,
  -64.5893,
  -64.5283,
  -64.4668,
  -64.4052,
  -64.3436,
  -64.2818,
  -64.2195,
  -64.156,
  -64.0908,
  -64.0232,
  -63.9527,
  -63.8788,
  -63.8012,
  -63.7194,
  -63.6338,
  -63.5446,
  -63.4527,
  -63.3573,
  -63.2617,
  -63.1654,
  -63.0687,
  -62.9726,
  -62.8772,
  -62.783,
  -62.6901,
  -62.5984,
  -62.5082,
  -62.4198,
  -62.3333,
  -62.2486,
  -62.1657,
  -62.0839,
  -62.0027,
  -61.9218,
  -61.8405,
  -61.7591,
  -61.6777,
  -61.596,
  -61.5146,
  -61.4335,
  -61.3532,
  -61.2741,
  -61.1963,
  -61.1202,
  -61.0463,
  -60.9751,
  -60.9071,
  -60.8427,
  -60.7824,
  -60.7265,
  -60.6755,
  -60.6295,
  -60.5885,
  -60.5523,
  -60.5202,
  -60.4921,
  -60.4675,
  -60.4457,
  -60.4259,
  -60.4061,
  -60.3871,
  -60.367,
  -60.3454,
  -60.3223,
  -60.2983,
  -60.2744,
  -60.2524,
  -60.233,
  -60.2166,
  -60.2032,
  -60.1927,
  -60.185,
  -60.1799,
  -50.3736,
  -50.5427,
  -50.711,
  -50.8794,
  -51.0506,
  -51.2271,
  -51.4097,
  -51.5992,
  -51.7955,
  -51.997,
  -52.2051,
  -52.4181,
  -52.6364,
  -52.8592,
  -53.0874,
  -53.3216,
  -53.5625,
  -53.8102,
  -54.0645,
  -54.3264,
  -54.5954,
  -54.8718,
  -55.1548,
  -55.4436,
  -55.7361,
  -56.0325,
  -56.3298,
  -56.6258,
  -56.9185,
  -57.2056,
  -57.4841,
  -57.7522,
  -58.0083,
  -58.2509,
  -58.4794,
  -58.6941,
  -58.8954,
  -59.0849,
  -59.2645,
  -59.4352,
  -59.601,
  -59.7623,
  -59.9196,
  -60.0734,
  -60.2233,
  -60.3689,
  -60.5098,
  -60.6458,
  -60.7766,
  -60.9024,
  -61.0236,
  -61.141,
  -61.2552,
  -61.3667,
  -61.4757,
  -61.581,
  -61.6839,
  -61.7831,
  -61.878,
  -61.9689,
  -62.0562,
  -62.141,
  -62.2242,
  -62.3063,
  -62.3871,
  -62.4672,
  -62.5464,
  -62.6244,
  -62.7011,
  -62.7768,
  -62.8519,
  -62.9268,
  -63.0016,
  -63.0786,
  -63.1578,
  -63.2394,
  -63.324,
  -63.4113,
  -63.5008,
  -63.5921,
  -63.6846,
  -63.7775,
  -63.8708,
  -63.9645,
  -64.0595,
  -64.1558,
  -64.2542,
  -64.3539,
  -64.4541,
  -64.5547,
  -64.6534,
  -64.7517,
  -64.8481,
  -64.9417,
  -65.0325,
  -65.121,
  -65.2071,
  -65.2912,
  -65.3738,
  -65.4555,
  -65.5379,
  -65.621,
  -65.7055,
  -65.7911,
  -65.877,
  -65.9633,
  -66.0494,
  -66.1347,
  -66.2189,
  -66.3009,
  -66.3826,
  -66.4629,
  -66.5415,
  -66.6175,
  -66.6908,
  -66.7609,
  -66.828,
  -66.892,
  -66.9535,
  -67.0134,
  -67.0718,
  -67.1297,
  -67.1874,
  -67.2454,
  -67.3035,
  -67.3624,
  -67.422,
  -67.4822,
  -67.5425,
  -67.6019,
  -67.6616,
  -67.7206,
  -67.7785,
  -67.8347,
  -67.89,
  -67.9446,
  -67.9987,
  -68.0523,
  -68.1048,
  -68.1557,
  -68.2047,
  -68.2519,
  -68.2967,
  -68.3387,
  -68.3782,
  -68.4143,
  -68.4471,
  -68.4764,
  -68.502,
  -68.5242,
  -68.543,
  -68.5578,
  -68.5705,
  -68.5797,
  -68.5859,
  -68.589,
  -68.5892,
  -68.5865,
  -68.5806,
  -68.5719,
  -68.5602,
  -68.5457,
  -68.5281,
  -68.5072,
  -68.4833,
  -68.4564,
  -68.4271,
  -68.3951,
  -68.3609,
  -68.3247,
  -68.2873,
  -68.2493,
  -68.2102,
  -68.1704,
  -68.1293,
  -68.086,
  -68.0424,
  -67.9971,
  -67.9499,
  -67.9004,
  -67.8484,
  -67.7941,
  -67.7374,
  -67.6775,
  -67.6143,
  -67.5471,
  -67.4767,
  -67.403,
  -67.326,
  -67.2467,
  -67.166,
  -67.0847,
  -67.0039,
  -66.9243,
  -66.8464,
  -66.7699,
  -66.6946,
  -66.6203,
  -66.5464,
  -66.4727,
  -66.3982,
  -66.3227,
  -66.245,
  -66.1671,
  -66.0884,
  -66.0098,
  -65.9316,
  -65.8543,
  -65.7783,
  -65.7037,
  -65.6303,
  -65.5576,
  -65.4853,
  -65.413,
  -65.3408,
  -65.2695,
  -65.2,
  -65.1326,
  -65.0677,
  -65.0053,
  -64.9447,
  -64.8856,
  -64.8275,
  -64.7697,
  -64.712,
  -64.6539,
  -64.5951,
  -64.5351,
  -64.4741,
  -64.412,
  -64.3495,
  -64.2872,
  -64.2252,
  -64.1618,
  -64.099,
  -64.0345,
  -63.9678,
  -63.8979,
  -63.8248,
  -63.7477,
  -63.6665,
  -63.5811,
  -63.4917,
  -63.399,
  -63.3037,
  -63.2065,
  -63.1085,
  -63.0099,
  -62.9115,
  -62.8132,
  -62.7162,
  -62.6205,
  -62.5265,
  -62.434,
  -62.3434,
  -62.2551,
  -62.1693,
  -62.0861,
  -62.0048,
  -61.9252,
  -61.8464,
  -61.7678,
  -61.6891,
  -61.6099,
  -61.5302,
  -61.4503,
  -61.3705,
  -61.2912,
  -61.2126,
  -61.1352,
  -61.0594,
  -60.9848,
  -60.9135,
  -60.8451,
  -60.7801,
  -60.7189,
  -60.6619,
  -60.6093,
  -60.5614,
  -60.5182,
  -60.4797,
  -60.4458,
  -60.4162,
  -60.3909,
  -60.3692,
  -60.3505,
  -60.3338,
  -60.3178,
  -60.3016,
  -60.2839,
  -60.2641,
  -60.2425,
  -60.2198,
  -60.1969,
  -60.1752,
  -60.156,
  -60.1397,
  -60.1263,
  -60.1159,
  -60.1088,
  -60.1049,
  -50.204,
  -50.3787,
  -50.5527,
  -50.7262,
  -50.903,
  -51.085,
  -51.2733,
  -51.468,
  -51.6693,
  -51.8765,
  -52.0893,
  -52.3068,
  -52.5292,
  -52.7566,
  -52.989,
  -53.2276,
  -53.4734,
  -53.7258,
  -53.9844,
  -54.2518,
  -54.5267,
  -54.809,
  -55.098,
  -55.3925,
  -55.6912,
  -55.992,
  -56.2928,
  -56.5916,
  -56.886,
  -57.1741,
  -57.453,
  -57.7205,
  -57.9752,
  -58.2151,
  -58.4416,
  -58.6539,
  -58.8531,
  -59.0404,
  -59.2177,
  -59.3871,
  -59.5507,
  -59.7096,
  -59.8648,
  -60.0165,
  -60.1645,
  -60.3082,
  -60.4476,
  -60.582,
  -60.7115,
  -60.8351,
  -60.955,
  -61.0711,
  -61.1841,
  -61.2942,
  -61.4018,
  -61.5067,
  -61.6085,
  -61.7068,
  -61.8011,
  -61.8917,
  -61.9791,
  -62.0642,
  -62.1481,
  -62.231,
  -62.3127,
  -62.3937,
  -62.4727,
  -62.5515,
  -62.6287,
  -62.7052,
  -62.7813,
  -62.8573,
  -62.9345,
  -63.0129,
  -63.0933,
  -63.176,
  -63.2616,
  -63.3498,
  -63.4402,
  -63.5327,
  -63.6267,
  -63.7215,
  -63.817,
  -63.9133,
  -64.0098,
  -64.1093,
  -64.2108,
  -64.3137,
  -64.417,
  -64.5205,
  -64.6233,
  -64.7243,
  -64.823,
  -64.9189,
  -65.0115,
  -65.1015,
  -65.1885,
  -65.2733,
  -65.3557,
  -65.4372,
  -65.5189,
  -65.6012,
  -65.6833,
  -65.7674,
  -65.8526,
  -65.9383,
  -66.0242,
  -66.1102,
  -66.1953,
  -66.2793,
  -66.3623,
  -66.4434,
  -66.5226,
  -66.5984,
  -66.6712,
  -66.7407,
  -66.8068,
  -66.8697,
  -66.9301,
  -66.9888,
  -67.0466,
  -67.1039,
  -67.1603,
  -67.2178,
  -67.2765,
  -67.3362,
  -67.3971,
  -67.459,
  -67.5212,
  -67.5835,
  -67.6456,
  -67.7067,
  -67.7666,
  -67.8248,
  -67.882,
  -67.9389,
  -67.995,
  -68.0505,
  -68.1043,
  -68.1568,
  -68.2076,
  -68.2563,
  -68.3024,
  -68.344,
  -68.3838,
  -68.4203,
  -68.4532,
  -68.4823,
  -68.5073,
  -68.5288,
  -68.5467,
  -68.5615,
  -68.5729,
  -68.5807,
  -68.5855,
  -68.5872,
  -68.5857,
  -68.5812,
  -68.5733,
  -68.5626,
  -68.5492,
  -68.533,
  -68.5139,
  -68.4915,
  -68.4665,
  -68.4389,
  -68.4079,
  -68.3757,
  -68.3411,
  -68.3051,
  -68.2683,
  -68.2303,
  -68.1914,
  -68.1514,
  -68.1107,
  -68.0689,
  -68.0254,
  -67.9802,
  -67.9326,
  -67.8828,
  -67.8306,
  -67.7761,
  -67.7191,
  -67.6589,
  -67.5959,
  -67.5298,
  -67.4601,
  -67.3874,
  -67.3114,
  -67.2333,
  -67.1539,
  -67.0738,
  -66.993,
  -66.9139,
  -66.8357,
  -66.7587,
  -66.6827,
  -66.6076,
  -66.5326,
  -66.4576,
  -66.3817,
  -66.3049,
  -66.2268,
  -66.1469,
  -66.0661,
  -65.9844,
  -65.9026,
  -65.821,
  -65.7397,
  -65.6589,
  -65.5788,
  -65.4988,
  -65.419,
  -65.3389,
  -65.2593,
  -65.1816,
  -65.1058,
  -65.0328,
  -64.963,
  -64.8963,
  -64.8321,
  -64.7687,
  -64.7077,
  -64.6469,
  -64.5866,
  -64.5261,
  -64.4649,
  -64.4032,
  -64.3403,
  -64.2771,
  -64.2136,
  -64.1503,
  -64.0875,
  -64.0245,
  -63.9605,
  -63.8949,
  -63.8262,
  -63.7541,
  -63.6778,
  -63.5973,
  -63.5125,
  -63.4231,
  -63.3301,
  -63.2336,
  -63.135,
  -63.0349,
  -62.9343,
  -62.8337,
  -62.7333,
  -62.6336,
  -62.5354,
  -62.4386,
  -62.3437,
  -62.2507,
  -62.1602,
  -62.0725,
  -61.9869,
  -61.9053,
  -61.8261,
  -61.749,
  -61.6731,
  -61.5978,
  -61.5223,
  -61.4459,
  -61.3691,
  -61.2917,
  -61.214,
  -61.1367,
  -61.0599,
  -60.9845,
  -60.9109,
  -60.8398,
  -60.7714,
  -60.7059,
  -60.6441,
  -60.5861,
  -60.5325,
  -60.4832,
  -60.4383,
  -60.3978,
  -60.3618,
  -60.3301,
  -60.3029,
  -60.2798,
  -60.2606,
  -60.2446,
  -60.2303,
  -60.2165,
  -60.202,
  -60.186,
  -60.1682,
  -60.1481,
  -60.1264,
  -60.1044,
  -60.0835,
  -60.0647,
  -60.0485,
  -60.0354,
  -60.0257,
  -60.0196,
  -60.0173,
  -50.0135,
  -50.1939,
  -50.373,
  -50.5528,
  -50.7353,
  -50.9221,
  -51.1155,
  -51.3154,
  -51.5214,
  -51.7336,
  -51.951,
  -52.1732,
  -52.4,
  -52.6312,
  -52.8687,
  -53.1121,
  -53.3625,
  -53.6203,
  -53.8852,
  -54.1578,
  -54.4381,
  -54.7259,
  -55.0203,
  -55.3201,
  -55.6236,
  -55.9285,
  -56.2325,
  -56.5336,
  -56.8287,
  -57.1179,
  -57.3974,
  -57.6649,
  -57.919,
  -58.1589,
  -58.384,
  -58.595,
  -58.7926,
  -58.9783,
  -59.1539,
  -59.3216,
  -59.4832,
  -59.64,
  -59.793,
  -59.9425,
  -60.0875,
  -60.2293,
  -60.3669,
  -60.4998,
  -60.6279,
  -60.7512,
  -60.8698,
  -60.9845,
  -61.0956,
  -61.2037,
  -61.3094,
  -61.4122,
  -61.5123,
  -61.6091,
  -61.7025,
  -61.7923,
  -61.8782,
  -61.9634,
  -62.0475,
  -62.1309,
  -62.2135,
  -62.295,
  -62.3756,
  -62.4553,
  -62.5337,
  -62.6116,
  -62.6893,
  -62.7674,
  -62.8464,
  -62.9266,
  -63.0085,
  -63.0924,
  -63.1788,
  -63.2671,
  -63.3587,
  -63.4524,
  -63.5478,
  -63.6445,
  -63.7423,
  -63.8413,
  -63.9419,
  -64.0445,
  -64.1495,
  -64.2558,
  -64.3626,
  -64.4694,
  -64.5751,
  -64.6792,
  -64.7805,
  -64.8788,
  -64.9735,
  -65.0647,
  -65.1515,
  -65.2369,
  -65.3202,
  -65.4016,
  -65.4821,
  -65.563,
  -65.6448,
  -65.7276,
  -65.8116,
  -65.8967,
  -65.9827,
  -66.0692,
  -66.1553,
  -66.2406,
  -66.3245,
  -66.4063,
  -66.4856,
  -66.5611,
  -66.6332,
  -66.7002,
  -66.7649,
  -66.8264,
  -66.8854,
  -66.9431,
  -66.9998,
  -67.0563,
  -67.1132,
  -67.1707,
  -67.2295,
  -67.2894,
  -67.3511,
  -67.4141,
  -67.4776,
  -67.5417,
  -67.6056,
  -67.669,
  -67.731,
  -67.792,
  -67.8522,
  -67.9116,
  -67.9689,
  -68.0264,
  -68.0825,
  -68.1369,
  -68.1893,
  -68.2391,
  -68.286,
  -68.3298,
  -68.3704,
  -68.4072,
  -68.4402,
  -68.4691,
  -68.4936,
  -68.5143,
  -68.5314,
  -68.5453,
  -68.5557,
  -68.5628,
  -68.5664,
  -68.5667,
  -68.5639,
  -68.5579,
  -68.5475,
  -68.5353,
  -68.52,
  -68.502,
  -68.4812,
  -68.4577,
  -68.4316,
  -68.4031,
  -68.3729,
  -68.3406,
  -68.3064,
  -68.2705,
  -68.2334,
  -68.1955,
  -68.1572,
  -68.1175,
  -68.0768,
  -68.0349,
  -67.9914,
  -67.9462,
  -67.8987,
  -67.8488,
  -67.7965,
  -67.742,
  -67.6852,
  -67.6245,
  -67.5622,
  -67.4967,
  -67.4282,
  -67.3569,
  -67.2828,
  -67.2066,
  -67.1287,
  -67.05,
  -66.9713,
  -66.893,
  -66.8152,
  -66.738,
  -66.6616,
  -66.5853,
  -66.5092,
  -66.4331,
  -66.3562,
  -66.2781,
  -66.1985,
  -66.117,
  -66.034,
  -65.9501,
  -65.8652,
  -65.78,
  -65.6942,
  -65.6081,
  -65.5202,
  -65.4331,
  -65.3457,
  -65.258,
  -65.1713,
  -65.0865,
  -65.004,
  -64.925,
  -64.8495,
  -64.7777,
  -64.7089,
  -64.6422,
  -64.5769,
  -64.5124,
  -64.4483,
  -64.3843,
  -64.3199,
  -64.2552,
  -64.1901,
  -64.1249,
  -64.0598,
  -63.9955,
  -63.9314,
  -63.8672,
  -63.8019,
  -63.7344,
  -63.6638,
  -63.589,
  -63.5096,
  -63.4256,
  -63.3368,
  -63.2436,
  -63.1468,
  -63.0458,
  -62.9441,
  -62.8413,
  -62.7383,
  -62.6357,
  -62.5338,
  -62.433,
  -62.3337,
  -62.2362,
  -62.141,
  -62.0482,
  -61.9582,
  -61.8716,
  -61.7887,
  -61.709,
  -61.6325,
  -61.5583,
  -61.4859,
  -61.4142,
  -61.3423,
  -61.2699,
  -61.1965,
  -61.1222,
  -61.0473,
  -60.9723,
  -60.8977,
  -60.8246,
  -60.7534,
  -60.6849,
  -60.6194,
  -60.5572,
  -60.4987,
  -60.4443,
  -60.394,
  -60.3481,
  -60.3062,
  -60.2685,
  -60.2348,
  -60.2053,
  -60.1801,
  -60.158,
  -60.141,
  -60.1267,
  -60.1136,
  -60.1008,
  -60.0875,
  -60.0726,
  -60.0557,
  -60.0364,
  -60.016,
  -59.9949,
  -59.9749,
  -59.9568,
  -59.9415,
  -59.9293,
  -59.9208,
  -59.9164,
  -59.9162,
  -49.8081,
  -49.9935,
  -50.1778,
  -50.3625,
  -50.5499,
  -50.7413,
  -50.9391,
  -51.1435,
  -51.3529,
  -51.5696,
  -51.7916,
  -52.0186,
  -52.2505,
  -52.4876,
  -52.7304,
  -52.979,
  -53.2343,
  -53.497,
  -53.7671,
  -54.0448,
  -54.3302,
  -54.6232,
  -54.9228,
  -55.2265,
  -55.5342,
  -55.8426,
  -56.1496,
  -56.4528,
  -56.7504,
  -57.0408,
  -57.3212,
  -57.5891,
  -57.8432,
  -58.0827,
  -58.3072,
  -58.5175,
  -58.7143,
  -58.8992,
  -59.0729,
  -59.2394,
  -59.3995,
  -59.5545,
  -59.7056,
  -59.853,
  -59.9968,
  -60.1369,
  -60.2728,
  -60.4043,
  -60.5309,
  -60.6527,
  -60.7698,
  -60.8824,
  -60.9911,
  -61.0967,
  -61.1987,
  -61.2991,
  -61.3967,
  -61.4913,
  -61.5829,
  -61.6716,
  -61.758,
  -61.8423,
  -61.9265,
  -62.0096,
  -62.0924,
  -62.1742,
  -62.2556,
  -62.3361,
  -62.4161,
  -62.496,
  -62.5757,
  -62.655,
  -62.7357,
  -62.8177,
  -62.9012,
  -62.9865,
  -63.0742,
  -63.1645,
  -63.2575,
  -63.3527,
  -63.4497,
  -63.5482,
  -63.6485,
  -63.7506,
  -63.8548,
  -63.9611,
  -64.0698,
  -64.1799,
  -64.2906,
  -64.4002,
  -64.5096,
  -64.6169,
  -64.7209,
  -64.8213,
  -64.9181,
  -65.0111,
  -65.1005,
  -65.1866,
  -65.2703,
  -65.3517,
  -65.4314,
  -65.5108,
  -65.5908,
  -65.6719,
  -65.7547,
  -65.8394,
  -65.9255,
  -66.0125,
  -66.0985,
  -66.1848,
  -66.2697,
  -66.3517,
  -66.4303,
  -66.505,
  -66.5755,
  -66.6419,
  -66.7047,
  -66.7643,
  -66.8218,
  -66.8782,
  -66.934,
  -66.9899,
  -67.0461,
  -67.1033,
  -67.1621,
  -67.2223,
  -67.2843,
  -67.3477,
  -67.4116,
  -67.4772,
  -67.5428,
  -67.6083,
  -67.673,
  -67.7372,
  -67.8004,
  -67.8625,
  -67.9233,
  -67.983,
  -68.0412,
  -68.0976,
  -68.1514,
  -68.2026,
  -68.2506,
  -68.2951,
  -68.3362,
  -68.3734,
  -68.4066,
  -68.4353,
  -68.4595,
  -68.4799,
  -68.4955,
  -68.5085,
  -68.518,
  -68.5242,
  -68.5272,
  -68.5266,
  -68.5227,
  -68.5151,
  -68.5044,
  -68.4907,
  -68.474,
  -68.4545,
  -68.4321,
  -68.4072,
  -68.3802,
  -68.3511,
  -68.3206,
  -68.2881,
  -68.2541,
  -68.2189,
  -68.1822,
  -68.1444,
  -68.1055,
  -68.0657,
  -68.024,
  -67.9819,
  -67.9383,
  -67.8927,
  -67.8451,
  -67.7954,
  -67.7434,
  -67.6893,
  -67.6328,
  -67.5739,
  -67.5126,
  -67.4483,
  -67.3813,
  -67.3118,
  -67.2399,
  -67.1659,
  -67.0902,
  -67.0134,
  -66.9359,
  -66.8583,
  -66.7813,
  -66.7044,
  -66.6276,
  -66.5508,
  -66.4738,
  -66.3966,
  -66.3173,
  -66.2381,
  -66.1569,
  -66.074,
  -65.9893,
  -65.9031,
  -65.8159,
  -65.7274,
  -65.6378,
  -65.5469,
  -65.4549,
  -65.3616,
  -65.2672,
  -65.1726,
  -65.0788,
  -64.9867,
  -64.8974,
  -64.8116,
  -64.7298,
  -64.6521,
  -64.5776,
  -64.5054,
  -64.4349,
  -64.3654,
  -64.2966,
  -64.228,
  -64.1594,
  -64.0909,
  -64.0225,
  -63.9545,
  -63.8873,
  -63.8201,
  -63.7542,
  -63.6882,
  -63.6209,
  -63.551,
  -63.4777,
  -63.3999,
  -63.3172,
  -63.2296,
  -63.1371,
  -63.0401,
  -62.9395,
  -62.8363,
  -62.7317,
  -62.6265,
  -62.5215,
  -62.4175,
  -62.3145,
  -62.2131,
  -62.1136,
  -62.0161,
  -61.921,
  -61.8289,
  -61.7404,
  -61.6555,
  -61.5744,
  -61.4971,
  -61.4233,
  -61.3526,
  -61.2838,
  -61.2162,
  -61.1488,
  -61.0808,
  -61.012,
  -60.9417,
  -60.8701,
  -60.7979,
  -60.7249,
  -60.6541,
  -60.5857,
  -60.5201,
  -60.4577,
  -60.3988,
  -60.344,
  -60.2933,
  -60.2467,
  -60.2042,
  -60.1655,
  -60.1304,
  -60.099,
  -60.0716,
  -60.0482,
  -60.0288,
  -60.0131,
  -59.9995,
  -59.9871,
  -59.9746,
  -59.9611,
  -59.9461,
  -59.9291,
  -59.9104,
  -59.8906,
  -59.8706,
  -59.8516,
  -59.8346,
  -59.8205,
  -59.8098,
  -59.8031,
  -59.801,
  -59.8035,
  -49.5906,
  -49.7803,
  -49.9692,
  -50.1575,
  -50.3489,
  -50.5446,
  -50.746,
  -50.9542,
  -51.169,
  -51.3897,
  -51.6163,
  -51.8481,
  -52.085,
  -52.3272,
  -52.5751,
  -52.8293,
  -53.0896,
  -53.3564,
  -53.6315,
  -53.914,
  -54.2043,
  -54.5017,
  -54.8057,
  -55.1144,
  -55.4257,
  -55.7372,
  -56.0467,
  -56.352,
  -56.6513,
  -56.943,
  -57.2246,
  -57.4933,
  -57.7469,
  -57.9865,
  -58.2111,
  -58.4214,
  -58.6181,
  -58.803,
  -58.9774,
  -59.1434,
  -59.3028,
  -59.4567,
  -59.6065,
  -59.7523,
  -59.8944,
  -60.0327,
  -60.1669,
  -60.2969,
  -60.4209,
  -60.5409,
  -60.6558,
  -60.7659,
  -60.8719,
  -60.9744,
  -61.0742,
  -61.1712,
  -61.2658,
  -61.3575,
  -61.4466,
  -61.5333,
  -61.6181,
  -61.7017,
  -61.7845,
  -61.867,
  -61.9492,
  -62.0301,
  -62.112,
  -62.1938,
  -62.2756,
  -62.3576,
  -62.4395,
  -62.5218,
  -62.6048,
  -62.6886,
  -62.7738,
  -62.8603,
  -62.9493,
  -63.0409,
  -63.1351,
  -63.2315,
  -63.3301,
  -63.4309,
  -63.5338,
  -63.6385,
  -63.7466,
  -63.8574,
  -63.9701,
  -64.0846,
  -64.1998,
  -64.3145,
  -64.4277,
  -64.5384,
  -64.6456,
  -64.749,
  -64.8485,
  -64.9439,
  -65.0352,
  -65.1227,
  -65.2068,
  -65.288,
  -65.367,
  -65.4439,
  -65.5218,
  -65.6013,
  -65.6828,
  -65.7663,
  -65.852,
  -65.9391,
  -66.0266,
  -66.1134,
  -66.1985,
  -66.2804,
  -66.3581,
  -66.4312,
  -66.4998,
  -66.5642,
  -66.625,
  -66.6827,
  -66.7385,
  -66.7937,
  -66.8485,
  -66.9032,
  -66.959,
  -67.016,
  -67.0746,
  -67.1348,
  -67.1971,
  -67.2609,
  -67.3264,
  -67.393,
  -67.4603,
  -67.5282,
  -67.5956,
  -67.6625,
  -67.7288,
  -67.7936,
  -67.857,
  -67.9191,
  -67.9795,
  -68.0378,
  -68.0933,
  -68.1459,
  -68.1937,
  -68.2389,
  -68.2807,
  -68.3182,
  -68.3515,
  -68.3802,
  -68.4042,
  -68.424,
  -68.4399,
  -68.4524,
  -68.4612,
  -68.4667,
  -68.4688,
  -68.4674,
  -68.4626,
  -68.4541,
  -68.4424,
  -68.4275,
  -68.4095,
  -68.3887,
  -68.3649,
  -68.3387,
  -68.3107,
  -68.2799,
  -68.2491,
  -68.2168,
  -68.183,
  -68.1479,
  -68.1113,
  -68.0737,
  -68.0346,
  -67.9944,
  -67.9531,
  -67.9104,
  -67.8664,
  -67.8207,
  -67.7731,
  -67.7236,
  -67.6719,
  -67.6185,
  -67.563,
  -67.5051,
  -67.445,
  -67.3824,
  -67.3173,
  -67.2496,
  -67.1798,
  -67.1083,
  -67.034,
  -66.9594,
  -66.8835,
  -66.8072,
  -66.7309,
  -66.6542,
  -66.5774,
  -66.5002,
  -66.4226,
  -66.3444,
  -66.2651,
  -66.1844,
  -66.1019,
  -66.0177,
  -65.9318,
  -65.8441,
  -65.7549,
  -65.6634,
  -65.5704,
  -65.4753,
  -65.378,
  -65.2792,
  -65.1789,
  -65.0782,
  -64.978,
  -64.8795,
  -64.7837,
  -64.691,
  -64.6024,
  -64.5166,
  -64.4355,
  -64.357,
  -64.2802,
  -64.2049,
  -64.1302,
  -64.0561,
  -63.9825,
  -63.9093,
  -63.8367,
  -63.7653,
  -63.6949,
  -63.6256,
  -63.5571,
  -63.4886,
  -63.4186,
  -63.346,
  -63.2696,
  -63.1886,
  -63.1026,
  -63.0113,
  -62.9151,
  -62.8146,
  -62.7107,
  -62.6046,
  -62.4976,
  -62.3903,
  -62.2838,
  -62.1784,
  -62.0748,
  -61.973,
  -61.8738,
  -61.777,
  -61.6829,
  -61.5912,
  -61.5047,
  -61.4221,
  -61.3438,
  -61.2695,
  -61.1992,
  -61.1322,
  -61.0675,
  -61.0044,
  -60.9418,
  -60.8787,
  -60.8145,
  -60.7486,
  -60.681,
  -60.6123,
  -60.5432,
  -60.4755,
  -60.4101,
  -60.3477,
  -60.2888,
  -60.2335,
  -60.1823,
  -60.1353,
  -60.0927,
  -60.0538,
  -60.0181,
  -59.9858,
  -59.9568,
  -59.9313,
  -59.9096,
  -59.8915,
  -59.8762,
  -59.8628,
  -59.8499,
  -59.8365,
  -59.822,
  -59.8059,
  -59.7883,
  -59.7693,
  -59.7498,
  -59.7306,
  -59.7129,
  -59.6974,
  -59.6852,
  -59.6766,
  -59.6717,
  -59.6724,
  -59.6782,
  -49.3614,
  -49.5556,
  -49.7485,
  -49.9415,
  -50.1368,
  -50.3361,
  -50.5408,
  -50.7521,
  -50.9704,
  -51.195,
  -51.4257,
  -51.6621,
  -51.9029,
  -52.1502,
  -52.4032,
  -52.6628,
  -52.9284,
  -53.2008,
  -53.4807,
  -53.7679,
  -54.0623,
  -54.3635,
  -54.6709,
  -54.9829,
  -55.2973,
  -55.6115,
  -55.9233,
  -56.2298,
  -56.5309,
  -56.8241,
  -57.1069,
  -57.377,
  -57.6325,
  -57.873,
  -58.0984,
  -58.3094,
  -58.5069,
  -58.6924,
  -58.8676,
  -59.0341,
  -59.1937,
  -59.3476,
  -59.4967,
  -59.6405,
  -59.7813,
  -59.9181,
  -60.0508,
  -60.1789,
  -60.302,
  -60.4196,
  -60.532,
  -60.639,
  -60.7418,
  -60.8407,
  -60.9366,
  -61.0297,
  -61.1203,
  -61.2083,
  -61.294,
  -61.3769,
  -61.4595,
  -61.5412,
  -61.6226,
  -61.7037,
  -61.785,
  -61.8666,
  -61.9488,
  -62.0317,
  -62.1151,
  -62.1988,
  -62.2828,
  -62.3671,
  -62.452,
  -62.5377,
  -62.6243,
  -62.7124,
  -62.8017,
  -62.8944,
  -62.9893,
  -63.0869,
  -63.1871,
  -63.2902,
  -63.3963,
  -63.5057,
  -63.6185,
  -63.734,
  -63.8522,
  -63.9716,
  -64.0915,
  -64.2107,
  -64.328,
  -64.443,
  -64.5543,
  -64.6614,
  -64.7634,
  -64.8618,
  -64.9557,
  -65.0449,
  -65.1298,
  -65.2111,
  -65.2891,
  -65.3656,
  -65.4416,
  -65.519,
  -65.5985,
  -65.6806,
  -65.7655,
  -65.8522,
  -65.9396,
  -66.0263,
  -66.1106,
  -66.1912,
  -66.2674,
  -66.3385,
  -66.4041,
  -66.466,
  -66.5245,
  -66.5804,
  -66.6347,
  -66.6886,
  -66.7429,
  -66.798,
  -66.8541,
  -66.9113,
  -66.9698,
  -67.0299,
  -67.0923,
  -67.1566,
  -67.2225,
  -67.29,
  -67.3589,
  -67.4288,
  -67.4988,
  -67.5682,
  -67.636,
  -67.7035,
  -67.7699,
  -67.8345,
  -67.8968,
  -67.9567,
  -68.0136,
  -68.0673,
  -68.1174,
  -68.1634,
  -68.2056,
  -68.2432,
  -68.2766,
  -68.3051,
  -68.3287,
  -68.3481,
  -68.3634,
  -68.3752,
  -68.3835,
  -68.3884,
  -68.3898,
  -68.3878,
  -68.3814,
  -68.3724,
  -68.3598,
  -68.3438,
  -68.3245,
  -68.3024,
  -68.2774,
  -68.2501,
  -68.221,
  -68.1906,
  -68.1594,
  -68.1272,
  -68.0935,
  -68.0583,
  -68.0215,
  -67.9834,
  -67.9443,
  -67.9036,
  -67.8618,
  -67.8183,
  -67.7737,
  -67.7279,
  -67.6804,
  -67.6316,
  -67.5804,
  -67.5266,
  -67.4724,
  -67.4158,
  -67.3573,
  -67.2963,
  -67.2332,
  -67.1681,
  -67.1005,
  -67.0312,
  -66.9603,
  -66.8879,
  -66.8142,
  -66.7395,
  -66.664,
  -66.5876,
  -66.5108,
  -66.4335,
  -66.3556,
  -66.2766,
  -66.1964,
  -66.1146,
  -66.0311,
  -65.9458,
  -65.8588,
  -65.7698,
  -65.6785,
  -65.5852,
  -65.4879,
  -65.3889,
  -65.2871,
  -65.1833,
  -65.078,
  -64.9718,
  -64.8663,
  -64.762,
  -64.6601,
  -64.5611,
  -64.4655,
  -64.3735,
  -64.2848,
  -64.199,
  -64.1151,
  -64.0327,
  -63.9513,
  -63.871,
  -63.7913,
  -63.7128,
  -63.6354,
  -63.5593,
  -63.4849,
  -63.4119,
  -63.3397,
  -63.2677,
  -63.1942,
  -63.1182,
  -63.0383,
  -62.954,
  -62.8643,
  -62.7696,
  -62.6688,
  -62.5651,
  -62.4582,
  -62.3497,
  -62.2404,
  -62.1315,
  -62.0237,
  -61.9173,
  -61.8132,
  -61.7115,
  -61.613,
  -61.5174,
  -61.4252,
  -61.337,
  -61.2529,
  -61.1735,
  -61.0988,
  -61.0286,
  -60.9624,
  -60.8996,
  -60.8395,
  -60.7811,
  -60.7234,
  -60.6653,
  -60.6061,
  -60.545,
  -60.482,
  -60.4174,
  -60.3523,
  -60.288,
  -60.2262,
  -60.1674,
  -60.1122,
  -60.0608,
  -60.0134,
  -59.9702,
  -59.9312,
  -59.8955,
  -59.8631,
  -59.8337,
  -59.8061,
  -59.7825,
  -59.7622,
  -59.7447,
  -59.7294,
  -59.7152,
  -59.7012,
  -59.6862,
  -59.67,
  -59.6521,
  -59.6331,
  -59.6133,
  -59.5936,
  -59.5751,
  -59.5586,
  -59.545,
  -59.5352,
  -59.5297,
  -59.5287,
  -59.5329,
  -59.5424,
  -49.1248,
  -49.3232,
  -49.5194,
  -49.7157,
  -49.914,
  -50.1163,
  -50.324,
  -50.5371,
  -50.7581,
  -50.9861,
  -51.2205,
  -51.461,
  -51.7075,
  -51.96,
  -52.218,
  -52.4822,
  -52.7528,
  -53.0302,
  -53.314,
  -53.6051,
  -53.9032,
  -54.2077,
  -54.5169,
  -54.8315,
  -55.1481,
  -55.4644,
  -55.7784,
  -56.088,
  -56.3912,
  -56.6861,
  -56.9706,
  -57.2422,
  -57.4993,
  -57.7414,
  -57.9684,
  -58.181,
  -58.3802,
  -58.5664,
  -58.7434,
  -58.9116,
  -59.0725,
  -59.2271,
  -59.3764,
  -59.5209,
  -59.6609,
  -59.7966,
  -59.9276,
  -60.0537,
  -60.1743,
  -60.2891,
  -60.3983,
  -60.502,
  -60.6009,
  -60.6949,
  -60.7865,
  -60.875,
  -60.961,
  -61.0448,
  -61.1264,
  -61.2068,
  -61.2865,
  -61.3657,
  -61.445,
  -61.5243,
  -61.6042,
  -61.6851,
  -61.7676,
  -61.8511,
  -61.9354,
  -62.0205,
  -62.1047,
  -62.1906,
  -62.2767,
  -62.3635,
  -62.4515,
  -62.5409,
  -62.6319,
  -62.7253,
  -62.8215,
  -62.9203,
  -63.0223,
  -63.1278,
  -63.2372,
  -63.3508,
  -63.4689,
  -63.5902,
  -63.7139,
  -63.8387,
  -63.9627,
  -64.0871,
  -64.2094,
  -64.3291,
  -64.4453,
  -64.5572,
  -64.6646,
  -64.7668,
  -64.8637,
  -64.9554,
  -65.0417,
  -65.1234,
  -65.201,
  -65.2758,
  -65.35,
  -65.425,
  -65.5023,
  -65.5824,
  -65.6657,
  -65.7502,
  -65.8367,
  -65.9223,
  -66.0051,
  -66.0836,
  -66.1573,
  -66.226,
  -66.2899,
  -66.3493,
  -66.4052,
  -66.4591,
  -66.5121,
  -66.5651,
  -66.619,
  -66.6743,
  -66.7307,
  -66.7882,
  -66.8472,
  -66.9078,
  -66.9703,
  -67.0338,
  -67.1002,
  -67.169,
  -67.2392,
  -67.3104,
  -67.3821,
  -67.454,
  -67.5257,
  -67.5961,
  -67.6646,
  -67.731,
  -67.7952,
  -67.8566,
  -67.9148,
  -67.9697,
  -68.0206,
  -68.0673,
  -68.1096,
  -68.1473,
  -68.1802,
  -68.2081,
  -68.2303,
  -68.2493,
  -68.2643,
  -68.2756,
  -68.2834,
  -68.2877,
  -68.2888,
  -68.2863,
  -68.2801,
  -68.2702,
  -68.2566,
  -68.2397,
  -68.2193,
  -68.1958,
  -68.1697,
  -68.1414,
  -68.1115,
  -68.0807,
  -68.049,
  -68.0166,
  -67.9828,
  -67.9477,
  -67.9106,
  -67.8719,
  -67.8308,
  -67.7894,
  -67.747,
  -67.7033,
  -67.6586,
  -67.6128,
  -67.5657,
  -67.5173,
  -67.4675,
  -67.4155,
  -67.3621,
  -67.307,
  -67.2504,
  -67.1916,
  -67.1305,
  -67.0674,
  -67.0024,
  -66.9357,
  -66.8669,
  -66.7968,
  -66.7251,
  -66.652,
  -66.5778,
  -66.5022,
  -66.4256,
  -66.3483,
  -66.2688,
  -66.1896,
  -66.1091,
  -66.0267,
  -65.9423,
  -65.8559,
  -65.7676,
  -65.6772,
  -65.5844,
  -65.4888,
  -65.3897,
  -65.2878,
  -65.1824,
  -65.0746,
  -64.9645,
  -64.8538,
  -64.7435,
  -64.6339,
  -64.5262,
  -64.4211,
  -64.3189,
  -64.2199,
  -64.1236,
  -64.03,
  -63.938,
  -63.8478,
  -63.759,
  -63.6716,
  -63.5855,
  -63.5009,
  -63.4167,
  -63.3358,
  -63.2564,
  -63.1788,
  -63.1022,
  -63.0256,
  -62.9481,
  -62.868,
  -62.7842,
  -62.696,
  -62.6027,
  -62.5044,
  -62.4014,
  -62.2947,
  -62.1852,
  -62.0742,
  -61.9632,
  -61.8531,
  -61.7439,
  -61.6368,
  -61.5327,
  -61.4316,
  -61.3341,
  -61.2402,
  -61.1506,
  -61.0654,
  -60.985,
  -60.9094,
  -60.8387,
  -60.7731,
  -60.7118,
  -60.6538,
  -60.5985,
  -60.5451,
  -60.4925,
  -60.4397,
  -60.3858,
  -60.329,
  -60.271,
  -60.2113,
  -60.1507,
  -60.091,
  -60.0333,
  -59.9787,
  -59.9276,
  -59.8803,
  -59.8366,
  -59.7971,
  -59.7614,
  -59.729,
  -59.6996,
  -59.6728,
  -59.6485,
  -59.6267,
  -59.6074,
  -59.5901,
  -59.5744,
  -59.559,
  -59.5432,
  -59.526,
  -59.5072,
  -59.487,
  -59.466,
  -59.4451,
  -59.4251,
  -59.407,
  -59.3919,
  -59.3805,
  -59.3734,
  -59.3711,
  -59.374,
  -59.3819,
  -59.3953,
  -48.881,
  -49.0832,
  -49.2814,
  -49.4805,
  -49.6813,
  -49.8859,
  -50.0956,
  -50.3119,
  -50.5352,
  -50.7659,
  -51.0038,
  -51.2481,
  -51.4986,
  -51.7555,
  -52.0182,
  -52.2866,
  -52.5603,
  -52.8417,
  -53.1297,
  -53.4238,
  -53.725,
  -54.0323,
  -54.3446,
  -54.6611,
  -54.9795,
  -55.2978,
  -55.6137,
  -55.9253,
  -56.2307,
  -56.5277,
  -56.8142,
  -57.087,
  -57.3465,
  -57.5911,
  -57.8207,
  -58.036,
  -58.2379,
  -58.428,
  -58.6077,
  -58.7786,
  -58.9418,
  -59.0982,
  -59.2486,
  -59.3935,
  -59.5331,
  -59.6677,
  -59.7969,
  -59.9196,
  -60.0375,
  -60.1491,
  -60.2545,
  -60.3541,
  -60.449,
  -60.5394,
  -60.6262,
  -60.7097,
  -60.7908,
  -60.8698,
  -60.9471,
  -61.0236,
  -61.0999,
  -61.1763,
  -61.253,
  -61.3305,
  -61.4079,
  -61.4877,
  -61.5694,
  -61.6527,
  -61.7372,
  -61.8226,
  -61.9083,
  -61.9945,
  -62.0814,
  -62.169,
  -62.2577,
  -62.3477,
  -62.4392,
  -62.5335,
  -62.6307,
  -62.7309,
  -62.8347,
  -62.9416,
  -63.0547,
  -63.173,
  -63.2961,
  -63.4232,
  -63.5526,
  -63.6832,
  -63.814,
  -63.9439,
  -64.072,
  -64.1973,
  -64.3195,
  -64.4371,
  -64.5501,
  -64.6572,
  -64.7585,
  -64.8533,
  -64.9418,
  -65.0242,
  -65.1005,
  -65.1741,
  -65.2462,
  -65.3188,
  -65.3934,
  -65.4712,
  -65.5521,
  -65.6354,
  -65.72,
  -65.8032,
  -65.8832,
  -65.959,
  -66.0298,
  -66.0953,
  -66.156,
  -66.2124,
  -66.266,
  -66.3181,
  -66.3699,
  -66.4215,
  -66.4756,
  -66.5311,
  -66.5881,
  -66.6465,
  -66.7062,
  -66.7674,
  -66.8301,
  -66.8951,
  -66.9625,
  -67.0319,
  -67.1031,
  -67.1758,
  -67.2494,
  -67.3236,
  -67.3974,
  -67.4697,
  -67.54,
  -67.6085,
  -67.6739,
  -67.7366,
  -67.7949,
  -67.8505,
  -67.9019,
  -67.9489,
  -67.9912,
  -68.0285,
  -68.0607,
  -68.0882,
  -68.1109,
  -68.1293,
  -68.1439,
  -68.155,
  -68.1625,
  -68.1664,
  -68.1668,
  -68.1635,
  -68.1564,
  -68.1458,
  -68.1313,
  -68.113,
  -68.0915,
  -68.067,
  -68.04,
  -68.0099,
  -67.9794,
  -67.9478,
  -67.9156,
  -67.8828,
  -67.8489,
  -67.8133,
  -67.7758,
  -67.7364,
  -67.6955,
  -67.6533,
  -67.6101,
  -67.5662,
  -67.5217,
  -67.4766,
  -67.4304,
  -67.3829,
  -67.3339,
  -67.2831,
  -67.2311,
  -67.1775,
  -67.1222,
  -67.0655,
  -67.0068,
  -66.9461,
  -66.8825,
  -66.8181,
  -66.7518,
  -66.6838,
  -66.6141,
  -66.5428,
  -66.4699,
  -66.3955,
  -66.3195,
  -66.2427,
  -66.1644,
  -66.0849,
  -66.0039,
  -65.9212,
  -65.8365,
  -65.7491,
  -65.6596,
  -65.5676,
  -65.4727,
  -65.3751,
  -65.2739,
  -65.1692,
  -65.0609,
  -64.9495,
  -64.8362,
  -64.7215,
  -64.6064,
  -64.4923,
  -64.3791,
  -64.267,
  -64.1585,
  -64.0524,
  -63.9487,
  -63.847,
  -63.7472,
  -63.649,
  -63.5522,
  -63.4573,
  -63.364,
  -63.2731,
  -63.1842,
  -63.0974,
  -63.0127,
  -62.9297,
  -62.8479,
  -62.7664,
  -62.6838,
  -62.5992,
  -62.5109,
  -62.4185,
  -62.3213,
  -62.2195,
  -62.1134,
  -62.0039,
  -61.892,
  -61.7791,
  -61.6662,
  -61.5544,
  -61.4444,
  -61.3371,
  -61.2331,
  -61.1327,
  -61.0367,
  -60.9443,
  -60.8576,
  -60.776,
  -60.6998,
  -60.6287,
  -60.5628,
  -60.5021,
  -60.4458,
  -60.3932,
  -60.3434,
  -60.2951,
  -60.2478,
  -60.2005,
  -60.1522,
  -60.102,
  -60.0497,
  -59.9955,
  -59.9406,
  -59.886,
  -59.8333,
  -59.7833,
  -59.7367,
  -59.6935,
  -59.6539,
  -59.6178,
  -59.5852,
  -59.5558,
  -59.529,
  -59.5046,
  -59.4822,
  -59.4618,
  -59.4431,
  -59.4256,
  -59.4089,
  -59.3919,
  -59.3737,
  -59.3538,
  -59.3324,
  -59.3096,
  -59.2866,
  -59.2641,
  -59.2437,
  -59.2263,
  -59.2114,
  -59.2022,
  -59.198,
  -59.1991,
  -59.2057,
  -59.2178,
  -59.2351,
  -48.6298,
  -48.8352,
  -49.0369,
  -49.2384,
  -49.4411,
  -49.6475,
  -49.8589,
  -50.0769,
  -50.3019,
  -50.5348,
  -50.7755,
  -51.0221,
  -51.2762,
  -51.5366,
  -51.8031,
  -52.0751,
  -52.353,
  -52.6377,
  -52.9284,
  -53.2254,
  -53.5286,
  -53.8378,
  -54.1519,
  -54.4697,
  -54.7896,
  -55.1095,
  -55.4265,
  -55.7406,
  -56.0484,
  -56.348,
  -56.637,
  -56.9138,
  -57.1765,
  -57.4246,
  -57.6581,
  -57.877,
  -58.0828,
  -58.2766,
  -58.46,
  -58.6345,
  -58.8009,
  -58.9599,
  -59.111,
  -59.2568,
  -59.3964,
  -59.5299,
  -59.6573,
  -59.7783,
  -59.8928,
  -60.0005,
  -60.1018,
  -60.1972,
  -60.2873,
  -60.3729,
  -60.4545,
  -60.533,
  -60.6088,
  -60.6829,
  -60.7548,
  -60.8272,
  -60.9002,
  -60.9736,
  -61.048,
  -61.1234,
  -61.2,
  -61.2783,
  -61.3585,
  -61.4404,
  -61.5237,
  -61.6082,
  -61.6933,
  -61.7791,
  -61.8657,
  -61.9535,
  -62.0421,
  -62.1313,
  -62.2235,
  -62.3185,
  -62.4166,
  -62.5179,
  -62.6237,
  -62.7346,
  -62.8512,
  -62.9738,
  -63.1017,
  -63.234,
  -63.3691,
  -63.5058,
  -63.6426,
  -63.7788,
  -63.9136,
  -64.0456,
  -64.1744,
  -64.2982,
  -64.4176,
  -64.5313,
  -64.6379,
  -64.737,
  -64.8281,
  -64.9117,
  -64.9892,
  -65.062,
  -65.1322,
  -65.2025,
  -65.2742,
  -65.3489,
  -65.4266,
  -65.5069,
  -65.5876,
  -65.6673,
  -65.7436,
  -65.8157,
  -65.8819,
  -65.9438,
  -66.0011,
  -66.0547,
  -66.1059,
  -66.1564,
  -66.2074,
  -66.2599,
  -66.3142,
  -66.3704,
  -66.4286,
  -66.4882,
  -66.5488,
  -66.6106,
  -66.6741,
  -66.7398,
  -66.8079,
  -66.8781,
  -66.9506,
  -67.0245,
  -67.0997,
  -67.1745,
  -67.2501,
  -67.3244,
  -67.3964,
  -67.4658,
  -67.5324,
  -67.5959,
  -67.6557,
  -67.7117,
  -67.7633,
  -67.8102,
  -67.852,
  -67.8889,
  -67.9206,
  -67.9473,
  -67.9694,
  -67.9873,
  -68.0017,
  -68.0123,
  -68.0191,
  -68.0224,
  -68.0219,
  -68.0169,
  -68.0089,
  -67.997,
  -67.9813,
  -67.9619,
  -67.9394,
  -67.914,
  -67.8862,
  -67.8563,
  -67.825,
  -67.7929,
  -67.7601,
  -67.7267,
  -67.692,
  -67.6559,
  -67.618,
  -67.578,
  -67.5363,
  -67.4934,
  -67.4496,
  -67.4059,
  -67.3619,
  -67.3177,
  -67.2726,
  -67.2253,
  -67.1775,
  -67.1281,
  -67.0772,
  -67.0253,
  -66.9717,
  -66.9168,
  -66.8602,
  -66.8018,
  -66.7417,
  -66.6797,
  -66.6159,
  -66.5501,
  -66.4823,
  -66.4127,
  -66.3413,
  -66.2686,
  -66.1941,
  -66.1179,
  -66.0402,
  -65.9607,
  -65.8796,
  -65.7966,
  -65.7114,
  -65.6235,
  -65.5327,
  -65.4392,
  -65.3412,
  -65.2412,
  -65.1374,
  -65.0302,
  -64.9198,
  -64.8057,
  -64.6897,
  -64.5714,
  -64.4524,
  -64.3335,
  -64.2155,
  -64.0986,
  -63.9834,
  -63.8703,
  -63.7594,
  -63.6502,
  -63.5426,
  -63.4366,
  -63.3323,
  -63.23,
  -63.1298,
  -63.032,
  -62.9368,
  -62.844,
  -62.7535,
  -62.6649,
  -62.5775,
  -62.4903,
  -62.4024,
  -62.3125,
  -62.2197,
  -62.1229,
  -62.0207,
  -61.9153,
  -61.8061,
  -61.694,
  -61.5799,
  -61.465,
  -61.3505,
  -61.2374,
  -61.1266,
  -61.0188,
  -60.915,
  -60.8156,
  -60.7214,
  -60.6325,
  -60.5491,
  -60.4716,
  -60.3997,
  -60.3337,
  -60.2732,
  -60.2176,
  -60.1668,
  -60.1196,
  -60.0752,
  -60.0322,
  -59.9904,
  -59.9488,
  -59.9063,
  -59.8623,
  -59.8161,
  -59.7684,
  -59.7195,
  -59.6711,
  -59.624,
  -59.5795,
  -59.5376,
  -59.4988,
  -59.4632,
  -59.4306,
  -59.401,
  -59.373,
  -59.3484,
  -59.3257,
  -59.3048,
  -59.2852,
  -59.2666,
  -59.2485,
  -59.2303,
  -59.2111,
  -59.1903,
  -59.1677,
  -59.1435,
  -59.1181,
  -59.0933,
  -59.0701,
  -59.0496,
  -59.0324,
  -59.0199,
  -59.0126,
  -59.0111,
  -59.0154,
  -59.0256,
  -59.0415,
  -59.0628,
  -48.374,
  -48.5817,
  -48.7858,
  -48.9885,
  -49.1929,
  -49.4005,
  -49.612,
  -49.8309,
  -50.057,
  -50.2913,
  -50.5339,
  -50.7839,
  -51.041,
  -51.3041,
  -51.5733,
  -51.8484,
  -52.129,
  -52.4155,
  -52.7082,
  -53.0067,
  -53.3115,
  -53.6209,
  -53.9361,
  -54.2552,
  -54.5767,
  -54.8987,
  -55.2189,
  -55.5356,
  -55.8465,
  -56.1491,
  -56.4414,
  -56.7217,
  -56.9887,
  -57.2413,
  -57.4793,
  -57.7031,
  -57.9125,
  -58.1111,
  -58.299,
  -58.4778,
  -58.6482,
  -58.8103,
  -58.965,
  -59.1121,
  -59.2519,
  -59.3845,
  -59.5096,
  -59.6276,
  -59.7383,
  -59.8418,
  -59.9385,
  -60.0289,
  -60.1127,
  -60.193,
  -60.2693,
  -60.3426,
  -60.4136,
  -60.4832,
  -60.5521,
  -60.6212,
  -60.691,
  -60.7621,
  -60.8342,
  -60.9073,
  -60.9817,
  -61.0576,
  -61.135,
  -61.2142,
  -61.295,
  -61.3761,
  -61.4592,
  -61.5439,
  -61.6296,
  -61.7167,
  -61.8052,
  -61.8954,
  -61.988,
  -62.0832,
  -62.182,
  -62.2848,
  -62.3924,
  -62.5058,
  -62.6254,
  -62.7516,
  -62.8838,
  -63.0209,
  -63.1614,
  -63.3029,
  -63.4464,
  -63.5896,
  -63.7317,
  -63.8715,
  -64.0083,
  -64.1411,
  -64.2687,
  -64.3896,
  -64.5025,
  -64.6065,
  -64.7011,
  -64.7869,
  -64.8652,
  -64.9376,
  -65.0065,
  -65.0745,
  -65.1433,
  -65.2133,
  -65.2868,
  -65.3623,
  -65.4383,
  -65.513,
  -65.5847,
  -65.6523,
  -65.7149,
  -65.773,
  -65.8268,
  -65.8775,
  -65.9268,
  -65.9759,
  -66.0265,
  -66.0788,
  -66.1339,
  -66.1912,
  -66.2506,
  -66.3115,
  -66.3733,
  -66.4353,
  -66.5,
  -66.5667,
  -66.6359,
  -66.7071,
  -66.7806,
  -66.8561,
  -66.9329,
  -67.0104,
  -67.0873,
  -67.1628,
  -67.236,
  -67.3062,
  -67.3733,
  -67.437,
  -67.4968,
  -67.5525,
  -67.6039,
  -67.6505,
  -67.692,
  -67.7283,
  -67.7594,
  -67.7844,
  -67.8059,
  -67.8233,
  -67.8366,
  -67.8463,
  -67.8522,
  -67.8547,
  -67.8532,
  -67.8478,
  -67.8385,
  -67.8252,
  -67.8083,
  -67.7878,
  -67.7643,
  -67.738,
  -67.7094,
  -67.679,
  -67.6471,
  -67.6142,
  -67.5806,
  -67.5462,
  -67.5109,
  -67.4739,
  -67.434,
  -67.3932,
  -67.351,
  -67.308,
  -67.2645,
  -67.2208,
  -67.1774,
  -67.1341,
  -67.0905,
  -67.0457,
  -66.9993,
  -66.9514,
  -66.9021,
  -66.8518,
  -66.8002,
  -66.7471,
  -66.6924,
  -66.6359,
  -66.5785,
  -66.519,
  -66.4576,
  -66.3938,
  -66.328,
  -66.2606,
  -66.1913,
  -66.12,
  -66.0461,
  -65.9712,
  -65.8944,
  -65.8153,
  -65.7343,
  -65.651,
  -65.565,
  -65.4763,
  -65.3844,
  -65.289,
  -65.1901,
  -65.0876,
  -64.9817,
  -64.8722,
  -64.7595,
  -64.6435,
  -64.5249,
  -64.4042,
  -64.2818,
  -64.1588,
  -64.0355,
  -63.9127,
  -63.7913,
  -63.6712,
  -63.5528,
  -63.4361,
  -63.321,
  -63.2079,
  -63.0967,
  -62.9876,
  -62.88,
  -62.7759,
  -62.6744,
  -62.5754,
  -62.4787,
  -62.3841,
  -62.2908,
  -62.1979,
  -62.1044,
  -62.0092,
  -61.9113,
  -61.81,
  -61.7049,
  -61.596,
  -61.4837,
  -61.3691,
  -61.2527,
  -61.136,
  -61.0198,
  -60.9054,
  -60.7939,
  -60.686,
  -60.5827,
  -60.4846,
  -60.3923,
  -60.3062,
  -60.2263,
  -60.1528,
  -60.0856,
  -60.0246,
  -59.9692,
  -59.9189,
  -59.873,
  -59.8309,
  -59.7916,
  -59.7544,
  -59.7172,
  -59.6814,
  -59.6452,
  -59.6077,
  -59.5685,
  -59.5277,
  -59.4858,
  -59.444,
  -59.4034,
  -59.3645,
  -59.328,
  -59.294,
  -59.2625,
  -59.2334,
  -59.2067,
  -59.1821,
  -59.1593,
  -59.1379,
  -59.1177,
  -59.0982,
  -59.079,
  -59.0597,
  -59.0397,
  -59.0184,
  -58.995,
  -58.9698,
  -58.9432,
  -58.9161,
  -58.8899,
  -58.866,
  -58.8452,
  -58.8285,
  -58.8168,
  -58.8108,
  -58.8111,
  -58.8179,
  -58.8311,
  -58.8504,
  -58.8752,
  -48.1135,
  -48.3219,
  -48.5268,
  -48.7304,
  -48.9356,
  -49.1437,
  -49.357,
  -49.5765,
  -49.8034,
  -50.0382,
  -50.2819,
  -50.5335,
  -50.7926,
  -51.0578,
  -51.329,
  -51.6048,
  -51.887,
  -52.1748,
  -52.4686,
  -52.7679,
  -53.0735,
  -53.3846,
  -53.701,
  -54.021,
  -54.3439,
  -54.6679,
  -54.9909,
  -55.3106,
  -55.6246,
  -55.9308,
  -56.2259,
  -56.5105,
  -56.7824,
  -57.0403,
  -57.2841,
  -57.5135,
  -57.7294,
  -57.9332,
  -58.126,
  -58.3095,
  -58.484,
  -58.65,
  -58.8075,
  -58.9563,
  -59.0963,
  -59.2276,
  -59.3494,
  -59.4637,
  -59.5702,
  -59.6691,
  -59.7608,
  -59.846,
  -59.9255,
  -60.0004,
  -60.0716,
  -60.1399,
  -60.2067,
  -60.2723,
  -60.3379,
  -60.4041,
  -60.4714,
  -60.5402,
  -60.6103,
  -60.6801,
  -60.7518,
  -60.8245,
  -60.8983,
  -60.9735,
  -61.0502,
  -61.1287,
  -61.2088,
  -61.2913,
  -61.3755,
  -61.4617,
  -61.5499,
  -61.6397,
  -61.732,
  -61.8274,
  -61.9266,
  -62.0304,
  -62.1387,
  -62.2544,
  -62.3767,
  -62.5057,
  -62.6412,
  -62.7822,
  -62.9275,
  -63.0759,
  -63.2262,
  -63.377,
  -63.5272,
  -63.6756,
  -63.8214,
  -63.9636,
  -64.1001,
  -64.2294,
  -64.3495,
  -64.4592,
  -64.5583,
  -64.6459,
  -64.726,
  -64.7989,
  -64.867,
  -64.9328,
  -64.9981,
  -65.0646,
  -65.133,
  -65.2026,
  -65.2724,
  -65.3412,
  -65.4072,
  -65.4694,
  -65.5273,
  -65.581,
  -65.6317,
  -65.68,
  -65.7277,
  -65.7758,
  -65.8249,
  -65.8778,
  -65.9337,
  -65.9925,
  -66.0535,
  -66.1158,
  -66.1794,
  -66.2439,
  -66.3101,
  -66.378,
  -66.4478,
  -66.5203,
  -66.5954,
  -66.6723,
  -66.7506,
  -66.8294,
  -66.9073,
  -66.9836,
  -67.0575,
  -67.1282,
  -67.1952,
  -67.2575,
  -67.3168,
  -67.3721,
  -67.4229,
  -67.4692,
  -67.5104,
  -67.5462,
  -67.5769,
  -67.6023,
  -67.623,
  -67.6395,
  -67.6516,
  -67.6601,
  -67.6648,
  -67.6656,
  -67.6626,
  -67.6554,
  -67.6444,
  -67.6296,
  -67.6111,
  -67.5895,
  -67.5648,
  -67.5378,
  -67.5077,
  -67.4767,
  -67.4439,
  -67.4101,
  -67.3757,
  -67.3402,
  -67.3036,
  -67.2654,
  -67.2253,
  -67.184,
  -67.1416,
  -67.0986,
  -67.0554,
  -67.0125,
  -66.9701,
  -66.9279,
  -66.8856,
  -66.8425,
  -66.798,
  -66.7522,
  -66.7048,
  -66.6562,
  -66.6063,
  -66.555,
  -66.5024,
  -66.4475,
  -66.3917,
  -66.3344,
  -66.2749,
  -66.2138,
  -66.1503,
  -66.0849,
  -66.0178,
  -65.9485,
  -65.8773,
  -65.8039,
  -65.7281,
  -65.65,
  -65.5691,
  -65.4854,
  -65.3988,
  -65.3088,
  -65.2152,
  -65.1179,
  -65.017,
  -64.9123,
  -64.804,
  -64.6922,
  -64.5771,
  -64.4593,
  -64.3385,
  -64.2154,
  -64.0901,
  -63.9622,
  -63.8343,
  -63.7059,
  -63.5779,
  -63.4509,
  -63.3252,
  -63.2013,
  -63.0795,
  -62.9599,
  -62.8427,
  -62.7277,
  -62.6154,
  -62.5057,
  -62.3986,
  -62.2936,
  -62.191,
  -62.0902,
  -61.991,
  -61.8923,
  -61.7933,
  -61.6929,
  -61.59,
  -61.4843,
  -61.3755,
  -61.2632,
  -61.148,
  -61.0307,
  -60.9122,
  -60.7937,
  -60.676,
  -60.5605,
  -60.4483,
  -60.3404,
  -60.2368,
  -60.1399,
  -60.0498,
  -59.9666,
  -59.8901,
  -59.8204,
  -59.7578,
  -59.7015,
  -59.6508,
  -59.6054,
  -59.5644,
  -59.5268,
  -59.4923,
  -59.4601,
  -59.4296,
  -59.3996,
  -59.3696,
  -59.3389,
  -59.3068,
  -59.2736,
  -59.2393,
  -59.2049,
  -59.1711,
  -59.1388,
  -59.1081,
  -59.0794,
  -59.0524,
  -59.027,
  -59.0031,
  -58.9806,
  -58.959,
  -58.9383,
  -58.9179,
  -58.8978,
  -58.8774,
  -58.8563,
  -58.8343,
  -58.8108,
  -58.785,
  -58.7575,
  -58.729,
  -58.7008,
  -58.6739,
  -58.6488,
  -58.6281,
  -58.6117,
  -58.6004,
  -58.5952,
  -58.5967,
  -58.6052,
  -58.6206,
  -58.6426,
  -58.6705,
  -47.8465,
  -48.0571,
  -48.2622,
  -48.466,
  -48.6712,
  -48.8798,
  -49.0933,
  -49.313,
  -49.54,
  -49.7748,
  -50.0178,
  -50.2703,
  -50.5299,
  -50.7965,
  -51.0692,
  -51.347,
  -51.6302,
  -51.9186,
  -52.2128,
  -52.5129,
  -52.8189,
  -53.131,
  -53.4482,
  -53.7694,
  -54.0941,
  -54.419,
  -54.7441,
  -55.0668,
  -55.3841,
  -55.6938,
  -55.9941,
  -56.2834,
  -56.5605,
  -56.8242,
  -57.074,
  -57.3096,
  -57.5314,
  -57.741,
  -57.9393,
  -58.1278,
  -58.3071,
  -58.4757,
  -58.6358,
  -58.7858,
  -58.9257,
  -59.0553,
  -59.175,
  -59.2852,
  -59.387,
  -59.4805,
  -59.5669,
  -59.6469,
  -59.7214,
  -59.7913,
  -59.8581,
  -59.9227,
  -59.986,
  -60.0477,
  -60.1108,
  -60.175,
  -60.2405,
  -60.3071,
  -60.3749,
  -60.4432,
  -60.5118,
  -60.5806,
  -60.6501,
  -60.7203,
  -60.7923,
  -60.8663,
  -60.9426,
  -61.0219,
  -61.1037,
  -61.1885,
  -61.2745,
  -61.3636,
  -61.4553,
  -61.5505,
  -61.65,
  -61.7545,
  -61.8649,
  -61.982,
  -62.1059,
  -62.2369,
  -62.3749,
  -62.5195,
  -62.6693,
  -62.8234,
  -62.9806,
  -63.1393,
  -63.2982,
  -63.4561,
  -63.6107,
  -63.7628,
  -63.909,
  -64.0474,
  -64.1757,
  -64.2923,
  -64.3969,
  -64.4898,
  -64.5725,
  -64.6465,
  -64.7141,
  -64.7775,
  -64.8391,
  -64.9006,
  -64.9629,
  -65.0259,
  -65.0886,
  -65.1507,
  -65.2101,
  -65.2651,
  -65.3179,
  -65.3675,
  -65.4151,
  -65.4613,
  -65.5072,
  -65.5549,
  -65.6051,
  -65.6589,
  -65.7158,
  -65.7759,
  -65.8385,
  -65.9028,
  -65.9687,
  -66.0353,
  -66.1029,
  -66.172,
  -66.2433,
  -66.3177,
  -66.3944,
  -66.4717,
  -66.5511,
  -66.6306,
  -66.7094,
  -66.7862,
  -66.8601,
  -66.9305,
  -66.9971,
  -67.0599,
  -67.1187,
  -67.1734,
  -67.2238,
  -67.2695,
  -67.3103,
  -67.3458,
  -67.3758,
  -67.4008,
  -67.4206,
  -67.4359,
  -67.4468,
  -67.4535,
  -67.4562,
  -67.4538,
  -67.4485,
  -67.4392,
  -67.4259,
  -67.4088,
  -67.3885,
  -67.3654,
  -67.3399,
  -67.3121,
  -67.2822,
  -67.2506,
  -67.2173,
  -67.1828,
  -67.147,
  -67.1102,
  -67.072,
  -67.0324,
  -66.9914,
  -66.9493,
  -66.9066,
  -66.8639,
  -66.8215,
  -66.7796,
  -66.7386,
  -66.6979,
  -66.6563,
  -66.6149,
  -66.5729,
  -66.5292,
  -66.4838,
  -66.437,
  -66.3894,
  -66.3401,
  -66.2893,
  -66.2374,
  -66.1837,
  -66.1286,
  -66.0713,
  -66.0123,
  -65.9511,
  -65.8879,
  -65.8227,
  -65.7555,
  -65.6861,
  -65.614,
  -65.5393,
  -65.4621,
  -65.3817,
  -65.2977,
  -65.21,
  -65.1183,
  -65.023,
  -64.9225,
  -64.8192,
  -64.712,
  -64.6012,
  -64.4873,
  -64.3701,
  -64.2501,
  -64.1273,
  -64.0018,
  -63.8738,
  -63.7434,
  -63.611,
  -63.4772,
  -63.3427,
  -63.2091,
  -63.0765,
  -62.9458,
  -62.8179,
  -62.6926,
  -62.5702,
  -62.4507,
  -62.3337,
  -62.2192,
  -62.107,
  -61.997,
  -61.8889,
  -61.7826,
  -61.6775,
  -61.5731,
  -61.4688,
  -61.3635,
  -61.2553,
  -61.1457,
  -61.0332,
  -60.9179,
  -60.8001,
  -60.6805,
  -60.5599,
  -60.4394,
  -60.3204,
  -60.2042,
  -60.0915,
  -59.9839,
  -59.8822,
  -59.7871,
  -59.699,
  -59.6184,
  -59.5453,
  -59.4795,
  -59.4208,
  -59.3684,
  -59.3216,
  -59.2801,
  -59.2428,
  -59.2095,
  -59.1792,
  -59.1518,
  -59.1264,
  -59.1025,
  -59.0789,
  -59.055,
  -59.0305,
  -59.005,
  -58.9788,
  -58.9521,
  -58.9256,
  -58.9003,
  -58.8759,
  -58.8527,
  -58.8296,
  -58.808,
  -58.787,
  -58.7663,
  -58.7458,
  -58.7252,
  -58.7043,
  -58.6829,
  -58.6609,
  -58.6379,
  -58.6139,
  -58.5882,
  -58.5607,
  -58.5318,
  -58.5021,
  -58.473,
  -58.4457,
  -58.4211,
  -58.4002,
  -58.3837,
  -58.3724,
  -58.3673,
  -58.3691,
  -58.3783,
  -58.395,
  -58.4189,
  -58.4494,
  -47.5753,
  -47.7861,
  -47.9912,
  -48.1946,
  -48.3992,
  -48.6064,
  -48.8195,
  -49.039,
  -49.2658,
  -49.5003,
  -49.7437,
  -49.9961,
  -50.2567,
  -50.5241,
  -50.7973,
  -51.0755,
  -51.3588,
  -51.6476,
  -51.942,
  -52.2429,
  -52.5488,
  -52.8616,
  -53.1804,
  -53.5033,
  -53.8294,
  -54.1569,
  -54.4844,
  -54.8091,
  -55.1291,
  -55.4422,
  -55.7465,
  -56.0404,
  -56.3229,
  -56.5923,
  -56.848,
  -57.0889,
  -57.317,
  -57.5325,
  -57.7364,
  -57.93,
  -58.1133,
  -58.2863,
  -58.4485,
  -58.5992,
  -58.7382,
  -58.8654,
  -58.9814,
  -59.087,
  -59.1835,
  -59.2715,
  -59.3524,
  -59.4263,
  -59.4962,
  -59.5624,
  -59.6258,
  -59.6876,
  -59.7487,
  -59.8097,
  -59.8715,
  -59.9344,
  -59.9984,
  -60.0632,
  -60.1288,
  -60.1943,
  -60.2594,
  -60.3238,
  -60.3879,
  -60.4529,
  -60.5184,
  -60.5873,
  -60.6591,
  -60.7346,
  -60.8137,
  -60.8961,
  -60.9813,
  -61.0692,
  -61.1602,
  -61.2549,
  -61.3541,
  -61.4586,
  -61.5694,
  -61.6869,
  -61.8118,
  -61.9443,
  -62.0843,
  -62.2306,
  -62.3846,
  -62.5444,
  -62.7084,
  -62.8751,
  -63.0432,
  -63.2113,
  -63.3774,
  -63.5398,
  -63.6964,
  -63.8446,
  -63.9819,
  -64.1066,
  -64.2178,
  -64.316,
  -64.4018,
  -64.4774,
  -64.5447,
  -64.6058,
  -64.6625,
  -64.7183,
  -64.7739,
  -64.8296,
  -64.885,
  -64.9391,
  -64.9912,
  -65.0412,
  -65.0889,
  -65.1344,
  -65.1788,
  -65.223,
  -65.2682,
  -65.3157,
  -65.3665,
  -65.4211,
  -65.4793,
  -65.5411,
  -65.6059,
  -65.6727,
  -65.7395,
  -65.8079,
  -65.8772,
  -65.9483,
  -66.0218,
  -66.098,
  -66.176,
  -66.2554,
  -66.3359,
  -66.416,
  -66.4951,
  -66.5718,
  -66.6453,
  -66.7153,
  -66.7814,
  -66.8436,
  -66.9017,
  -66.9559,
  -67.006,
  -67.0513,
  -67.0918,
  -67.1258,
  -67.1555,
  -67.1798,
  -67.1989,
  -67.2129,
  -67.222,
  -67.2266,
  -67.2268,
  -67.2226,
  -67.2145,
  -67.202,
  -67.1857,
  -67.1662,
  -67.1438,
  -67.1191,
  -67.0923,
  -67.0635,
  -67.033,
  -67.0006,
  -66.9666,
  -66.9308,
  -66.8937,
  -66.8554,
  -66.8157,
  -66.7736,
  -66.7314,
  -66.6885,
  -66.6458,
  -66.6036,
  -66.5621,
  -66.5214,
  -66.4816,
  -66.4428,
  -66.4041,
  -66.3651,
  -66.3247,
  -66.2832,
  -66.2403,
  -66.1961,
  -66.1505,
  -66.1031,
  -66.0545,
  -66.0046,
  -65.9529,
  -65.8997,
  -65.8445,
  -65.7873,
  -65.7284,
  -65.6674,
  -65.6043,
  -65.5376,
  -65.4695,
  -65.3991,
  -65.3256,
  -65.2489,
  -65.1684,
  -65.0841,
  -64.9958,
  -64.9026,
  -64.8053,
  -64.7034,
  -64.5972,
  -64.4875,
  -64.3742,
  -64.2579,
  -64.1381,
  -64.0158,
  -63.8909,
  -63.763,
  -63.6323,
  -63.4982,
  -63.3615,
  -63.2227,
  -63.0827,
  -62.9429,
  -62.804,
  -62.6673,
  -62.5337,
  -62.4039,
  -62.2764,
  -62.1532,
  -62.0326,
  -61.9144,
  -61.7982,
  -61.6838,
  -61.5709,
  -61.4597,
  -61.3495,
  -61.2401,
  -61.1307,
  -61.0209,
  -60.9098,
  -60.7966,
  -60.6811,
  -60.5631,
  -60.443,
  -60.3213,
  -60.1989,
  -60.077,
  -59.9569,
  -59.84,
  -59.7274,
  -59.6204,
  -59.5198,
  -59.4266,
  -59.3408,
  -59.263,
  -59.1929,
  -59.1303,
  -59.0748,
  -59.0255,
  -58.9819,
  -58.9432,
  -58.9092,
  -58.8781,
  -58.8516,
  -58.8282,
  -58.8075,
  -58.789,
  -58.7719,
  -58.7549,
  -58.7377,
  -58.7201,
  -58.7017,
  -58.683,
  -58.6643,
  -58.6461,
  -58.6285,
  -58.6112,
  -58.5941,
  -58.5767,
  -58.5586,
  -58.5397,
  -58.5199,
  -58.4992,
  -58.4775,
  -58.4548,
  -58.431,
  -58.4063,
  -58.3803,
  -58.353,
  -58.324,
  -58.294,
  -58.2636,
  -58.2341,
  -58.2064,
  -58.1814,
  -58.1601,
  -58.143,
  -58.131,
  -58.1252,
  -58.1263,
  -58.1353,
  -58.1524,
  -58.1776,
  -58.21,
  -47.2962,
  -47.5065,
  -47.7113,
  -47.9139,
  -48.1175,
  -48.3249,
  -48.5375,
  -48.756,
  -48.9822,
  -49.2162,
  -49.4589,
  -49.7106,
  -49.9712,
  -50.2392,
  -50.5118,
  -50.7904,
  -51.0739,
  -51.3631,
  -51.658,
  -51.9601,
  -52.2687,
  -52.5835,
  -52.9041,
  -53.2287,
  -53.5561,
  -53.8849,
  -54.2135,
  -54.5397,
  -54.8618,
  -55.1775,
  -55.484,
  -55.7819,
  -56.069,
  -56.3438,
  -56.6053,
  -56.8532,
  -57.0873,
  -57.3087,
  -57.518,
  -57.7157,
  -57.9026,
  -58.0781,
  -58.2413,
  -58.3917,
  -58.5289,
  -58.652,
  -58.7635,
  -58.8639,
  -58.9545,
  -59.0368,
  -59.1125,
  -59.1828,
  -59.2491,
  -59.3125,
  -59.3741,
  -59.4346,
  -59.4951,
  -59.5558,
  -59.6173,
  -59.6795,
  -59.7424,
  -59.8057,
  -59.868,
  -59.9303,
  -59.9914,
  -60.0509,
  -60.1098,
  -60.1689,
  -60.2295,
  -60.2929,
  -60.3597,
  -60.4311,
  -60.5065,
  -60.5861,
  -60.6693,
  -60.7556,
  -60.8452,
  -60.939,
  -61.0377,
  -61.1407,
  -61.2509,
  -61.3683,
  -61.4935,
  -61.6267,
  -61.7682,
  -61.9184,
  -62.0763,
  -62.2412,
  -62.4122,
  -62.5872,
  -62.7649,
  -62.9431,
  -63.1199,
  -63.2931,
  -63.4606,
  -63.6196,
  -63.7668,
  -63.8996,
  -64.0185,
  -64.1226,
  -64.2124,
  -64.2896,
  -64.3564,
  -64.4152,
  -64.4685,
  -64.5187,
  -64.5673,
  -64.6151,
  -64.6624,
  -64.7085,
  -64.7536,
  -64.7972,
  -64.8396,
  -64.8809,
  -64.9226,
  -64.9654,
  -65.01,
  -65.0568,
  -65.1081,
  -65.1642,
  -65.2243,
  -65.2883,
  -65.3551,
  -65.4239,
  -65.4938,
  -65.5644,
  -65.636,
  -65.7094,
  -65.785,
  -65.8627,
  -65.9423,
  -66.0229,
  -66.1039,
  -66.1843,
  -66.2633,
  -66.3398,
  -66.4128,
  -66.4822,
  -66.5465,
  -66.6082,
  -66.6661,
  -66.7196,
  -66.7693,
  -66.8143,
  -66.8546,
  -66.8895,
  -66.9189,
  -66.9426,
  -66.9606,
  -66.9731,
  -66.9801,
  -66.982,
  -66.9792,
  -66.9716,
  -66.9599,
  -66.944,
  -66.9244,
  -66.9018,
  -66.8769,
  -66.8503,
  -66.8211,
  -66.7912,
  -66.7597,
  -66.7262,
  -66.6911,
  -66.6542,
  -66.6156,
  -66.5754,
  -66.5338,
  -66.4912,
  -66.4479,
  -66.4044,
  -66.3616,
  -66.3195,
  -66.2791,
  -66.2399,
  -66.2018,
  -66.1645,
  -66.1278,
  -66.0909,
  -66.0529,
  -66.0135,
  -65.9728,
  -65.9307,
  -65.8873,
  -65.8415,
  -65.7953,
  -65.7473,
  -65.6974,
  -65.6459,
  -65.5929,
  -65.5377,
  -65.4805,
  -65.421,
  -65.3596,
  -65.2957,
  -65.2287,
  -65.1592,
  -65.0864,
  -65.0104,
  -64.9301,
  -64.8452,
  -64.756,
  -64.6615,
  -64.562,
  -64.4579,
  -64.3492,
  -64.2365,
  -64.1201,
  -64.0009,
  -63.8789,
  -63.754,
  -63.6266,
  -63.4948,
  -63.361,
  -63.2235,
  -63.0825,
  -62.9391,
  -62.7941,
  -62.649,
  -62.5049,
  -62.3633,
  -62.2253,
  -62.0914,
  -61.9619,
  -61.836,
  -61.7128,
  -61.5919,
  -61.4728,
  -61.3551,
  -61.2387,
  -61.1233,
  -61.0087,
  -60.895,
  -60.7815,
  -60.6677,
  -60.553,
  -60.4366,
  -60.3185,
  -60.1982,
  -60.0761,
  -59.9528,
  -59.8292,
  -59.7063,
  -59.5856,
  -59.4685,
  -59.3554,
  -59.2493,
  -59.1503,
  -59.0589,
  -58.9758,
  -58.9006,
  -58.8332,
  -58.7733,
  -58.7202,
  -58.6732,
  -58.6318,
  -58.5955,
  -58.5637,
  -58.5362,
  -58.5129,
  -58.4931,
  -58.4767,
  -58.463,
  -58.4515,
  -58.4412,
  -58.4311,
  -58.4208,
  -58.4103,
  -58.3995,
  -58.3887,
  -58.3778,
  -58.3668,
  -58.3556,
  -58.3436,
  -58.3303,
  -58.3152,
  -58.2982,
  -58.2794,
  -58.2587,
  -58.2363,
  -58.2124,
  -58.1873,
  -58.1609,
  -58.1335,
  -58.105,
  -58.0751,
  -58.0445,
  -58.0126,
  -57.9828,
  -57.9546,
  -57.9289,
  -57.9066,
  -57.8882,
  -57.8748,
  -57.8674,
  -57.8671,
  -57.875,
  -57.8916,
  -57.917,
  -57.9507,
  -47.0101,
  -47.2193,
  -47.4233,
  -47.6251,
  -47.8275,
  -48.0336,
  -48.2452,
  -48.4627,
  -48.6879,
  -48.9201,
  -49.1622,
  -49.4132,
  -49.6739,
  -49.9421,
  -50.2162,
  -50.4954,
  -50.7798,
  -51.07,
  -51.3667,
  -51.6705,
  -51.9815,
  -52.2991,
  -52.622,
  -52.9485,
  -53.2761,
  -53.6053,
  -53.934,
  -54.2605,
  -54.5833,
  -54.9004,
  -55.2102,
  -55.511,
  -55.8018,
  -56.081,
  -56.3473,
  -56.6008,
  -56.8408,
  -57.0675,
  -57.2815,
  -57.483,
  -57.6712,
  -57.8476,
  -58.0103,
  -58.1589,
  -58.2928,
  -58.4127,
  -58.5196,
  -58.6141,
  -58.6989,
  -58.7757,
  -58.8464,
  -58.9131,
  -58.9768,
  -59.0389,
  -59.1002,
  -59.1612,
  -59.2215,
  -59.2832,
  -59.3451,
  -59.4074,
  -59.4697,
  -59.5316,
  -59.5924,
  -59.6515,
  -59.7082,
  -59.7629,
  -59.8161,
  -59.8693,
  -59.9239,
  -59.9814,
  -60.043,
  -60.1098,
  -60.1815,
  -60.2567,
  -60.3373,
  -60.4213,
  -60.5094,
  -60.6025,
  -60.7,
  -60.8028,
  -60.912,
  -61.0286,
  -61.1535,
  -61.2869,
  -61.4301,
  -61.5826,
  -61.7445,
  -61.9147,
  -62.0924,
  -62.2756,
  -62.4624,
  -62.6501,
  -62.8378,
  -63.0224,
  -63.2013,
  -63.3713,
  -63.5295,
  -63.673,
  -63.8004,
  -63.9108,
  -64.0049,
  -64.0842,
  -64.1505,
  -64.2068,
  -64.2556,
  -64.3,
  -64.3418,
  -64.3816,
  -64.4206,
  -64.4591,
  -64.4958,
  -64.5333,
  -64.5704,
  -64.6081,
  -64.6471,
  -64.6884,
  -64.7328,
  -64.7812,
  -64.834,
  -64.8916,
  -64.9536,
  -65.0198,
  -65.0884,
  -65.1591,
  -65.231,
  -65.3041,
  -65.3787,
  -65.4544,
  -65.5318,
  -65.6109,
  -65.6907,
  -65.7724,
  -65.8539,
  -65.9345,
  -66.0131,
  -66.0891,
  -66.1618,
  -66.2304,
  -66.2952,
  -66.3562,
  -66.4136,
  -66.4673,
  -66.5166,
  -66.5615,
  -66.6017,
  -66.6365,
  -66.6657,
  -66.6887,
  -66.7052,
  -66.7156,
  -66.7203,
  -66.7193,
  -66.7119,
  -66.7006,
  -66.6846,
  -66.6648,
  -66.6416,
  -66.6157,
  -66.588,
  -66.559,
  -66.529,
  -66.4978,
  -66.465,
  -66.4304,
  -66.3938,
  -66.3553,
  -66.315,
  -66.2727,
  -66.2291,
  -66.1847,
  -66.1402,
  -66.0963,
  -66.0532,
  -66.0117,
  -65.9721,
  -65.9344,
  -65.8973,
  -65.8617,
  -65.8266,
  -65.7914,
  -65.7556,
  -65.719,
  -65.6803,
  -65.64,
  -65.5989,
  -65.5566,
  -65.5131,
  -65.4671,
  -65.4193,
  -65.3697,
  -65.318,
  -65.2649,
  -65.2088,
  -65.1506,
  -65.0899,
  -65.0269,
  -64.9614,
  -64.8923,
  -64.82,
  -64.7437,
  -64.6636,
  -64.5788,
  -64.488,
  -64.3911,
  -64.2898,
  -64.1832,
  -64.0721,
  -63.9564,
  -63.837,
  -63.7144,
  -63.5894,
  -63.4624,
  -63.3317,
  -63.1978,
  -63.0602,
  -62.919,
  -62.7744,
  -62.6265,
  -62.4772,
  -62.3278,
  -62.1799,
  -62.0347,
  -61.8935,
  -61.7569,
  -61.625,
  -61.4972,
  -61.3725,
  -61.2497,
  -61.1288,
  -61.0088,
  -60.8897,
  -60.7714,
  -60.6536,
  -60.5362,
  -60.4185,
  -60.3014,
  -60.1836,
  -60.0647,
  -59.9443,
  -59.8222,
  -59.6987,
  -59.574,
  -59.4495,
  -59.3263,
  -59.2056,
  -59.0891,
  -58.9778,
  -58.8732,
  -58.7761,
  -58.687,
  -58.6062,
  -58.5337,
  -58.4689,
  -58.4114,
  -58.3602,
  -58.3151,
  -58.2753,
  -58.2405,
  -58.2106,
  -58.1851,
  -58.1642,
  -58.1475,
  -58.1348,
  -58.1255,
  -58.1189,
  -58.1144,
  -58.1108,
  -58.1076,
  -58.1044,
  -58.1012,
  -58.0977,
  -58.0928,
  -58.0883,
  -58.0829,
  -58.0759,
  -58.0667,
  -58.0548,
  -58.0399,
  -58.0224,
  -58.0023,
  -57.9798,
  -57.9553,
  -57.9291,
  -57.9017,
  -57.8731,
  -57.8438,
  -57.8136,
  -57.7826,
  -57.7517,
  -57.7212,
  -57.6923,
  -57.6655,
  -57.6416,
  -57.6214,
  -57.6058,
  -57.5961,
  -57.5936,
  -57.5995,
  -57.6148,
  -57.6396,
  -57.674,
  -46.7138,
  -46.922,
  -47.1247,
  -47.3255,
  -47.5258,
  -47.7305,
  -47.9405,
  -48.1568,
  -48.3806,
  -48.613,
  -48.8546,
  -49.1056,
  -49.3662,
  -49.6349,
  -49.9102,
  -50.191,
  -50.4775,
  -50.7701,
  -51.0698,
  -51.3756,
  -51.6899,
  -52.0107,
  -52.3362,
  -52.6646,
  -52.9935,
  -53.322,
  -53.6499,
  -53.9754,
  -54.2975,
  -54.6145,
  -54.9248,
  -55.2272,
  -55.5204,
  -55.8032,
  -56.0723,
  -56.3306,
  -56.5756,
  -56.8069,
  -57.0246,
  -57.2285,
  -57.4185,
  -57.5942,
  -57.7549,
  -57.9,
  -58.0297,
  -58.1445,
  -58.2453,
  -58.3344,
  -58.4135,
  -58.4853,
  -58.5513,
  -58.6152,
  -58.6778,
  -58.7402,
  -58.8026,
  -58.8657,
  -58.9292,
  -58.9926,
  -59.0557,
  -59.1186,
  -59.1806,
  -59.2411,
  -59.2993,
  -59.355,
  -59.4076,
  -59.4572,
  -59.5047,
  -59.5507,
  -59.5994,
  -59.6513,
  -59.7078,
  -59.7698,
  -59.8374,
  -59.9101,
  -59.9873,
  -60.0692,
  -60.1552,
  -60.2471,
  -60.3429,
  -60.4439,
  -60.5516,
  -60.6668,
  -60.7909,
  -60.9249,
  -61.0685,
  -61.2237,
  -61.3896,
  -61.5653,
  -61.7496,
  -61.9409,
  -62.1369,
  -62.3358,
  -62.5347,
  -62.7309,
  -62.9216,
  -63.1033,
  -63.2727,
  -63.4263,
  -63.5624,
  -63.6798,
  -63.7784,
  -63.8596,
  -63.9256,
  -63.9785,
  -64.0232,
  -64.0618,
  -64.0964,
  -64.1287,
  -64.1599,
  -64.1903,
  -64.221,
  -64.2522,
  -64.2845,
  -64.3187,
  -64.3554,
  -64.3956,
  -64.4401,
  -64.4894,
  -64.5438,
  -64.6031,
  -64.6671,
  -64.7349,
  -64.8053,
  -64.8766,
  -64.9509,
  -65.0266,
  -65.1036,
  -65.1816,
  -65.261,
  -65.3416,
  -65.4234,
  -65.5058,
  -65.5875,
  -65.6682,
  -65.7465,
  -65.822,
  -65.894,
  -65.9621,
  -66.0267,
  -66.0874,
  -66.1446,
  -66.1981,
  -66.2474,
  -66.2924,
  -66.3315,
  -66.3662,
  -66.395,
  -66.4167,
  -66.4317,
  -66.4399,
  -66.4417,
  -66.4371,
  -66.4268,
  -66.4112,
  -66.391,
  -66.367,
  -66.3399,
  -66.3105,
  -66.2798,
  -66.2483,
  -66.2161,
  -66.1831,
  -66.1487,
  -66.1125,
  -66.0741,
  -66.0335,
  -65.9909,
  -65.9453,
  -65.8996,
  -65.8533,
  -65.8075,
  -65.7627,
  -65.7196,
  -65.6788,
  -65.6402,
  -65.604,
  -65.5694,
  -65.5356,
  -65.5023,
  -65.4688,
  -65.435,
  -65.4001,
  -65.3636,
  -65.3259,
  -65.2869,
  -65.2469,
  -65.2056,
  -65.1621,
  -65.1167,
  -65.0688,
  -65.0187,
  -64.9662,
  -64.911,
  -64.8526,
  -64.7925,
  -64.7299,
  -64.6644,
  -64.5957,
  -64.5236,
  -64.4475,
  -64.367,
  -64.2812,
  -64.1896,
  -64.0923,
  -63.9889,
  -63.8802,
  -63.7662,
  -63.6476,
  -63.5253,
  -63.3997,
  -63.2716,
  -63.1409,
  -63.0069,
  -62.8696,
  -62.7282,
  -62.5829,
  -62.4341,
  -62.2824,
  -62.1296,
  -61.9771,
  -61.8267,
  -61.6795,
  -61.5355,
  -61.3975,
  -61.2642,
  -61.1354,
  -61.0099,
  -60.8864,
  -60.7643,
  -60.643,
  -60.5224,
  -60.4022,
  -60.2821,
  -60.1624,
  -60.0429,
  -59.9233,
  -59.8032,
  -59.6821,
  -59.5599,
  -59.4364,
  -59.3116,
  -59.1862,
  -59.0614,
  -58.9385,
  -58.8187,
  -58.7034,
  -58.5938,
  -58.4911,
  -58.3961,
  -58.3095,
  -58.2313,
  -58.1614,
  -58.0992,
  -58.0439,
  -57.9946,
  -57.951,
  -57.9126,
  -57.8782,
  -57.8496,
  -57.8257,
  -57.8067,
  -57.7926,
  -57.7831,
  -57.7775,
  -57.7753,
  -57.7755,
  -57.7775,
  -57.7806,
  -57.7839,
  -57.7874,
  -57.7904,
  -57.7931,
  -57.7947,
  -57.7948,
  -57.7927,
  -57.7875,
  -57.779,
  -57.7668,
  -57.7511,
  -57.7321,
  -57.7101,
  -57.6856,
  -57.659,
  -57.6311,
  -57.6021,
  -57.5726,
  -57.5422,
  -57.511,
  -57.4797,
  -57.4489,
  -57.4189,
  -57.3906,
  -57.3647,
  -57.3421,
  -57.3238,
  -57.3111,
  -57.3057,
  -57.3088,
  -57.3218,
  -57.3454,
  -57.3798,
  -46.4057,
  -46.612,
  -46.8132,
  -47.0125,
  -47.2126,
  -47.4154,
  -47.6235,
  -47.8385,
  -48.0611,
  -48.2925,
  -48.5338,
  -48.785,
  -49.046,
  -49.3164,
  -49.5927,
  -49.8764,
  -50.1665,
  -50.4633,
  -50.7674,
  -51.0788,
  -51.3966,
  -51.7204,
  -52.0481,
  -52.3774,
  -52.7059,
  -53.0333,
  -53.3593,
  -53.6828,
  -54.0028,
  -54.3175,
  -54.6275,
  -54.9305,
  -55.225,
  -55.5101,
  -55.7836,
  -56.0453,
  -56.2939,
  -56.5281,
  -56.7477,
  -56.952,
  -57.1411,
  -57.3142,
  -57.4713,
  -57.6116,
  -57.7348,
  -57.8438,
  -57.9391,
  -58.0225,
  -58.0968,
  -58.1649,
  -58.2293,
  -58.2923,
  -58.3553,
  -58.4192,
  -58.4843,
  -58.5504,
  -58.6166,
  -58.6824,
  -58.7474,
  -58.811,
  -58.8728,
  -58.9309,
  -58.987,
  -59.0393,
  -59.0878,
  -59.1328,
  -59.1749,
  -59.2161,
  -59.2589,
  -59.3051,
  -59.3565,
  -59.4136,
  -59.476,
  -59.5445,
  -59.6187,
  -59.6976,
  -59.7819,
  -59.8707,
  -59.964,
  -60.0629,
  -60.1689,
  -60.2828,
  -60.4064,
  -60.5411,
  -60.6874,
  -60.8456,
  -61.0159,
  -61.1973,
  -61.3885,
  -61.5878,
  -61.7932,
  -62.0023,
  -62.2124,
  -62.4204,
  -62.6229,
  -62.816,
  -62.9955,
  -63.1593,
  -63.3042,
  -63.4284,
  -63.5318,
  -63.6152,
  -63.6813,
  -63.7335,
  -63.7743,
  -63.8072,
  -63.8349,
  -63.8597,
  -63.8829,
  -63.9058,
  -63.9297,
  -63.9551,
  -63.9827,
  -64.0136,
  -64.0483,
  -64.0881,
  -64.1318,
  -64.1819,
  -64.2377,
  -64.2988,
  -64.3644,
  -64.4335,
  -64.5052,
  -64.5797,
  -64.6562,
  -64.7342,
  -64.813,
  -64.893,
  -64.9742,
  -65.0562,
  -65.139,
  -65.2216,
  -65.3036,
  -65.3841,
  -65.4622,
  -65.5374,
  -65.6079,
  -65.6757,
  -65.7402,
  -65.801,
  -65.8584,
  -65.9119,
  -65.9613,
  -66.0064,
  -66.0465,
  -66.0808,
  -66.1085,
  -66.129,
  -66.1422,
  -66.1478,
  -66.1463,
  -66.138,
  -66.1234,
  -66.1033,
  -66.0787,
  -66.0504,
  -66.0191,
  -65.986,
  -65.9522,
  -65.9168,
  -65.8822,
  -65.8466,
  -65.81,
  -65.7716,
  -65.7309,
  -65.6877,
  -65.6423,
  -65.5951,
  -65.5471,
  -65.499,
  -65.4518,
  -65.4062,
  -65.3631,
  -65.3229,
  -65.2856,
  -65.2508,
  -65.2176,
  -65.1853,
  -65.1538,
  -65.122,
  -65.0897,
  -65.0563,
  -65.0217,
  -64.9855,
  -64.949,
  -64.9115,
  -64.8722,
  -64.8312,
  -64.7882,
  -64.742,
  -64.6932,
  -64.641,
  -64.5861,
  -64.5287,
  -64.4686,
  -64.406,
  -64.3402,
  -64.2714,
  -64.1994,
  -64.1231,
  -64.0422,
  -63.9554,
  -63.8627,
  -63.7638,
  -63.6584,
  -63.5473,
  -63.4306,
  -63.3091,
  -63.1837,
  -63.0552,
  -62.9237,
  -62.7879,
  -62.6501,
  -62.5087,
  -62.3632,
  -62.2139,
  -62.061,
  -61.9059,
  -61.7503,
  -61.5958,
  -61.444,
  -61.296,
  -61.1527,
  -61.0147,
  -60.8816,
  -60.7527,
  -60.627,
  -60.5035,
  -60.3811,
  -60.2593,
  -60.1378,
  -60.0164,
  -59.8952,
  -59.7741,
  -59.653,
  -59.5317,
  -59.4099,
  -59.2874,
  -59.1637,
  -59.0392,
  -58.9138,
  -58.7883,
  -58.6641,
  -58.542,
  -58.4227,
  -58.3092,
  -58.2019,
  -58.1018,
  -58.0096,
  -57.9259,
  -57.8506,
  -57.7833,
  -57.7236,
  -57.6705,
  -57.6233,
  -57.5812,
  -57.5441,
  -57.5118,
  -57.4845,
  -57.4621,
  -57.4448,
  -57.4326,
  -57.4254,
  -57.4227,
  -57.4236,
  -57.4275,
  -57.4339,
  -57.4418,
  -57.4508,
  -57.46,
  -57.4691,
  -57.4775,
  -57.4847,
  -57.4902,
  -57.4928,
  -57.4919,
  -57.487,
  -57.4779,
  -57.4645,
  -57.4472,
  -57.4263,
  -57.4023,
  -57.376,
  -57.3482,
  -57.3192,
  -57.2887,
  -57.2585,
  -57.2276,
  -57.1961,
  -57.1645,
  -57.1334,
  -57.1033,
  -57.0752,
  -57.0499,
  -57.0284,
  -57.0123,
  -57.0032,
  -57.0031,
  -57.0136,
  -57.0358,
  -57.0701,
  -46.086,
  -46.2902,
  -46.4901,
  -46.6877,
  -46.8862,
  -47.0873,
  -47.2938,
  -47.5068,
  -47.7271,
  -47.9577,
  -48.1987,
  -48.4504,
  -48.7128,
  -48.9851,
  -49.2662,
  -49.5545,
  -49.8501,
  -50.1527,
  -50.4621,
  -50.7785,
  -51.1009,
  -51.4272,
  -51.7564,
  -52.0843,
  -52.4117,
  -52.737,
  -53.0604,
  -53.3807,
  -53.6978,
  -54.0115,
  -54.3201,
  -54.6226,
  -54.9179,
  -55.2042,
  -55.4796,
  -55.7431,
  -55.9936,
  -56.2291,
  -56.4486,
  -56.6507,
  -56.8368,
  -57.0061,
  -57.158,
  -57.2927,
  -57.411,
  -57.5138,
  -57.6033,
  -57.6818,
  -57.7523,
  -57.818,
  -57.8812,
  -57.9444,
  -58.0091,
  -58.0758,
  -58.1445,
  -58.2134,
  -58.2832,
  -58.3522,
  -58.4191,
  -58.4839,
  -58.5457,
  -58.6037,
  -58.6576,
  -58.707,
  -58.7518,
  -58.7922,
  -58.8294,
  -58.8657,
  -58.9033,
  -58.9442,
  -58.9898,
  -59.0415,
  -59.098,
  -59.1621,
  -59.2321,
  -59.3084,
  -59.3891,
  -59.4755,
  -59.5671,
  -59.6636,
  -59.7674,
  -59.8801,
  -60.0038,
  -60.1397,
  -60.2882,
  -60.4503,
  -60.6255,
  -60.8126,
  -61.011,
  -61.2185,
  -61.4321,
  -61.6515,
  -61.8728,
  -62.0923,
  -62.3063,
  -62.5106,
  -62.7017,
  -62.8753,
  -63.0284,
  -63.1595,
  -63.2676,
  -63.3539,
  -63.4207,
  -63.4711,
  -63.5086,
  -63.5364,
  -63.5576,
  -63.5749,
  -63.5907,
  -63.6055,
  -63.623,
  -63.6428,
  -63.666,
  -63.6938,
  -63.7269,
  -63.7662,
  -63.811,
  -63.8617,
  -63.9187,
  -63.9813,
  -64.0482,
  -64.1184,
  -64.1916,
  -64.2674,
  -64.3455,
  -64.4254,
  -64.506,
  -64.5875,
  -64.67,
  -64.7522,
  -64.8358,
  -64.9189,
  -65.0009,
  -65.0812,
  -65.1592,
  -65.2342,
  -65.3056,
  -65.3736,
  -65.4381,
  -65.4994,
  -65.5572,
  -65.611,
  -65.6606,
  -65.7057,
  -65.7454,
  -65.7791,
  -65.8055,
  -65.8242,
  -65.8349,
  -65.8375,
  -65.8325,
  -65.819,
  -65.8,
  -65.7752,
  -65.7458,
  -65.7129,
  -65.6773,
  -65.6405,
  -65.603,
  -65.5655,
  -65.5279,
  -65.4895,
  -65.45,
  -65.4087,
  -65.3651,
  -65.319,
  -65.2704,
  -65.2204,
  -65.1698,
  -65.1197,
  -65.0714,
  -65.0251,
  -64.982,
  -64.9425,
  -64.9056,
  -64.8724,
  -64.8406,
  -64.8101,
  -64.7798,
  -64.7493,
  -64.7189,
  -64.6869,
  -64.6546,
  -64.6214,
  -64.5872,
  -64.5526,
  -64.5155,
  -64.4766,
  -64.4352,
  -64.3909,
  -64.3434,
  -64.2914,
  -64.2365,
  -64.1782,
  -64.1176,
  -64.0547,
  -63.9884,
  -63.9193,
  -63.8466,
  -63.7699,
  -63.6886,
  -63.5999,
  -63.5057,
  -63.4048,
  -63.2976,
  -63.1842,
  -63.0647,
  -62.9407,
  -62.8122,
  -62.6802,
  -62.5453,
  -62.4066,
  -62.2643,
  -62.1181,
  -61.9683,
  -61.8149,
  -61.6581,
  -61.5,
  -61.3421,
  -61.1866,
  -61.0345,
  -60.8871,
  -60.7451,
  -60.6082,
  -60.4761,
  -60.3482,
  -60.2231,
  -60.1001,
  -59.9783,
  -59.8567,
  -59.735,
  -59.6125,
  -59.4909,
  -59.3693,
  -59.2477,
  -59.1256,
  -59.0032,
  -58.8797,
  -58.7554,
  -58.6303,
  -58.5049,
  -58.3801,
  -58.2569,
  -58.1366,
  -58.0201,
  -57.9092,
  -57.8049,
  -57.7081,
  -57.6192,
  -57.5387,
  -57.4666,
  -57.4023,
  -57.3451,
  -57.2943,
  -57.2491,
  -57.2087,
  -57.1731,
  -57.142,
  -57.1159,
  -57.0949,
  -57.0791,
  -57.0687,
  -57.0632,
  -57.0624,
  -57.0659,
  -57.0725,
  -57.0818,
  -57.0933,
  -57.1066,
  -57.1195,
  -57.1332,
  -57.1464,
  -57.1585,
  -57.1686,
  -57.1758,
  -57.1793,
  -57.1782,
  -57.1724,
  -57.1619,
  -57.1468,
  -57.1277,
  -57.1052,
  -57.0798,
  -57.0526,
  -57.0243,
  -56.9953,
  -56.9655,
  -56.935,
  -56.9035,
  -56.8714,
  -56.8391,
  -56.8073,
  -56.7768,
  -56.7487,
  -56.7237,
  -56.704,
  -56.6909,
  -56.6869,
  -56.6944,
  -56.7148,
  -56.7489,
  -45.7556,
  -45.957,
  -46.1544,
  -46.3491,
  -46.5456,
  -46.7455,
  -46.9503,
  -47.1621,
  -47.3825,
  -47.6126,
  -47.8534,
  -48.1058,
  -48.3706,
  -48.6456,
  -48.9309,
  -49.2248,
  -49.5264,
  -49.8355,
  -50.1502,
  -50.4718,
  -50.7975,
  -51.1262,
  -51.4557,
  -51.7838,
  -52.1096,
  -52.4323,
  -52.7521,
  -53.0689,
  -53.3831,
  -53.6938,
  -54.0009,
  -54.3028,
  -54.5979,
  -54.8838,
  -55.1602,
  -55.4242,
  -55.6741,
  -55.9082,
  -56.1257,
  -56.3254,
  -56.5073,
  -56.6711,
  -56.8173,
  -56.946,
  -57.058,
  -57.1552,
  -57.2396,
  -57.3142,
  -57.382,
  -57.4452,
  -57.5087,
  -57.5734,
  -57.641,
  -57.7115,
  -57.7843,
  -57.8582,
  -57.932,
  -58.004,
  -58.0735,
  -58.1394,
  -58.2014,
  -58.2588,
  -58.3109,
  -58.358,
  -58.3995,
  -58.4364,
  -58.469,
  -58.5009,
  -58.5342,
  -58.5696,
  -58.6098,
  -58.6558,
  -58.708,
  -58.7672,
  -58.8329,
  -58.9043,
  -58.9816,
  -59.0647,
  -59.1528,
  -59.247,
  -59.3494,
  -59.4613,
  -59.5856,
  -59.7219,
  -59.8743,
  -60.0407,
  -60.2214,
  -60.4149,
  -60.6208,
  -60.8367,
  -61.0606,
  -61.2902,
  -61.5222,
  -61.7523,
  -61.9769,
  -62.1916,
  -62.3921,
  -62.5746,
  -62.7355,
  -62.8729,
  -62.9859,
  -63.075,
  -63.142,
  -63.1913,
  -63.2258,
  -63.2491,
  -63.2644,
  -63.2753,
  -63.2844,
  -63.2933,
  -63.3046,
  -63.3192,
  -63.3385,
  -63.3634,
  -63.3949,
  -63.4328,
  -63.4775,
  -63.5287,
  -63.5865,
  -63.6499,
  -63.7177,
  -63.7879,
  -63.8624,
  -63.9395,
  -64.0183,
  -64.0992,
  -64.181,
  -64.2638,
  -64.3474,
  -64.4313,
  -64.5154,
  -64.5986,
  -64.6808,
  -64.7612,
  -64.8391,
  -64.9142,
  -64.9858,
  -65.0544,
  -65.1198,
  -65.1818,
  -65.2402,
  -65.2944,
  -65.3442,
  -65.3879,
  -65.427,
  -65.4596,
  -65.4843,
  -65.5008,
  -65.5086,
  -65.5078,
  -65.4988,
  -65.4818,
  -65.458,
  -65.4283,
  -65.3938,
  -65.3561,
  -65.3161,
  -65.2751,
  -65.2339,
  -65.1927,
  -65.1515,
  -65.1095,
  -65.0665,
  -65.0216,
  -64.9745,
  -64.9248,
  -64.8721,
  -64.8192,
  -64.7661,
  -64.7141,
  -64.6646,
  -64.6178,
  -64.575,
  -64.5365,
  -64.5017,
  -64.4699,
  -64.4396,
  -64.4103,
  -64.3819,
  -64.3526,
  -64.3233,
  -64.2931,
  -64.2627,
  -64.2321,
  -64.2008,
  -64.1684,
  -64.1336,
  -64.0967,
  -64.0575,
  -64.0144,
  -63.9674,
  -63.9149,
  -63.8594,
  -63.801,
  -63.7395,
  -63.6757,
  -63.6084,
  -63.5387,
  -63.4658,
  -63.3885,
  -63.3061,
  -63.2172,
  -63.1218,
  -63.0195,
  -62.9102,
  -62.7944,
  -62.6723,
  -62.5454,
  -62.4143,
  -62.2791,
  -62.1401,
  -61.9969,
  -61.85,
  -61.6991,
  -61.5446,
  -61.3869,
  -61.2266,
  -61.066,
  -60.9068,
  -60.7509,
  -60.5986,
  -60.4525,
  -60.3125,
  -60.1779,
  -60.0478,
  -59.9215,
  -59.7979,
  -59.6763,
  -59.5557,
  -59.4352,
  -59.3143,
  -59.1933,
  -59.0723,
  -58.9512,
  -58.8297,
  -58.7079,
  -58.5855,
  -58.4623,
  -58.3379,
  -58.2128,
  -58.0879,
  -57.9644,
  -57.8432,
  -57.7254,
  -57.6119,
  -57.5043,
  -57.4036,
  -57.3106,
  -57.2255,
  -57.1486,
  -57.0797,
  -57.0183,
  -56.9635,
  -56.9148,
  -56.8705,
  -56.8318,
  -56.7978,
  -56.7682,
  -56.7436,
  -56.7238,
  -56.7097,
  -56.7007,
  -56.6966,
  -56.697,
  -56.7016,
  -56.7099,
  -56.7214,
  -56.7356,
  -56.7516,
  -56.7688,
  -56.7863,
  -56.8035,
  -56.8197,
  -56.8339,
  -56.8452,
  -56.8528,
  -56.8557,
  -56.8533,
  -56.8458,
  -56.8334,
  -56.8164,
  -56.7956,
  -56.7721,
  -56.7464,
  -56.7194,
  -56.6914,
  -56.6626,
  -56.6329,
  -56.6018,
  -56.5693,
  -56.536,
  -56.5024,
  -56.4698,
  -56.4389,
  -56.4106,
  -56.387,
  -56.3698,
  -56.3622,
  -56.3667,
  -56.384,
  -56.4181,
  -45.4149,
  -45.6129,
  -45.8074,
  -46.0008,
  -46.1956,
  -46.3941,
  -46.5983,
  -46.8095,
  -47.0294,
  -47.2594,
  -47.5012,
  -47.7546,
  -48.0212,
  -48.2989,
  -48.5884,
  -48.8877,
  -49.1958,
  -49.5113,
  -49.8328,
  -50.1589,
  -50.4874,
  -50.8165,
  -51.1449,
  -51.4713,
  -51.7945,
  -52.1141,
  -52.4302,
  -52.7436,
  -53.0534,
  -53.362,
  -53.6674,
  -53.9684,
  -54.2633,
  -54.5501,
  -54.826,
  -55.0885,
  -55.336,
  -55.567,
  -55.7801,
  -55.9751,
  -56.1513,
  -56.3091,
  -56.4492,
  -56.571,
  -56.6776,
  -56.77,
  -56.8508,
  -56.9227,
  -56.989,
  -57.0529,
  -57.1174,
  -57.1846,
  -57.2557,
  -57.3302,
  -57.4073,
  -57.4857,
  -57.5633,
  -57.6388,
  -57.7107,
  -57.7781,
  -57.8395,
  -57.8966,
  -57.9478,
  -57.993,
  -58.0324,
  -58.0671,
  -58.0981,
  -58.1272,
  -58.1561,
  -58.1873,
  -58.2222,
  -58.2627,
  -58.3095,
  -58.3635,
  -58.4242,
  -58.491,
  -58.5641,
  -58.642,
  -58.7267,
  -58.8185,
  -58.9194,
  -59.0311,
  -59.156,
  -59.2966,
  -59.4526,
  -59.6243,
  -59.8108,
  -60.0116,
  -60.2253,
  -60.4496,
  -60.6824,
  -60.9216,
  -61.1629,
  -61.4027,
  -61.6365,
  -61.8591,
  -62.0679,
  -62.258,
  -62.4256,
  -62.5686,
  -62.6863,
  -62.7784,
  -62.8475,
  -62.8964,
  -62.9289,
  -62.9486,
  -62.9594,
  -62.9645,
  -62.9675,
  -62.9705,
  -62.9762,
  -62.9861,
  -63.0017,
  -63.0238,
  -63.0517,
  -63.0879,
  -63.1317,
  -63.1828,
  -63.2409,
  -63.3044,
  -63.3729,
  -63.4449,
  -63.52,
  -63.5974,
  -63.6767,
  -63.7579,
  -63.8404,
  -63.9238,
  -64.0079,
  -64.0921,
  -64.1764,
  -64.2598,
  -64.3419,
  -64.4223,
  -64.5005,
  -64.5753,
  -64.6478,
  -64.7173,
  -64.7837,
  -64.8467,
  -64.9063,
  -64.9611,
  -65.0111,
  -65.0555,
  -65.0936,
  -65.1245,
  -65.1469,
  -65.1607,
  -65.1652,
  -65.1605,
  -65.1471,
  -65.1254,
  -65.0964,
  -65.0613,
  -65.0215,
  -64.9785,
  -64.9336,
  -64.887,
  -64.8413,
  -64.796,
  -64.7505,
  -64.7044,
  -64.6571,
  -64.608,
  -64.5567,
  -64.5033,
  -64.4481,
  -64.3922,
  -64.3367,
  -64.2832,
  -64.2328,
  -64.1859,
  -64.1436,
  -64.1058,
  -64.0722,
  -64.0418,
  -64.0129,
  -63.9852,
  -63.9577,
  -63.9302,
  -63.9026,
  -63.8746,
  -63.8456,
  -63.8173,
  -63.7887,
  -63.7589,
  -63.7265,
  -63.6915,
  -63.6533,
  -63.6112,
  -63.5652,
  -63.5137,
  -63.4584,
  -63.3992,
  -63.3368,
  -63.2724,
  -63.2046,
  -63.1341,
  -63.0603,
  -62.9823,
  -62.8991,
  -62.8091,
  -62.7124,
  -62.6085,
  -62.4973,
  -62.3795,
  -62.2551,
  -62.1254,
  -61.991,
  -61.8516,
  -61.7086,
  -61.561,
  -61.4092,
  -61.2534,
  -61.0942,
  -60.9324,
  -60.7693,
  -60.6067,
  -60.4467,
  -60.2911,
  -60.1412,
  -59.9973,
  -59.8596,
  -59.7277,
  -59.6006,
  -59.477,
  -59.3557,
  -59.2361,
  -59.1172,
  -58.9983,
  -58.8792,
  -58.7596,
  -58.6399,
  -58.5202,
  -58.4001,
  -58.2794,
  -58.1577,
  -58.035,
  -57.9116,
  -57.7877,
  -57.6644,
  -57.5418,
  -57.4234,
  -57.3088,
  -57.1993,
  -57.0957,
  -56.9991,
  -56.9101,
  -56.8289,
  -56.7556,
  -56.6896,
  -56.6307,
  -56.5781,
  -56.5312,
  -56.4896,
  -56.4526,
  -56.4203,
  -56.3925,
  -56.3693,
  -56.3511,
  -56.3381,
  -56.3303,
  -56.3272,
  -56.3283,
  -56.3336,
  -56.3429,
  -56.3559,
  -56.3717,
  -56.3896,
  -56.409,
  -56.4295,
  -56.4501,
  -56.4698,
  -56.4876,
  -56.5026,
  -56.5138,
  -56.5203,
  -56.5211,
  -56.5164,
  -56.5064,
  -56.492,
  -56.4739,
  -56.4517,
  -56.428,
  -56.4028,
  -56.3767,
  -56.3495,
  -56.321,
  -56.2906,
  -56.2584,
  -56.2243,
  -56.1895,
  -56.1549,
  -56.1214,
  -56.0901,
  -56.0631,
  -56.0425,
  -56.0315,
  -56.0334,
  -56.0502,
  -56.0837,
  -45.069,
  -45.2634,
  -45.4548,
  -45.6458,
  -45.8392,
  -46.0368,
  -46.241,
  -46.4514,
  -46.6723,
  -46.9033,
  -47.1459,
  -47.4012,
  -47.67,
  -47.9504,
  -48.2441,
  -48.5479,
  -48.8607,
  -49.1813,
  -49.5072,
  -49.8361,
  -50.1652,
  -50.4932,
  -50.8186,
  -51.1424,
  -51.4623,
  -51.7779,
  -52.0908,
  -52.4011,
  -52.7093,
  -53.0156,
  -53.3197,
  -53.6201,
  -53.914,
  -54.1996,
  -54.4741,
  -54.7337,
  -54.9772,
  -55.2032,
  -55.4097,
  -55.5987,
  -55.7691,
  -55.9206,
  -56.0548,
  -56.1726,
  -56.2751,
  -56.3643,
  -56.4428,
  -56.5134,
  -56.5793,
  -56.644,
  -56.7104,
  -56.7805,
  -56.8551,
  -56.9338,
  -57.0142,
  -57.0967,
  -57.1783,
  -57.257,
  -57.3313,
  -57.4005,
  -57.4639,
  -57.5213,
  -57.5722,
  -57.6168,
  -57.6554,
  -57.6889,
  -57.7188,
  -57.7459,
  -57.7722,
  -57.7996,
  -57.8304,
  -57.8652,
  -57.9075,
  -57.9565,
  -58.0118,
  -58.074,
  -58.1427,
  -58.2173,
  -58.2982,
  -58.3875,
  -58.4866,
  -58.5987,
  -58.7254,
  -58.8688,
  -59.0292,
  -59.2064,
  -59.3997,
  -59.6069,
  -59.8286,
  -60.0598,
  -60.3012,
  -60.5483,
  -60.7978,
  -61.0454,
  -61.2868,
  -61.5175,
  -61.7331,
  -61.9292,
  -62.1024,
  -62.2502,
  -62.3716,
  -62.4668,
  -62.5372,
  -62.5862,
  -62.6175,
  -62.6346,
  -62.6417,
  -62.6416,
  -62.6398,
  -62.6381,
  -62.6391,
  -62.6448,
  -62.6565,
  -62.675,
  -62.701,
  -62.735,
  -62.7771,
  -62.8273,
  -62.8846,
  -62.948,
  -63.0163,
  -63.0885,
  -63.1636,
  -63.2409,
  -63.3201,
  -63.4011,
  -63.4833,
  -63.5657,
  -63.6497,
  -63.7338,
  -63.8176,
  -63.9007,
  -63.9829,
  -64.0637,
  -64.1426,
  -64.2194,
  -64.2932,
  -64.3643,
  -64.4324,
  -64.4969,
  -64.5574,
  -64.6129,
  -64.6631,
  -64.7072,
  -64.7442,
  -64.7732,
  -64.7929,
  -64.8033,
  -64.8039,
  -64.7937,
  -64.7755,
  -64.7483,
  -64.7137,
  -64.6728,
  -64.6272,
  -64.5784,
  -64.528,
  -64.4772,
  -64.4267,
  -64.3763,
  -64.3259,
  -64.2749,
  -64.2227,
  -64.169,
  -64.1133,
  -64.0558,
  -63.9971,
  -63.9384,
  -63.8809,
  -63.826,
  -63.7748,
  -63.7277,
  -63.6858,
  -63.6481,
  -63.6156,
  -63.5864,
  -63.5589,
  -63.5326,
  -63.5068,
  -63.4811,
  -63.4556,
  -63.43,
  -63.4048,
  -63.3797,
  -63.3539,
  -63.3267,
  -63.2964,
  -63.2632,
  -63.2263,
  -63.1851,
  -63.1392,
  -63.0879,
  -63.0325,
  -62.9735,
  -62.9109,
  -62.8457,
  -62.7771,
  -62.706,
  -62.6317,
  -62.552,
  -62.4677,
  -62.3766,
  -62.2787,
  -62.1735,
  -62.061,
  -61.9411,
  -61.8145,
  -61.6823,
  -61.545,
  -61.4031,
  -61.2563,
  -61.1041,
  -60.9476,
  -60.7872,
  -60.6236,
  -60.458,
  -60.2923,
  -60.1283,
  -59.9684,
  -59.8136,
  -59.6653,
  -59.524,
  -59.3895,
  -59.2607,
  -59.1368,
  -59.0164,
  -58.8981,
  -58.781,
  -58.6644,
  -58.5467,
  -58.43,
  -58.3131,
  -58.1956,
  -58.0779,
  -57.96,
  -57.8411,
  -57.7211,
  -57.6002,
  -57.4784,
  -57.3564,
  -57.2356,
  -57.117,
  -57.0021,
  -56.8918,
  -56.7867,
  -56.6878,
  -56.5958,
  -56.5108,
  -56.4333,
  -56.363,
  -56.2997,
  -56.2427,
  -56.1919,
  -56.1462,
  -56.1059,
  -56.0705,
  -56.0399,
  -56.0138,
  -55.9924,
  -55.9756,
  -55.9638,
  -55.9568,
  -55.9542,
  -55.9558,
  -55.9612,
  -55.9708,
  -55.9835,
  -56.0005,
  -56.0199,
  -56.0412,
  -56.0641,
  -56.0875,
  -56.1102,
  -56.1313,
  -56.1495,
  -56.1637,
  -56.173,
  -56.1767,
  -56.1748,
  -56.1675,
  -56.1557,
  -56.14,
  -56.1214,
  -56.1003,
  -56.0775,
  -56.0536,
  -56.0285,
  -56.002,
  -55.9728,
  -55.9411,
  -55.9069,
  -55.8714,
  -55.8356,
  -55.8001,
  -55.7668,
  -55.7373,
  -55.7142,
  -55.7009,
  -55.7008,
  -55.7166,
  -55.7499,
  -44.7205,
  -44.9113,
  -45.0985,
  -45.2872,
  -45.4797,
  -45.6773,
  -45.882,
  -46.0949,
  -46.3175,
  -46.5504,
  -46.795,
  -47.0521,
  -47.3224,
  -47.6048,
  -47.9,
  -48.2061,
  -48.5218,
  -48.8435,
  -49.1709,
  -49.5003,
  -49.8282,
  -50.1531,
  -50.4756,
  -50.7958,
  -51.1119,
  -51.424,
  -51.7335,
  -52.0409,
  -52.3467,
  -52.6512,
  -52.9542,
  -53.2534,
  -53.5457,
  -53.8292,
  -54.1006,
  -54.3565,
  -54.595,
  -54.8153,
  -55.017,
  -55.1998,
  -55.3642,
  -55.5104,
  -55.6398,
  -55.7534,
  -55.8534,
  -55.941,
  -56.0188,
  -56.0893,
  -56.1551,
  -56.2213,
  -56.2899,
  -56.3629,
  -56.4409,
  -56.5237,
  -56.6093,
  -56.6958,
  -56.7808,
  -56.8623,
  -56.9392,
  -57.0104,
  -57.0755,
  -57.134,
  -57.1859,
  -57.231,
  -57.2703,
  -57.3034,
  -57.3332,
  -57.3598,
  -57.3848,
  -57.4104,
  -57.4389,
  -57.4717,
  -57.51,
  -57.5549,
  -57.6062,
  -57.664,
  -57.7279,
  -57.7984,
  -57.8759,
  -57.9623,
  -58.0603,
  -58.1725,
  -58.2996,
  -58.4455,
  -58.6099,
  -58.7922,
  -58.9915,
  -59.2061,
  -59.435,
  -59.6745,
  -59.9229,
  -60.1763,
  -60.4319,
  -60.6856,
  -60.9324,
  -61.1681,
  -61.3882,
  -61.5887,
  -61.7661,
  -61.9175,
  -62.0421,
  -62.1386,
  -62.2104,
  -62.2599,
  -62.2907,
  -62.3066,
  -62.3117,
  -62.3098,
  -62.3047,
  -62.2997,
  -62.297,
  -62.299,
  -62.3067,
  -62.3212,
  -62.3437,
  -62.3747,
  -62.4144,
  -62.4624,
  -62.518,
  -62.5804,
  -62.647,
  -62.7186,
  -62.7931,
  -62.8697,
  -62.948,
  -63.0279,
  -63.1094,
  -63.192,
  -63.2751,
  -63.3584,
  -63.4414,
  -63.5244,
  -63.6065,
  -63.6879,
  -63.7678,
  -63.8458,
  -63.9216,
  -63.9947,
  -64.0649,
  -64.1313,
  -64.193,
  -64.2486,
  -64.299,
  -64.3427,
  -64.3783,
  -64.4048,
  -64.4217,
  -64.4282,
  -64.4242,
  -64.4099,
  -64.3858,
  -64.3528,
  -64.3119,
  -64.2646,
  -64.2126,
  -64.1575,
  -64.1013,
  -64.0445,
  -63.9882,
  -63.9322,
  -63.8762,
  -63.8199,
  -63.7625,
  -63.7037,
  -63.6423,
  -63.5805,
  -63.5185,
  -63.4571,
  -63.3975,
  -63.3413,
  -63.2893,
  -63.2425,
  -63.201,
  -63.1649,
  -63.1335,
  -63.1053,
  -63.0794,
  -63.0548,
  -63.0308,
  -63.0075,
  -62.9846,
  -62.9624,
  -62.9406,
  -62.9189,
  -62.8964,
  -62.8716,
  -62.8438,
  -62.8121,
  -62.7762,
  -62.7356,
  -62.6886,
  -62.638,
  -62.5828,
  -62.524,
  -62.4616,
  -62.3959,
  -62.3273,
  -62.2557,
  -62.1808,
  -62.1012,
  -62.0159,
  -61.9242,
  -61.8252,
  -61.7188,
  -61.605,
  -61.4837,
  -61.3554,
  -61.2211,
  -61.0812,
  -60.936,
  -60.7854,
  -60.6297,
  -60.4689,
  -60.3041,
  -60.1367,
  -59.9679,
  -59.8001,
  -59.6353,
  -59.4747,
  -59.3214,
  -59.1754,
  -59.0367,
  -58.9053,
  -58.7799,
  -58.6594,
  -58.5423,
  -58.4273,
  -58.3133,
  -58.1997,
  -58.0859,
  -57.9723,
  -57.8586,
  -57.7444,
  -57.6297,
  -57.5142,
  -57.398,
  -57.2805,
  -57.1618,
  -57.0426,
  -56.9236,
  -56.8065,
  -56.6921,
  -56.5815,
  -56.4758,
  -56.3756,
  -56.2817,
  -56.1942,
  -56.1132,
  -56.0388,
  -55.9709,
  -55.9095,
  -55.8539,
  -55.8029,
  -55.7586,
  -55.7193,
  -55.685,
  -55.6557,
  -55.6313,
  -55.6114,
  -55.596,
  -55.5851,
  -55.5786,
  -55.5764,
  -55.578,
  -55.5836,
  -55.5933,
  -55.6071,
  -55.625,
  -55.6459,
  -55.669,
  -55.6939,
  -55.7198,
  -55.7453,
  -55.769,
  -55.7898,
  -55.8066,
  -55.8184,
  -55.8244,
  -55.8248,
  -55.8201,
  -55.811,
  -55.7981,
  -55.7821,
  -55.7637,
  -55.7435,
  -55.7221,
  -55.6995,
  -55.6751,
  -55.6477,
  -55.6173,
  -55.5839,
  -55.5486,
  -55.5126,
  -55.4768,
  -55.4426,
  -55.412,
  -55.3867,
  -55.3722,
  -55.3708,
  -55.3857,
  -55.4188,
  -44.3728,
  -44.5601,
  -44.7455,
  -44.9324,
  -45.1239,
  -45.322,
  -45.5283,
  -45.7435,
  -45.9683,
  -46.2038,
  -46.4504,
  -46.7094,
  -46.9794,
  -47.2622,
  -47.5569,
  -47.8626,
  -48.1775,
  -48.4995,
  -48.8254,
  -49.1524,
  -49.4768,
  -49.7976,
  -50.1147,
  -50.4296,
  -50.7417,
  -51.0504,
  -51.3564,
  -51.6598,
  -51.9633,
  -52.2662,
  -52.5677,
  -52.8655,
  -53.1567,
  -53.4376,
  -53.7053,
  -53.9567,
  -54.19,
  -54.4047,
  -54.6005,
  -54.7779,
  -54.9371,
  -55.0791,
  -55.2045,
  -55.3165,
  -55.4152,
  -55.5026,
  -55.5809,
  -55.6528,
  -55.7212,
  -55.7895,
  -55.8604,
  -55.936,
  -56.0172,
  -56.1036,
  -56.193,
  -56.2828,
  -56.3711,
  -56.4556,
  -56.5349,
  -56.6076,
  -56.6751,
  -56.7356,
  -56.7895,
  -56.8369,
  -56.8785,
  -56.9147,
  -56.9461,
  -56.9742,
  -56.9999,
  -57.0256,
  -57.0532,
  -57.0849,
  -57.1211,
  -57.1638,
  -57.2119,
  -57.2669,
  -57.3261,
  -57.3936,
  -57.4683,
  -57.5522,
  -57.6487,
  -57.7602,
  -57.8891,
  -58.0367,
  -58.2038,
  -58.3908,
  -58.5954,
  -58.8162,
  -59.0508,
  -59.2962,
  -59.5496,
  -59.8076,
  -60.0673,
  -60.3242,
  -60.5732,
  -60.8118,
  -61.0345,
  -61.2373,
  -61.417,
  -61.5708,
  -61.6974,
  -61.7965,
  -61.8696,
  -61.92,
  -61.951,
  -61.9669,
  -61.9714,
  -61.9686,
  -61.9622,
  -61.9551,
  -61.9497,
  -61.9484,
  -61.9522,
  -61.9619,
  -61.9804,
  -62.0076,
  -62.0437,
  -62.0885,
  -62.1415,
  -62.2018,
  -62.2679,
  -62.3382,
  -62.4112,
  -62.4865,
  -62.5632,
  -62.6417,
  -62.7216,
  -62.8025,
  -62.8841,
  -62.9659,
  -63.0481,
  -63.1307,
  -63.2132,
  -63.2954,
  -63.3755,
  -63.4554,
  -63.5335,
  -63.6091,
  -63.6815,
  -63.7498,
  -63.8131,
  -63.8708,
  -63.9215,
  -63.9643,
  -63.9983,
  -64.0223,
  -64.0356,
  -64.0379,
  -64.0287,
  -64.0085,
  -63.9781,
  -63.9383,
  -63.8904,
  -63.8361,
  -63.7771,
  -63.7153,
  -63.6513,
  -63.588,
  -63.5254,
  -63.4631,
  -63.4013,
  -63.3392,
  -63.2763,
  -63.2122,
  -63.147,
  -63.0812,
  -63.0155,
  -62.9515,
  -62.8901,
  -62.8326,
  -62.7799,
  -62.7329,
  -62.6917,
  -62.6562,
  -62.6256,
  -62.5985,
  -62.5741,
  -62.5514,
  -62.5298,
  -62.509,
  -62.4885,
  -62.4702,
  -62.4528,
  -62.4351,
  -62.4159,
  -62.3943,
  -62.3688,
  -62.3389,
  -62.3038,
  -62.2634,
  -62.2177,
  -62.1673,
  -62.1127,
  -62.0543,
  -61.9922,
  -61.9268,
  -61.8586,
  -61.7869,
  -61.7115,
  -61.631,
  -61.5449,
  -61.4525,
  -61.3528,
  -61.2456,
  -61.1306,
  -61.0085,
  -60.8795,
  -60.7437,
  -60.6011,
  -60.4534,
  -60.2996,
  -60.1407,
  -59.9767,
  -59.8085,
  -59.6379,
  -59.4669,
  -59.2978,
  -59.1327,
  -58.9737,
  -58.8221,
  -58.6787,
  -58.5427,
  -58.4142,
  -58.2921,
  -58.1749,
  -58.0612,
  -57.9496,
  -57.8392,
  -57.729,
  -57.6189,
  -57.5088,
  -57.3985,
  -57.2881,
  -57.1767,
  -57.0646,
  -56.9513,
  -56.837,
  -56.7216,
  -56.6059,
  -56.4901,
  -56.3774,
  -56.2679,
  -56.1624,
  -56.062,
  -55.9668,
  -55.8775,
  -55.7943,
  -55.717,
  -55.6452,
  -55.5792,
  -55.5187,
  -55.4638,
  -55.4145,
  -55.3706,
  -55.3322,
  -55.2989,
  -55.2707,
  -55.2473,
  -55.2285,
  -55.2141,
  -55.2039,
  -55.1976,
  -55.1952,
  -55.1967,
  -55.2022,
  -55.212,
  -55.2261,
  -55.2446,
  -55.2671,
  -55.2922,
  -55.3193,
  -55.3474,
  -55.3753,
  -55.4015,
  -55.4245,
  -55.4433,
  -55.4569,
  -55.4649,
  -55.4675,
  -55.4642,
  -55.4576,
  -55.4473,
  -55.4341,
  -55.4183,
  -55.4008,
  -55.3821,
  -55.3623,
  -55.3405,
  -55.3158,
  -55.2873,
  -55.2556,
  -55.2218,
  -55.187,
  -55.1519,
  -55.1185,
  -55.0882,
  -55.064,
  -55.0494,
  -55.0476,
  -55.0621,
  -55.0948,
  -44.0312,
  -44.2153,
  -44.3984,
  -44.5837,
  -44.7747,
  -44.9739,
  -45.1819,
  -45.3987,
  -45.6264,
  -45.8644,
  -46.1131,
  -46.3726,
  -46.643,
  -46.9243,
  -47.2162,
  -47.5183,
  -47.8292,
  -48.147,
  -48.4687,
  -48.7907,
  -49.1097,
  -49.4237,
  -49.7352,
  -50.0443,
  -50.3507,
  -50.655,
  -50.9577,
  -51.259,
  -51.5602,
  -51.861,
  -52.1603,
  -52.4557,
  -52.7437,
  -53.021,
  -53.2847,
  -53.5314,
  -53.7599,
  -53.9686,
  -54.1595,
  -54.3324,
  -54.4881,
  -54.6275,
  -54.7527,
  -54.8646,
  -54.9643,
  -55.0531,
  -55.1333,
  -55.2072,
  -55.2782,
  -55.3488,
  -55.4222,
  -55.5006,
  -55.5845,
  -55.6728,
  -55.7652,
  -55.858,
  -55.9492,
  -56.0365,
  -56.1188,
  -56.1953,
  -56.2655,
  -56.3293,
  -56.3864,
  -56.4378,
  -56.4832,
  -56.523,
  -56.5583,
  -56.5896,
  -56.6187,
  -56.6467,
  -56.6753,
  -56.7073,
  -56.7447,
  -56.7874,
  -56.835,
  -56.8882,
  -56.9467,
  -57.0123,
  -57.0849,
  -57.168,
  -57.2632,
  -57.3731,
  -57.5006,
  -57.6484,
  -57.8175,
  -58.0066,
  -58.215,
  -58.4394,
  -58.6775,
  -58.9267,
  -59.1832,
  -59.4437,
  -59.7048,
  -59.9632,
  -60.2138,
  -60.4527,
  -60.6757,
  -60.8788,
  -61.0589,
  -61.2131,
  -61.3402,
  -61.44,
  -61.5141,
  -61.5655,
  -61.5975,
  -61.6144,
  -61.6189,
  -61.6169,
  -61.6107,
  -61.6032,
  -61.5963,
  -61.5921,
  -61.5927,
  -61.5995,
  -61.614,
  -61.6368,
  -61.6684,
  -61.709,
  -61.7584,
  -61.8156,
  -61.879,
  -61.9469,
  -62.018,
  -62.0911,
  -62.1658,
  -62.242,
  -62.3186,
  -62.3972,
  -62.4767,
  -62.5572,
  -62.6387,
  -62.7211,
  -62.8043,
  -62.8875,
  -62.9703,
  -63.0524,
  -63.133,
  -63.2111,
  -63.2859,
  -63.3562,
  -63.421,
  -63.4793,
  -63.53,
  -63.5718,
  -63.6037,
  -63.6246,
  -63.6339,
  -63.6312,
  -63.6153,
  -63.5889,
  -63.5515,
  -63.5045,
  -63.4491,
  -63.3871,
  -63.3205,
  -63.2511,
  -63.1807,
  -63.1105,
  -63.041,
  -62.9722,
  -62.9039,
  -62.8359,
  -62.7675,
  -62.6981,
  -62.6283,
  -62.5584,
  -62.4895,
  -62.4229,
  -62.3598,
  -62.3011,
  -62.2478,
  -62.1994,
  -62.1582,
  -62.1229,
  -62.0926,
  -62.0667,
  -62.0437,
  -62.0229,
  -62.004,
  -61.9867,
  -61.9711,
  -61.9574,
  -61.9444,
  -61.9314,
  -61.9163,
  -61.8978,
  -61.8751,
  -61.8467,
  -61.8125,
  -61.7724,
  -61.727,
  -61.6769,
  -61.6226,
  -61.5648,
  -61.5033,
  -61.4385,
  -61.3708,
  -61.2995,
  -61.2228,
  -61.1419,
  -61.0553,
  -60.9623,
  -60.862,
  -60.7544,
  -60.639,
  -60.5167,
  -60.3874,
  -60.2515,
  -60.1088,
  -59.9598,
  -59.8044,
  -59.6435,
  -59.4773,
  -59.3072,
  -59.135,
  -58.9629,
  -58.7933,
  -58.6285,
  -58.4704,
  -58.3204,
  -58.1792,
  -58.046,
  -57.9201,
  -57.8007,
  -57.6867,
  -57.5764,
  -57.4683,
  -57.3616,
  -57.2542,
  -57.148,
  -57.0415,
  -56.935,
  -56.8281,
  -56.7204,
  -56.6117,
  -56.502,
  -56.3913,
  -56.2802,
  -56.169,
  -56.0591,
  -55.9516,
  -55.8476,
  -55.748,
  -55.653,
  -55.5629,
  -55.4781,
  -55.3984,
  -55.3239,
  -55.2542,
  -55.1894,
  -55.1294,
  -55.0747,
  -55.0255,
  -54.982,
  -54.9443,
  -54.9118,
  -54.8843,
  -54.8617,
  -54.8434,
  -54.8294,
  -54.8191,
  -54.8126,
  -54.8098,
  -54.811,
  -54.8153,
  -54.8252,
  -54.8399,
  -54.8594,
  -54.8833,
  -54.9107,
  -54.9402,
  -54.9705,
  -55.0006,
  -55.0289,
  -55.0538,
  -55.0741,
  -55.0891,
  -55.0989,
  -55.1034,
  -55.1033,
  -55.0992,
  -55.0916,
  -55.0808,
  -55.0678,
  -55.053,
  -55.0371,
  -55.0203,
  -55.0015,
  -54.9796,
  -54.9542,
  -54.9255,
  -54.8945,
  -54.8621,
  -54.8295,
  -54.7978,
  -54.7694,
  -54.7467,
  -54.733,
  -54.7317,
  -54.7459,
  -54.778,
  -43.6974,
  -43.8786,
  -44.0589,
  -44.2432,
  -44.434,
  -44.6339,
  -44.8435,
  -45.0636,
  -45.2939,
  -45.5336,
  -45.7831,
  -46.0416,
  -46.3099,
  -46.5873,
  -46.8737,
  -47.1694,
  -47.473,
  -47.784,
  -48.099,
  -48.4142,
  -48.7262,
  -49.0347,
  -49.3395,
  -49.6425,
  -49.9432,
  -50.2427,
  -50.5407,
  -50.8385,
  -51.1364,
  -51.4344,
  -51.7304,
  -52.0212,
  -52.3051,
  -52.5781,
  -52.8369,
  -53.0793,
  -53.3034,
  -53.5089,
  -53.6964,
  -53.8663,
  -54.0198,
  -54.1586,
  -54.2843,
  -54.3977,
  -54.4997,
  -54.5913,
  -54.6746,
  -54.7508,
  -54.8249,
  -54.8985,
  -54.9747,
  -55.0556,
  -55.1421,
  -55.2336,
  -55.3283,
  -55.4236,
  -55.5173,
  -55.6072,
  -55.6926,
  -55.7724,
  -55.8464,
  -55.914,
  -55.9761,
  -56.0323,
  -56.082,
  -56.1278,
  -56.1688,
  -56.2061,
  -56.2403,
  -56.2734,
  -56.3068,
  -56.3435,
  -56.3838,
  -56.4289,
  -56.4786,
  -56.5327,
  -56.5921,
  -56.6577,
  -56.7308,
  -56.8132,
  -56.9074,
  -57.0155,
  -57.1421,
  -57.2889,
  -57.4568,
  -57.6466,
  -57.8552,
  -58.0811,
  -58.3206,
  -58.5706,
  -58.828,
  -59.0882,
  -59.349,
  -59.6061,
  -59.8553,
  -60.0925,
  -60.3134,
  -60.5146,
  -60.6926,
  -60.8453,
  -60.9702,
  -61.0694,
  -61.1436,
  -61.1958,
  -61.2292,
  -61.248,
  -61.2558,
  -61.2559,
  -61.2515,
  -61.2447,
  -61.2374,
  -61.2318,
  -61.2297,
  -61.2332,
  -61.2436,
  -61.2618,
  -61.2885,
  -61.3241,
  -61.3688,
  -61.4209,
  -61.4804,
  -61.545,
  -61.6129,
  -61.6833,
  -61.7556,
  -61.8289,
  -61.9035,
  -61.9794,
  -62.0569,
  -62.1361,
  -62.2171,
  -62.3,
  -62.3842,
  -62.4691,
  -62.5541,
  -62.6386,
  -62.7216,
  -62.8021,
  -62.879,
  -62.9512,
  -63.0159,
  -63.0743,
  -63.124,
  -63.1642,
  -63.1934,
  -63.2107,
  -63.2155,
  -63.2073,
  -63.1865,
  -63.1533,
  -63.1087,
  -63.0538,
  -62.9902,
  -62.92,
  -62.8452,
  -62.7679,
  -62.6897,
  -62.6119,
  -62.5352,
  -62.4594,
  -62.3851,
  -62.3111,
  -62.2371,
  -62.162,
  -62.0877,
  -62.0143,
  -61.9425,
  -61.8736,
  -61.8087,
  -61.7491,
  -61.695,
  -61.6472,
  -61.6056,
  -61.5702,
  -61.5401,
  -61.5147,
  -61.493,
  -61.4742,
  -61.4581,
  -61.4447,
  -61.434,
  -61.4251,
  -61.4173,
  -61.409,
  -61.3984,
  -61.3835,
  -61.363,
  -61.3363,
  -61.3022,
  -61.2627,
  -61.2175,
  -61.1675,
  -61.1134,
  -61.0559,
  -60.9955,
  -60.9317,
  -60.8646,
  -60.7936,
  -60.718,
  -60.6371,
  -60.5501,
  -60.4568,
  -60.3563,
  -60.2487,
  -60.1338,
  -60.0118,
  -59.8832,
  -59.7479,
  -59.6059,
  -59.4569,
  -59.3016,
  -59.1403,
  -58.9738,
  -58.8034,
  -58.6313,
  -58.4595,
  -58.2893,
  -58.1255,
  -57.9688,
  -57.8206,
  -57.681,
  -57.55,
  -57.4265,
  -57.3095,
  -57.1981,
  -57.0908,
  -56.9859,
  -56.8827,
  -56.78,
  -56.6774,
  -56.5747,
  -56.4718,
  -56.3682,
  -56.264,
  -56.159,
  -56.0531,
  -55.9466,
  -55.8401,
  -55.7341,
  -55.6298,
  -55.5282,
  -55.4303,
  -55.3366,
  -55.2473,
  -55.1622,
  -55.0815,
  -55.0048,
  -54.9323,
  -54.864,
  -54.7998,
  -54.7393,
  -54.6846,
  -54.6355,
  -54.5922,
  -54.5547,
  -54.5229,
  -54.496,
  -54.4736,
  -54.4553,
  -54.4408,
  -54.4301,
  -54.423,
  -54.4195,
  -54.4201,
  -54.4251,
  -54.4353,
  -54.4509,
  -54.4718,
  -54.4976,
  -54.5273,
  -54.5595,
  -54.5922,
  -54.6242,
  -54.6543,
  -54.6808,
  -54.7023,
  -54.7185,
  -54.7295,
  -54.7358,
  -54.7378,
  -54.736,
  -54.7309,
  -54.7228,
  -54.7124,
  -54.7005,
  -54.6878,
  -54.674,
  -54.6584,
  -54.6401,
  -54.6185,
  -54.5939,
  -54.5667,
  -54.5381,
  -54.5079,
  -54.4797,
  -54.4541,
  -54.4339,
  -54.422,
  -54.4218,
  -54.4363,
  -54.4676,
  -43.3718,
  -43.5502,
  -43.73,
  -43.9137,
  -44.104,
  -44.3041,
  -44.5149,
  -44.7363,
  -44.9676,
  -45.208,
  -45.4564,
  -45.7113,
  -45.975,
  -46.246,
  -46.5247,
  -46.8121,
  -47.108,
  -47.4104,
  -47.7168,
  -48.0241,
  -48.3287,
  -48.6297,
  -48.9276,
  -49.2241,
  -49.5186,
  -49.8127,
  -50.1049,
  -50.3983,
  -50.6921,
  -50.9859,
  -51.2777,
  -51.5647,
  -51.8436,
  -52.111,
  -52.365,
  -52.603,
  -52.8231,
  -53.0255,
  -53.2104,
  -53.3787,
  -53.5319,
  -53.6716,
  -53.7981,
  -53.9142,
  -54.0195,
  -54.1151,
  -54.2025,
  -54.2838,
  -54.3616,
  -54.4386,
  -54.5179,
  -54.6016,
  -54.6903,
  -54.7837,
  -54.8802,
  -54.9776,
  -55.0735,
  -55.1663,
  -55.254,
  -55.3375,
  -55.4158,
  -55.4887,
  -55.5562,
  -55.6187,
  -55.6762,
  -55.7295,
  -55.7783,
  -55.8233,
  -55.8651,
  -55.9051,
  -55.9455,
  -55.9882,
  -56.0346,
  -56.0849,
  -56.1392,
  -56.1966,
  -56.2594,
  -56.3282,
  -56.4039,
  -56.4879,
  -56.583,
  -56.6913,
  -56.8167,
  -56.9613,
  -57.1272,
  -57.3139,
  -57.5204,
  -57.7445,
  -57.982,
  -58.2301,
  -58.485,
  -58.7431,
  -59.0008,
  -59.2538,
  -59.4994,
  -59.7324,
  -59.9494,
  -60.1462,
  -60.3198,
  -60.4686,
  -60.5912,
  -60.6884,
  -60.7617,
  -60.8138,
  -60.8484,
  -60.8695,
  -60.8803,
  -60.8836,
  -60.8818,
  -60.8768,
  -60.8704,
  -60.8644,
  -60.8598,
  -60.8608,
  -60.8674,
  -60.8809,
  -60.9025,
  -60.933,
  -60.9723,
  -61.02,
  -61.0746,
  -61.1349,
  -61.1991,
  -61.266,
  -61.3347,
  -61.4048,
  -61.4765,
  -61.5499,
  -61.6257,
  -61.7039,
  -61.7852,
  -61.8691,
  -61.9541,
  -62.0413,
  -62.1287,
  -62.2154,
  -62.3007,
  -62.3833,
  -62.4617,
  -62.5346,
  -62.6005,
  -62.6583,
  -62.7065,
  -62.7439,
  -62.7696,
  -62.7825,
  -62.7823,
  -62.7684,
  -62.7411,
  -62.7008,
  -62.6485,
  -62.5855,
  -62.5136,
  -62.4349,
  -62.3517,
  -62.2652,
  -62.1789,
  -62.0932,
  -62.009,
  -61.9266,
  -61.8457,
  -61.766,
  -61.687,
  -61.6084,
  -61.5305,
  -61.454,
  -61.3798,
  -61.3092,
  -61.2429,
  -61.1822,
  -61.1276,
  -61.0793,
  -61.0371,
  -61.0011,
  -60.9708,
  -60.9457,
  -60.9249,
  -60.908,
  -60.8952,
  -60.8849,
  -60.8788,
  -60.8753,
  -60.8729,
  -60.8696,
  -60.8632,
  -60.852,
  -60.8343,
  -60.8094,
  -60.7773,
  -60.7383,
  -60.6933,
  -60.6435,
  -60.5896,
  -60.5326,
  -60.4726,
  -60.4096,
  -60.3434,
  -60.273,
  -60.1978,
  -60.1168,
  -60.0299,
  -59.9366,
  -59.8366,
  -59.7296,
  -59.6155,
  -59.4949,
  -59.3669,
  -59.2335,
  -59.0934,
  -58.9464,
  -58.7928,
  -58.6331,
  -58.4682,
  -58.2996,
  -58.129,
  -57.9589,
  -57.7915,
  -57.6295,
  -57.4747,
  -57.328,
  -57.19,
  -57.0604,
  -56.9389,
  -56.8238,
  -56.7145,
  -56.6094,
  -56.5073,
  -56.4071,
  -56.3075,
  -56.2083,
  -56.1089,
  -56.0091,
  -55.9087,
  -55.8077,
  -55.7063,
  -55.604,
  -55.5017,
  -55.3989,
  -55.2984,
  -55.2002,
  -55.1049,
  -55.0132,
  -54.9251,
  -54.8411,
  -54.7611,
  -54.6844,
  -54.6105,
  -54.5397,
  -54.4724,
  -54.4089,
  -54.3497,
  -54.2953,
  -54.2464,
  -54.2032,
  -54.1662,
  -54.1346,
  -54.108,
  -54.0855,
  -54.0667,
  -54.0513,
  -54.0395,
  -54.0312,
  -54.0268,
  -54.0266,
  -54.0314,
  -54.0419,
  -54.0587,
  -54.0813,
  -54.1091,
  -54.1413,
  -54.1761,
  -54.2114,
  -54.2455,
  -54.2771,
  -54.3047,
  -54.3274,
  -54.3437,
  -54.3559,
  -54.3637,
  -54.3675,
  -54.3679,
  -54.3653,
  -54.3601,
  -54.3527,
  -54.3442,
  -54.3347,
  -54.3244,
  -54.3125,
  -54.298,
  -54.2808,
  -54.2606,
  -54.238,
  -54.2138,
  -54.1892,
  -54.1653,
  -54.1437,
  -54.1268,
  -54.1174,
  -54.1188,
  -54.1335,
  -54.1641,
  -43.0556,
  -43.232,
  -43.4101,
  -43.593,
  -43.7829,
  -43.9826,
  -44.1921,
  -44.4134,
  -44.6442,
  -44.8828,
  -45.128,
  -45.3791,
  -45.6361,
  -45.8988,
  -46.1683,
  -46.4458,
  -46.7314,
  -47.0241,
  -47.3209,
  -47.6198,
  -47.9168,
  -48.2095,
  -48.5003,
  -48.7895,
  -49.0785,
  -49.3667,
  -49.6547,
  -49.9429,
  -50.2317,
  -50.52,
  -50.8058,
  -51.0868,
  -51.3595,
  -51.6213,
  -51.8698,
  -52.1032,
  -52.3189,
  -52.5187,
  -52.7021,
  -52.8701,
  -53.0242,
  -53.1657,
  -53.2957,
  -53.4152,
  -53.5246,
  -53.6246,
  -53.7167,
  -53.8027,
  -53.885,
  -53.9659,
  -54.0489,
  -54.1354,
  -54.2252,
  -54.3203,
  -54.4184,
  -54.5176,
  -54.6158,
  -54.7113,
  -54.8033,
  -54.8911,
  -54.9745,
  -55.0531,
  -55.1268,
  -55.1964,
  -55.2621,
  -55.3242,
  -55.3825,
  -55.4366,
  -55.4873,
  -55.5354,
  -55.5843,
  -55.6359,
  -55.6907,
  -55.7489,
  -55.8103,
  -55.8756,
  -55.9453,
  -56.02,
  -56.1006,
  -56.1897,
  -56.2874,
  -56.3967,
  -56.5221,
  -56.6645,
  -56.8269,
  -57.0092,
  -57.2102,
  -57.4283,
  -57.661,
  -57.9043,
  -58.155,
  -58.4087,
  -58.6616,
  -58.9104,
  -59.1503,
  -59.3774,
  -59.588,
  -59.7784,
  -59.9454,
  -60.0879,
  -60.2054,
  -60.2983,
  -60.369,
  -60.4199,
  -60.4552,
  -60.4773,
  -60.4912,
  -60.4978,
  -60.499,
  -60.4967,
  -60.4923,
  -60.4869,
  -60.4833,
  -60.4823,
  -60.4856,
  -60.4952,
  -60.512,
  -60.5371,
  -60.5706,
  -60.6124,
  -60.6617,
  -60.7168,
  -60.7766,
  -60.8392,
  -60.904,
  -60.9698,
  -61.0386,
  -61.1097,
  -61.1839,
  -61.2619,
  -61.3441,
  -61.4298,
  -61.518,
  -61.6077,
  -61.6979,
  -61.7871,
  -61.8743,
  -61.9582,
  -62.0371,
  -62.1099,
  -62.1751,
  -62.231,
  -62.2766,
  -62.3103,
  -62.3315,
  -62.3392,
  -62.333,
  -62.3119,
  -62.2778,
  -62.2302,
  -62.1702,
  -62.0991,
  -62.0189,
  -61.9319,
  -61.8404,
  -61.7464,
  -61.652,
  -61.5584,
  -61.4669,
  -61.3777,
  -61.2908,
  -61.2057,
  -61.122,
  -61.0398,
  -60.9588,
  -60.88,
  -60.8041,
  -60.7321,
  -60.6652,
  -60.604,
  -60.5479,
  -60.4989,
  -60.4562,
  -60.4198,
  -60.3891,
  -60.3638,
  -60.3437,
  -60.3285,
  -60.3186,
  -60.3132,
  -60.3121,
  -60.3138,
  -60.3167,
  -60.3181,
  -60.3159,
  -60.3081,
  -60.2931,
  -60.2702,
  -60.239,
  -60.2006,
  -60.1559,
  -60.1062,
  -60.0524,
  -59.9953,
  -59.9358,
  -59.8736,
  -59.807,
  -59.7373,
  -59.6623,
  -59.5819,
  -59.4955,
  -59.4028,
  -59.3035,
  -59.1978,
  -59.0857,
  -58.9673,
  -58.8429,
  -58.7124,
  -58.5757,
  -58.4322,
  -58.282,
  -58.1259,
  -57.9645,
  -57.7995,
  -57.6326,
  -57.4656,
  -57.3012,
  -57.1417,
  -56.9891,
  -56.8443,
  -56.7076,
  -56.5792,
  -56.4584,
  -56.3448,
  -56.2369,
  -56.1334,
  -56.0324,
  -55.9344,
  -55.8375,
  -55.7409,
  -55.6442,
  -55.5471,
  -55.4491,
  -55.3511,
  -55.2528,
  -55.1539,
  -55.0554,
  -54.9581,
  -54.863,
  -54.7706,
  -54.6813,
  -54.5955,
  -54.5133,
  -54.4347,
  -54.3593,
  -54.2863,
  -54.2153,
  -54.1463,
  -54.0802,
  -54.0175,
  -53.9588,
  -53.9052,
  -53.8569,
  -53.8144,
  -53.7775,
  -53.7461,
  -53.7194,
  -53.6965,
  -53.677,
  -53.6603,
  -53.6469,
  -53.636,
  -53.6302,
  -53.6293,
  -53.6338,
  -53.6448,
  -53.6628,
  -53.6873,
  -53.7175,
  -53.7521,
  -53.7894,
  -53.8272,
  -53.8634,
  -53.8962,
  -53.9247,
  -53.9483,
  -53.9668,
  -53.9802,
  -53.9894,
  -53.9951,
  -53.9979,
  -53.998,
  -53.9959,
  -53.9921,
  -53.9871,
  -53.9814,
  -53.9747,
  -53.9667,
  -53.9565,
  -53.9438,
  -53.9283,
  -53.9106,
  -53.8912,
  -53.8714,
  -53.8522,
  -53.8352,
  -53.8223,
  -53.8161,
  -53.8195,
  -53.8348,
  -53.8644,
  -42.7452,
  -42.9189,
  -43.0957,
  -43.2776,
  -43.4667,
  -43.6652,
  -43.8745,
  -44.0938,
  -44.3221,
  -44.5568,
  -44.7969,
  -45.0411,
  -45.2896,
  -45.543,
  -45.8024,
  -46.0679,
  -46.3423,
  -46.6239,
  -46.9105,
  -47.1997,
  -47.4881,
  -47.7746,
  -48.0588,
  -48.3424,
  -48.6263,
  -48.9091,
  -49.1914,
  -49.4742,
  -49.757,
  -50.0389,
  -50.318,
  -50.5908,
  -50.8565,
  -51.1115,
  -51.3541,
  -51.5827,
  -51.7956,
  -51.9933,
  -52.1758,
  -52.344,
  -52.4992,
  -52.6428,
  -52.776,
  -52.8991,
  -53.0125,
  -53.1171,
  -53.2131,
  -53.304,
  -53.3911,
  -53.4767,
  -53.5634,
  -53.6526,
  -53.7458,
  -53.8432,
  -53.9431,
  -54.0444,
  -54.145,
  -54.2436,
  -54.3393,
  -54.4318,
  -54.5205,
  -54.605,
  -54.6856,
  -54.762,
  -54.8363,
  -54.9075,
  -54.9754,
  -55.0392,
  -55.1003,
  -55.1594,
  -55.2191,
  -55.2811,
  -55.3459,
  -55.4138,
  -55.4852,
  -55.56,
  -55.6388,
  -55.722,
  -55.811,
  -55.907,
  -56.0098,
  -56.1227,
  -56.2486,
  -56.3907,
  -56.5507,
  -56.728,
  -56.9239,
  -57.1364,
  -57.3623,
  -57.5985,
  -57.8417,
  -58.089,
  -58.3356,
  -58.5771,
  -58.8099,
  -59.0293,
  -59.2316,
  -59.4132,
  -59.5706,
  -59.7049,
  -59.8147,
  -59.9013,
  -59.9673,
  -60.0157,
  -60.0503,
  -60.0744,
  -60.0903,
  -60.0998,
  -60.1045,
  -60.1052,
  -60.1033,
  -60.0998,
  -60.0963,
  -60.0945,
  -60.0957,
  -60.102,
  -60.1147,
  -60.1349,
  -60.162,
  -60.1979,
  -60.2416,
  -60.2914,
  -60.346,
  -60.4038,
  -60.4642,
  -60.5273,
  -60.5933,
  -60.6626,
  -60.7359,
  -60.8142,
  -60.8977,
  -60.9855,
  -61.0764,
  -61.1688,
  -61.2619,
  -61.3533,
  -61.4421,
  -61.5264,
  -61.605,
  -61.6754,
  -61.7383,
  -61.7911,
  -61.8327,
  -61.8618,
  -61.8776,
  -61.8795,
  -61.8672,
  -61.8403,
  -61.7991,
  -61.7444,
  -61.6769,
  -61.5978,
  -61.5097,
  -61.4144,
  -61.3147,
  -61.2127,
  -61.1103,
  -61.0094,
  -60.9107,
  -60.8151,
  -60.7224,
  -60.6314,
  -60.5439,
  -60.4588,
  -60.3758,
  -60.2955,
  -60.2186,
  -60.1461,
  -60.0791,
  -60.0176,
  -59.9622,
  -59.9126,
  -59.8694,
  -59.8324,
  -59.8011,
  -59.7756,
  -59.7561,
  -59.7428,
  -59.7354,
  -59.7336,
  -59.7365,
  -59.7431,
  -59.7507,
  -59.7567,
  -59.7584,
  -59.7538,
  -59.7404,
  -59.719,
  -59.6887,
  -59.6508,
  -59.6063,
  -59.5564,
  -59.5025,
  -59.4457,
  -59.3864,
  -59.3247,
  -59.2594,
  -59.1899,
  -59.1157,
  -59.0361,
  -58.9507,
  -58.8592,
  -58.7615,
  -58.658,
  -58.5486,
  -58.4336,
  -58.313,
  -58.1866,
  -58.0542,
  -57.9153,
  -57.7701,
  -57.6189,
  -57.4625,
  -57.3023,
  -57.1402,
  -56.9771,
  -56.8165,
  -56.6606,
  -56.5111,
  -56.3684,
  -56.2332,
  -56.1058,
  -55.9858,
  -55.8729,
  -55.7659,
  -55.6637,
  -55.5648,
  -55.4683,
  -55.3732,
  -55.2787,
  -55.1838,
  -55.0886,
  -54.9931,
  -54.8973,
  -54.8012,
  -54.7051,
  -54.6095,
  -54.5161,
  -54.4254,
  -54.3378,
  -54.2537,
  -54.1733,
  -54.0965,
  -54.0229,
  -53.952,
  -53.8827,
  -53.815,
  -53.7488,
  -53.6836,
  -53.6223,
  -53.565,
  -53.5126,
  -53.4658,
  -53.4243,
  -53.3881,
  -53.357,
  -53.3299,
  -53.3064,
  -53.2856,
  -53.2674,
  -53.252,
  -53.2402,
  -53.2328,
  -53.2309,
  -53.2352,
  -53.2465,
  -53.2656,
  -53.2919,
  -53.3246,
  -53.3617,
  -53.4013,
  -53.4412,
  -53.4792,
  -53.5134,
  -53.5429,
  -53.5672,
  -53.5866,
  -53.6012,
  -53.6118,
  -53.6196,
  -53.6251,
  -53.6286,
  -53.6302,
  -53.6303,
  -53.6295,
  -53.6278,
  -53.6252,
  -53.6214,
  -53.6154,
  -53.607,
  -53.5952,
  -53.5822,
  -53.5679,
  -53.5531,
  -53.5389,
  -53.5267,
  -53.5181,
  -53.5152,
  -53.5204,
  -53.5363,
  -53.5649,
  -42.4369,
  -42.6117,
  -42.7871,
  -42.9671,
  -43.1549,
  -43.3518,
  -43.5584,
  -43.7744,
  -43.9982,
  -44.2273,
  -44.4596,
  -44.6958,
  -44.9348,
  -45.1779,
  -45.4264,
  -45.6816,
  -45.9441,
  -46.2141,
  -46.4898,
  -46.7693,
  -47.0496,
  -47.3288,
  -47.6073,
  -47.8854,
  -48.1635,
  -48.4403,
  -48.7174,
  -48.9941,
  -49.2704,
  -49.5451,
  -49.8162,
  -50.0822,
  -50.34,
  -50.5879,
  -50.8241,
  -51.0476,
  -51.2573,
  -51.4524,
  -51.6339,
  -51.8022,
  -51.9587,
  -52.1031,
  -52.2387,
  -52.3648,
  -52.4821,
  -52.591,
  -52.6925,
  -52.7885,
  -52.8806,
  -52.971,
  -53.0614,
  -53.1543,
  -53.2504,
  -53.3501,
  -53.4525,
  -53.5561,
  -53.6595,
  -53.7604,
  -53.86,
  -53.9572,
  -54.0511,
  -54.142,
  -54.2298,
  -54.3151,
  -54.3982,
  -54.4786,
  -54.5557,
  -54.6297,
  -54.7011,
  -54.7714,
  -54.8426,
  -54.9155,
  -54.9917,
  -55.0712,
  -55.1528,
  -55.2391,
  -55.3294,
  -55.4241,
  -55.5235,
  -55.6286,
  -55.7398,
  -55.8595,
  -55.99,
  -56.1336,
  -56.2916,
  -56.4651,
  -56.6559,
  -56.8615,
  -57.0799,
  -57.3084,
  -57.544,
  -57.7829,
  -58.0204,
  -58.254,
  -58.4783,
  -58.6884,
  -58.8808,
  -59.0522,
  -59.2001,
  -59.324,
  -59.4241,
  -59.5024,
  -59.5618,
  -59.6058,
  -59.638,
  -59.6612,
  -59.6781,
  -59.6897,
  -59.6969,
  -59.7007,
  -59.7015,
  -59.6992,
  -59.6971,
  -59.6951,
  -59.6952,
  -59.6992,
  -59.7085,
  -59.7244,
  -59.7475,
  -59.7784,
  -59.8164,
  -59.8607,
  -59.9098,
  -59.9626,
  -60.0188,
  -60.0783,
  -60.1417,
  -60.2095,
  -60.2823,
  -60.3612,
  -60.4461,
  -60.5351,
  -60.6287,
  -60.7241,
  -60.8197,
  -60.9131,
  -61.0026,
  -61.0866,
  -61.1637,
  -61.2325,
  -61.2917,
  -61.3401,
  -61.3766,
  -61.4001,
  -61.4099,
  -61.4053,
  -61.3863,
  -61.3526,
  -61.3046,
  -61.2427,
  -61.1677,
  -61.0813,
  -60.9858,
  -60.8821,
  -60.7751,
  -60.6656,
  -60.556,
  -60.4479,
  -60.3428,
  -60.2412,
  -60.1433,
  -60.0491,
  -59.9583,
  -59.871,
  -59.7868,
  -59.706,
  -59.6291,
  -59.5569,
  -59.4902,
  -59.4291,
  -59.3736,
  -59.324,
  -59.2804,
  -59.2429,
  -59.2113,
  -59.1858,
  -59.1667,
  -59.1536,
  -59.1481,
  -59.1492,
  -59.1558,
  -59.1661,
  -59.1777,
  -59.1876,
  -59.1928,
  -59.1907,
  -59.1802,
  -59.1601,
  -59.1307,
  -59.093,
  -59.0483,
  -58.9982,
  -58.9442,
  -58.8873,
  -58.8282,
  -58.7665,
  -58.7017,
  -58.6329,
  -58.5594,
  -58.481,
  -58.3973,
  -58.3076,
  -58.2125,
  -58.1121,
  -58.0057,
  -57.8949,
  -57.7789,
  -57.6574,
  -57.5304,
  -57.3972,
  -57.2578,
  -57.1124,
  -56.9622,
  -56.8081,
  -56.6517,
  -56.495,
  -56.3399,
  -56.1881,
  -56.0419,
  -55.9019,
  -55.7684,
  -55.6418,
  -55.5226,
  -55.4103,
  -55.304,
  -55.2022,
  -55.1041,
  -55.0087,
  -54.9147,
  -54.8212,
  -54.7279,
  -54.634,
  -54.54,
  -54.4457,
  -54.3511,
  -54.2559,
  -54.1628,
  -54.0721,
  -53.9849,
  -53.9011,
  -53.8211,
  -53.7449,
  -53.6729,
  -53.6039,
  -53.537,
  -53.4717,
  -53.4074,
  -53.3444,
  -53.2832,
  -53.2244,
  -53.1693,
  -53.1186,
  -53.0738,
  -53.0341,
  -52.999,
  -52.9681,
  -52.9407,
  -52.9163,
  -52.8943,
  -52.8744,
  -52.857,
  -52.8432,
  -52.8341,
  -52.8311,
  -52.835,
  -52.8468,
  -52.867,
  -52.895,
  -52.9297,
  -52.9691,
  -53.0107,
  -53.0524,
  -53.092,
  -53.1274,
  -53.1566,
  -53.1817,
  -53.2017,
  -53.2175,
  -53.2299,
  -53.24,
  -53.2486,
  -53.256,
  -53.262,
  -53.2668,
  -53.2704,
  -53.2732,
  -53.2751,
  -53.2752,
  -53.2734,
  -53.2691,
  -53.2627,
  -53.2544,
  -53.2449,
  -53.235,
  -53.2259,
  -53.2185,
  -53.2142,
  -53.2148,
  -53.2223,
  -53.2388,
  -53.266,
  -42.132,
  -42.3061,
  -42.4807,
  -42.6593,
  -42.8449,
  -43.038,
  -43.2411,
  -43.4526,
  -43.6704,
  -43.8924,
  -44.1178,
  -44.3454,
  -44.5746,
  -44.8072,
  -45.045,
  -45.2886,
  -45.5393,
  -45.7978,
  -46.0623,
  -46.3314,
  -46.6023,
  -46.8753,
  -47.148,
  -47.421,
  -47.6938,
  -47.9661,
  -48.2375,
  -48.5082,
  -48.7773,
  -49.044,
  -49.3069,
  -49.5648,
  -49.8146,
  -50.0543,
  -50.2846,
  -50.5013,
  -50.7069,
  -50.9002,
  -51.0801,
  -51.2476,
  -51.4046,
  -51.5512,
  -51.6886,
  -51.8169,
  -51.937,
  -52.0493,
  -52.155,
  -52.2555,
  -52.3525,
  -52.4475,
  -52.5424,
  -52.6381,
  -52.7377,
  -52.8404,
  -52.9453,
  -53.0518,
  -53.158,
  -53.2634,
  -53.3671,
  -53.4689,
  -53.5685,
  -53.6657,
  -53.7608,
  -53.854,
  -53.9454,
  -54.0344,
  -54.1207,
  -54.2045,
  -54.2853,
  -54.3663,
  -54.4489,
  -54.5335,
  -54.6217,
  -54.7129,
  -54.8079,
  -54.9071,
  -55.0107,
  -55.1182,
  -55.2299,
  -55.3461,
  -55.4678,
  -55.5965,
  -55.7335,
  -55.8803,
  -56.0386,
  -56.2096,
  -56.3967,
  -56.5972,
  -56.8083,
  -57.0294,
  -57.2571,
  -57.4877,
  -57.7177,
  -57.9424,
  -58.1572,
  -58.3573,
  -58.5388,
  -58.6986,
  -58.8346,
  -58.9466,
  -59.0356,
  -59.1039,
  -59.1548,
  -59.1924,
  -59.2191,
  -59.2396,
  -59.2558,
  -59.2682,
  -59.277,
  -59.2831,
  -59.2863,
  -59.2874,
  -59.2865,
  -59.2854,
  -59.2853,
  -59.2877,
  -59.2946,
  -59.3069,
  -59.326,
  -59.3522,
  -59.3853,
  -59.4241,
  -59.4679,
  -59.5159,
  -59.5667,
  -59.6228,
  -59.6837,
  -59.7501,
  -59.8229,
  -59.9027,
  -59.9892,
  -60.0813,
  -60.1774,
  -60.2751,
  -60.3726,
  -60.4671,
  -60.5568,
  -60.6394,
  -60.7138,
  -60.7788,
  -60.8332,
  -60.8761,
  -60.9065,
  -60.9236,
  -60.9266,
  -60.9143,
  -60.8884,
  -60.8481,
  -60.7933,
  -60.7247,
  -60.6432,
  -60.5504,
  -60.4485,
  -60.3394,
  -60.2258,
  -60.1099,
  -59.9938,
  -59.8797,
  -59.7687,
  -59.6618,
  -59.5593,
  -59.4613,
  -59.3679,
  -59.2792,
  -59.1946,
  -59.1142,
  -59.0379,
  -58.9668,
  -58.901,
  -58.8397,
  -58.7849,
  -58.7356,
  -58.6922,
  -58.6547,
  -58.6228,
  -58.5974,
  -58.5788,
  -58.5677,
  -58.5639,
  -58.5669,
  -58.5758,
  -58.5888,
  -58.6032,
  -58.6158,
  -58.6236,
  -58.6238,
  -58.6148,
  -58.5952,
  -58.5662,
  -58.5283,
  -58.4832,
  -58.4326,
  -58.3783,
  -58.3213,
  -58.2611,
  -58.1995,
  -58.135,
  -58.067,
  -57.9951,
  -57.9184,
  -57.8371,
  -57.7504,
  -57.6589,
  -57.5624,
  -57.4614,
  -57.3559,
  -57.2453,
  -57.1296,
  -57.0083,
  -56.8812,
  -56.7482,
  -56.6094,
  -56.4656,
  -56.3182,
  -56.1684,
  -56.0178,
  -55.868,
  -55.7214,
  -55.5791,
  -55.4418,
  -55.3106,
  -55.1855,
  -55.0672,
  -54.9555,
  -54.8485,
  -54.747,
  -54.6492,
  -54.5544,
  -54.4612,
  -54.3687,
  -54.2762,
  -54.1832,
  -54.0899,
  -53.9964,
  -53.9024,
  -53.8093,
  -53.7177,
  -53.629,
  -53.544,
  -53.4628,
  -53.3858,
  -53.3129,
  -53.2443,
  -53.1793,
  -53.1164,
  -53.0546,
  -52.994,
  -52.9347,
  -52.877,
  -52.8218,
  -52.7699,
  -52.7221,
  -52.6793,
  -52.6415,
  -52.6077,
  -52.5771,
  -52.5494,
  -52.5241,
  -52.5006,
  -52.4783,
  -52.4592,
  -52.4436,
  -52.4332,
  -52.4292,
  -52.4327,
  -52.445,
  -52.4662,
  -52.4957,
  -52.532,
  -52.5731,
  -52.6166,
  -52.6597,
  -52.7005,
  -52.7369,
  -52.7679,
  -52.7934,
  -52.814,
  -52.8309,
  -52.8453,
  -52.8581,
  -52.8702,
  -52.882,
  -52.893,
  -52.9032,
  -52.9119,
  -52.9196,
  -52.9259,
  -52.93,
  -52.932,
  -52.9316,
  -52.9293,
  -52.9253,
  -52.9205,
  -52.9157,
  -52.9115,
  -52.9089,
  -52.9087,
  -52.9128,
  -52.9225,
  -52.9397,
  -52.9661,
  -41.8276,
  -42.0028,
  -42.175,
  -42.348,
  -42.5324,
  -42.7232,
  -42.9231,
  -43.1293,
  -43.3406,
  -43.5545,
  -43.7715,
  -43.9902,
  -44.21,
  -44.4328,
  -44.6601,
  -44.8919,
  -45.1313,
  -45.3782,
  -45.6311,
  -45.8909,
  -46.1544,
  -46.4204,
  -46.6871,
  -46.9549,
  -47.2223,
  -47.489,
  -47.7541,
  -48.0176,
  -48.2794,
  -48.5381,
  -48.7914,
  -49.0404,
  -49.2816,
  -49.5143,
  -49.7376,
  -49.9504,
  -50.1517,
  -50.3417,
  -50.5193,
  -50.6859,
  -50.8423,
  -50.9892,
  -51.1275,
  -51.2575,
  -51.3795,
  -51.4934,
  -51.6023,
  -51.7068,
  -51.808,
  -51.9076,
  -52.0071,
  -52.1081,
  -52.2118,
  -52.3175,
  -52.4257,
  -52.5351,
  -52.6443,
  -52.7532,
  -52.8609,
  -52.9672,
  -53.0721,
  -53.1756,
  -53.2768,
  -53.3776,
  -53.4768,
  -53.574,
  -53.6689,
  -53.7619,
  -53.8536,
  -53.9456,
  -54.0387,
  -54.1348,
  -54.2344,
  -54.3382,
  -54.446,
  -54.5585,
  -54.6756,
  -54.7962,
  -54.9209,
  -55.0484,
  -55.1815,
  -55.32,
  -55.4651,
  -55.6179,
  -55.7805,
  -55.954,
  -56.1394,
  -56.3363,
  -56.5434,
  -56.7582,
  -56.9791,
  -57.2025,
  -57.4244,
  -57.6402,
  -57.8452,
  -58.0346,
  -58.2045,
  -58.3507,
  -58.4736,
  -58.5726,
  -58.6492,
  -58.7066,
  -58.7479,
  -58.7773,
  -58.7985,
  -58.8148,
  -58.8286,
  -58.8398,
  -58.849,
  -58.8561,
  -58.8614,
  -58.8642,
  -58.8647,
  -58.8644,
  -58.8644,
  -58.8661,
  -58.8712,
  -58.88,
  -58.8959,
  -58.9181,
  -58.9466,
  -58.9804,
  -59.0192,
  -59.0625,
  -59.1106,
  -59.1634,
  -59.2222,
  -59.2876,
  -59.3604,
  -59.4411,
  -59.5289,
  -59.6228,
  -59.7206,
  -59.82,
  -59.9186,
  -60.0133,
  -60.1017,
  -60.1818,
  -60.2516,
  -60.3118,
  -60.3605,
  -60.3972,
  -60.4208,
  -60.4312,
  -60.4274,
  -60.4093,
  -60.3767,
  -60.33,
  -60.2692,
  -60.1949,
  -60.1079,
  -60.0097,
  -59.9023,
  -59.788,
  -59.669,
  -59.5477,
  -59.4263,
  -59.307,
  -59.1912,
  -59.0798,
  -58.9724,
  -58.8714,
  -58.7761,
  -58.6866,
  -58.6021,
  -58.5225,
  -58.4476,
  -58.3779,
  -58.3137,
  -58.2548,
  -58.2011,
  -58.1526,
  -58.1098,
  -58.0728,
  -58.0413,
  -58.0162,
  -57.9981,
  -57.9875,
  -57.9847,
  -57.9889,
  -57.9991,
  -58.0131,
  -58.0289,
  -58.0429,
  -58.052,
  -58.0522,
  -58.0439,
  -58.0248,
  -57.9956,
  -57.9571,
  -57.9115,
  -57.8604,
  -57.8056,
  -57.7483,
  -57.689,
  -57.6276,
  -57.5638,
  -57.4969,
  -57.4267,
  -57.3527,
  -57.2747,
  -57.1921,
  -57.1053,
  -57.0142,
  -56.9185,
  -56.8184,
  -56.7138,
  -56.6041,
  -56.489,
  -56.3681,
  -56.2412,
  -56.1088,
  -55.9717,
  -55.8301,
  -55.6867,
  -55.5422,
  -55.3984,
  -55.2571,
  -55.1191,
  -54.9857,
  -54.8573,
  -54.7344,
  -54.6177,
  -54.5069,
  -54.4012,
  -54.2999,
  -54.2023,
  -54.1079,
  -54.0154,
  -53.9233,
  -53.8313,
  -53.7388,
  -53.6458,
  -53.5527,
  -53.4593,
  -53.3666,
  -53.2757,
  -53.1878,
  -53.1036,
  -53.0238,
  -52.9486,
  -52.8778,
  -52.8113,
  -52.7491,
  -52.6896,
  -52.6312,
  -52.5732,
  -52.5178,
  -52.4644,
  -52.4133,
  -52.3654,
  -52.3208,
  -52.2805,
  -52.2443,
  -52.2117,
  -52.1817,
  -52.1537,
  -52.1272,
  -52.1026,
  -52.0796,
  -52.0592,
  -52.0425,
  -52.0311,
  -52.0265,
  -52.0302,
  -52.043,
  -52.0651,
  -52.0958,
  -52.1338,
  -52.1764,
  -52.2212,
  -52.2655,
  -52.3069,
  -52.344,
  -52.3755,
  -52.4012,
  -52.4223,
  -52.4403,
  -52.4566,
  -52.4723,
  -52.4882,
  -52.5047,
  -52.5212,
  -52.5369,
  -52.5516,
  -52.5647,
  -52.5755,
  -52.5828,
  -52.5885,
  -52.5918,
  -52.5932,
  -52.5934,
  -52.5934,
  -52.5934,
  -52.5941,
  -52.5963,
  -52.6004,
  -52.6078,
  -52.6197,
  -52.6377,
  -52.6632,
  -41.5279,
  -41.703,
  -41.8724,
  -42.0408,
  -42.2176,
  -42.398,
  -42.6018,
  -42.8051,
  -43.0096,
  -43.2151,
  -43.4236,
  -43.6327,
  -43.8435,
  -44.0576,
  -44.2759,
  -44.4992,
  -44.7278,
  -44.9631,
  -45.2051,
  -45.4552,
  -45.7087,
  -45.9683,
  -46.2286,
  -46.4903,
  -46.7505,
  -47.0106,
  -47.2689,
  -47.5251,
  -47.7791,
  -48.0297,
  -48.2757,
  -48.5156,
  -48.7485,
  -48.9741,
  -49.1905,
  -49.3977,
  -49.5944,
  -49.7805,
  -49.9559,
  -50.1202,
  -50.2746,
  -50.421,
  -50.5594,
  -50.69,
  -50.8132,
  -50.9297,
  -51.0411,
  -51.1487,
  -51.2537,
  -51.3577,
  -51.4618,
  -51.5673,
  -51.675,
  -51.7844,
  -51.8957,
  -52.008,
  -52.1191,
  -52.2311,
  -52.3424,
  -52.4534,
  -52.5635,
  -52.6731,
  -52.782,
  -52.8898,
  -52.9962,
  -53.101,
  -53.2041,
  -53.3058,
  -53.4067,
  -53.5085,
  -53.6122,
  -53.7192,
  -53.8302,
  -53.9448,
  -54.0651,
  -54.1905,
  -54.3205,
  -54.4542,
  -54.5914,
  -54.7326,
  -54.8774,
  -55.0268,
  -55.1817,
  -55.3427,
  -55.5114,
  -55.6889,
  -55.8758,
  -56.0721,
  -56.2768,
  -56.4882,
  -56.7047,
  -56.9209,
  -57.1359,
  -57.3433,
  -57.5387,
  -57.7173,
  -57.8751,
  -58.0093,
  -58.1188,
  -58.2043,
  -58.2681,
  -58.3136,
  -58.3444,
  -58.3645,
  -58.3781,
  -58.3885,
  -58.398,
  -58.4067,
  -58.4146,
  -58.4217,
  -58.4264,
  -58.4302,
  -58.4319,
  -58.4322,
  -58.4324,
  -58.4337,
  -58.4376,
  -58.4456,
  -58.4588,
  -58.4777,
  -58.502,
  -58.5317,
  -58.566,
  -58.6051,
  -58.6497,
  -58.6998,
  -58.7565,
  -58.8211,
  -58.8938,
  -58.9752,
  -59.063,
  -59.158,
  -59.2568,
  -59.3567,
  -59.4551,
  -59.5487,
  -59.6348,
  -59.7116,
  -59.7777,
  -59.8324,
  -59.875,
  -59.905,
  -59.9218,
  -59.9253,
  -59.9146,
  -59.8899,
  -59.8514,
  -59.7989,
  -59.733,
  -59.6541,
  -59.5628,
  -59.4607,
  -59.3485,
  -59.2303,
  -59.1073,
  -58.9818,
  -58.8561,
  -58.7327,
  -58.613,
  -58.4981,
  -58.3887,
  -58.2851,
  -58.1884,
  -58.0984,
  -58.0144,
  -57.936,
  -57.8629,
  -57.7951,
  -57.7327,
  -57.6757,
  -57.6237,
  -57.5766,
  -57.535,
  -57.4988,
  -57.4681,
  -57.4436,
  -57.425,
  -57.4148,
  -57.4123,
  -57.4167,
  -57.4266,
  -57.4404,
  -57.4559,
  -57.4697,
  -57.4787,
  -57.4802,
  -57.4713,
  -57.4517,
  -57.4219,
  -57.383,
  -57.3366,
  -57.2849,
  -57.2297,
  -57.1719,
  -57.1127,
  -57.0518,
  -56.9892,
  -56.924,
  -56.8565,
  -56.786,
  -56.7123,
  -56.6349,
  -56.5534,
  -56.4671,
  -56.3774,
  -56.2834,
  -56.1846,
  -56.081,
  -55.972,
  -55.8571,
  -55.7364,
  -55.6102,
  -55.4793,
  -55.345,
  -55.208,
  -55.0696,
  -54.9316,
  -54.7957,
  -54.6628,
  -54.5336,
  -54.4089,
  -54.2892,
  -54.1746,
  -54.0654,
  -53.9605,
  -53.8597,
  -53.7622,
  -53.6681,
  -53.5759,
  -53.4844,
  -53.3926,
  -53.3002,
  -53.2073,
  -53.1133,
  -53.0203,
  -52.9279,
  -52.8372,
  -52.7497,
  -52.6658,
  -52.5863,
  -52.5114,
  -52.4412,
  -52.3759,
  -52.3153,
  -52.2579,
  -52.2026,
  -52.149,
  -52.0974,
  -52.0483,
  -52.0015,
  -51.9574,
  -51.9165,
  -51.8784,
  -51.8437,
  -51.8117,
  -51.782,
  -51.7533,
  -51.7258,
  -51.6996,
  -51.6755,
  -51.6541,
  -51.6371,
  -51.6256,
  -51.6213,
  -51.6255,
  -51.6391,
  -51.6623,
  -51.6941,
  -51.7331,
  -51.7771,
  -51.8228,
  -51.8672,
  -51.9092,
  -51.9465,
  -51.9783,
  -52.0043,
  -52.0257,
  -52.0448,
  -52.0627,
  -52.0815,
  -52.1013,
  -52.1225,
  -52.1446,
  -52.1664,
  -52.1873,
  -52.206,
  -52.2218,
  -52.2343,
  -52.2438,
  -52.2506,
  -52.2558,
  -52.2604,
  -52.265,
  -52.2699,
  -52.2754,
  -52.2823,
  -52.2906,
  -52.3014,
  -52.3158,
  -52.3349,
  -52.3601,
  -41.2292,
  -41.4027,
  -41.5709,
  -41.7397,
  -41.9136,
  -42.096,
  -42.2855,
  -42.4807,
  -42.678,
  -42.8772,
  -43.0777,
  -43.2791,
  -43.4824,
  -43.6899,
  -43.9002,
  -44.1149,
  -44.3346,
  -44.5593,
  -44.7915,
  -45.0289,
  -45.2744,
  -45.5237,
  -45.7769,
  -46.0306,
  -46.2844,
  -46.5367,
  -46.7872,
  -47.0357,
  -47.2813,
  -47.5234,
  -47.7608,
  -47.9926,
  -48.2174,
  -48.4352,
  -48.6442,
  -48.8461,
  -49.0379,
  -49.2199,
  -49.3917,
  -49.5538,
  -49.7075,
  -49.8533,
  -49.9915,
  -50.1222,
  -50.2459,
  -50.3635,
  -50.4765,
  -50.5864,
  -50.6948,
  -50.8028,
  -50.91,
  -51.0198,
  -51.1312,
  -51.2442,
  -51.3587,
  -51.4737,
  -51.5886,
  -51.7033,
  -51.8184,
  -51.9332,
  -52.0482,
  -52.1635,
  -52.2784,
  -52.3927,
  -52.5058,
  -52.6179,
  -52.7285,
  -52.8371,
  -52.9468,
  -53.0579,
  -53.1716,
  -53.289,
  -53.4107,
  -53.5375,
  -53.6694,
  -53.8068,
  -53.9486,
  -54.094,
  -54.2429,
  -54.3957,
  -54.552,
  -54.713,
  -54.8779,
  -55.0481,
  -55.2237,
  -55.407,
  -55.5979,
  -55.7964,
  -56.0018,
  -56.2128,
  -56.4268,
  -56.6405,
  -56.8496,
  -57.0499,
  -57.2362,
  -57.4039,
  -57.5498,
  -57.6711,
  -57.7672,
  -57.8394,
  -57.8902,
  -57.9236,
  -57.9431,
  -57.9523,
  -57.9577,
  -57.9613,
  -57.9652,
  -57.97,
  -57.9753,
  -57.9809,
  -57.9857,
  -57.9893,
  -57.9912,
  -57.9917,
  -57.9919,
  -57.9926,
  -57.9957,
  -58.0023,
  -58.0133,
  -58.0293,
  -58.0503,
  -58.0759,
  -58.1064,
  -58.1406,
  -58.1818,
  -58.2295,
  -58.2849,
  -58.3486,
  -58.4213,
  -58.5031,
  -58.5922,
  -58.6877,
  -58.7864,
  -58.8857,
  -58.9825,
  -59.0737,
  -59.1565,
  -59.2291,
  -59.2902,
  -59.3391,
  -59.3755,
  -59.3988,
  -59.4089,
  -59.4057,
  -59.3876,
  -59.3571,
  -59.3131,
  -59.2559,
  -59.1859,
  -59.1034,
  -59.0094,
  -58.9047,
  -58.7911,
  -58.6707,
  -58.5454,
  -58.4171,
  -58.2884,
  -58.1618,
  -58.0393,
  -57.9219,
  -57.8103,
  -57.7052,
  -57.6075,
  -57.5173,
  -57.4339,
  -57.3568,
  -57.2854,
  -57.2187,
  -57.1587,
  -57.1036,
  -57.0535,
  -57.0083,
  -56.9682,
  -56.9333,
  -56.9037,
  -56.8803,
  -56.863,
  -56.8529,
  -56.8501,
  -56.8535,
  -56.8619,
  -56.8736,
  -56.8868,
  -56.8989,
  -56.9064,
  -56.9064,
  -56.8965,
  -56.876,
  -56.8453,
  -56.8056,
  -56.7587,
  -56.7067,
  -56.6511,
  -56.5926,
  -56.5336,
  -56.4739,
  -56.4124,
  -56.3495,
  -56.2856,
  -56.2193,
  -56.1505,
  -56.0787,
  -56.0034,
  -55.9244,
  -55.8409,
  -55.7531,
  -55.6603,
  -55.5626,
  -55.4596,
  -55.3504,
  -55.2353,
  -55.1147,
  -54.9898,
  -54.8614,
  -54.7305,
  -54.5984,
  -54.4662,
  -54.3359,
  -54.2086,
  -54.0844,
  -53.9639,
  -53.8479,
  -53.7355,
  -53.6282,
  -53.5247,
  -53.4248,
  -53.3279,
  -53.2339,
  -53.1418,
  -53.0506,
  -52.9589,
  -52.8666,
  -52.774,
  -52.6812,
  -52.5885,
  -52.4966,
  -52.4063,
  -52.3188,
  -52.2349,
  -52.1548,
  -52.0795,
  -52.0089,
  -51.9436,
  -51.8831,
  -51.8271,
  -51.7739,
  -51.7235,
  -51.675,
  -51.6295,
  -51.5865,
  -51.546,
  -51.508,
  -51.472,
  -51.438,
  -51.4059,
  -51.3754,
  -51.3458,
  -51.3161,
  -51.2884,
  -51.2632,
  -51.2415,
  -51.2247,
  -51.2141,
  -51.2109,
  -51.2164,
  -51.2314,
  -51.256,
  -51.2891,
  -51.3291,
  -51.3739,
  -51.4207,
  -51.4664,
  -51.5088,
  -51.5464,
  -51.5781,
  -51.6045,
  -51.6261,
  -51.6459,
  -51.666,
  -51.6876,
  -51.7112,
  -51.737,
  -51.7646,
  -51.7927,
  -51.8197,
  -51.8443,
  -51.8656,
  -51.8828,
  -51.8963,
  -51.9071,
  -51.9162,
  -51.925,
  -51.9342,
  -51.944,
  -51.9543,
  -51.9656,
  -51.9782,
  -51.9927,
  -52.0099,
  -52.0307,
  -52.0564,
  -40.936,
  -41.1096,
  -41.2782,
  -41.4445,
  -41.6169,
  -41.7889,
  -41.9735,
  -42.1622,
  -42.3486,
  -42.5416,
  -42.7375,
  -42.9336,
  -43.1328,
  -43.3332,
  -43.5351,
  -43.7435,
  -43.9551,
  -44.1714,
  -44.3927,
  -44.6213,
  -44.856,
  -45.0965,
  -45.3397,
  -45.5839,
  -45.8285,
  -46.0713,
  -46.313,
  -46.5524,
  -46.789,
  -47.0216,
  -47.2504,
  -47.4735,
  -47.6905,
  -47.9012,
  -48.1048,
  -48.3008,
  -48.4877,
  -48.6655,
  -48.8338,
  -48.9935,
  -49.1453,
  -49.2902,
  -49.428,
  -49.5587,
  -49.6828,
  -49.8002,
  -49.9142,
  -50.0258,
  -50.1369,
  -50.2481,
  -50.3601,
  -50.4735,
  -50.5882,
  -50.7045,
  -50.8217,
  -50.9392,
  -51.0563,
  -51.1738,
  -51.2917,
  -51.4104,
  -51.5299,
  -51.6491,
  -51.7698,
  -51.8901,
  -52.0097,
  -52.1284,
  -52.2457,
  -52.3628,
  -52.4806,
  -52.6004,
  -52.7234,
  -52.8504,
  -52.9825,
  -53.1197,
  -53.2617,
  -53.4093,
  -53.5613,
  -53.7173,
  -53.8759,
  -54.0391,
  -54.2061,
  -54.3769,
  -54.5525,
  -54.7323,
  -54.9173,
  -55.1083,
  -55.3051,
  -55.5084,
  -55.7172,
  -55.9301,
  -56.1443,
  -56.356,
  -56.5613,
  -56.7551,
  -56.9332,
  -57.0908,
  -57.2241,
  -57.3327,
  -57.4156,
  -57.4747,
  -57.5131,
  -57.5345,
  -57.5429,
  -57.5433,
  -57.5399,
  -57.536,
  -57.5335,
  -57.5334,
  -57.5351,
  -57.5378,
  -57.5405,
  -57.5428,
  -57.5438,
  -57.5436,
  -57.543,
  -57.5432,
  -57.5442,
  -57.5493,
  -57.5584,
  -57.5717,
  -57.5895,
  -57.6118,
  -57.6388,
  -57.671,
  -57.7094,
  -57.7548,
  -57.8087,
  -57.8718,
  -57.9445,
  -58.026,
  -58.115,
  -58.2099,
  -58.3074,
  -58.4048,
  -58.4991,
  -58.5873,
  -58.6647,
  -58.7325,
  -58.7881,
  -58.8313,
  -58.8616,
  -58.8786,
  -58.8825,
  -58.8731,
  -58.8504,
  -58.8148,
  -58.7662,
  -58.7053,
  -58.6323,
  -58.5477,
  -58.4521,
  -58.3466,
  -58.2323,
  -58.1114,
  -57.9852,
  -57.8556,
  -57.725,
  -57.5966,
  -57.4723,
  -57.3521,
  -57.239,
  -57.1329,
  -57.0347,
  -56.9447,
  -56.862,
  -56.7863,
  -56.7165,
  -56.6528,
  -56.5949,
  -56.542,
  -56.494,
  -56.4507,
  -56.4124,
  -56.3792,
  -56.351,
  -56.3282,
  -56.3114,
  -56.3012,
  -56.2973,
  -56.2985,
  -56.3041,
  -56.3125,
  -56.3218,
  -56.3303,
  -56.3338,
  -56.3311,
  -56.3191,
  -56.2972,
  -56.2657,
  -56.2255,
  -56.1784,
  -56.1263,
  -56.0712,
  -56.0142,
  -55.956,
  -55.8976,
  -55.8384,
  -55.7787,
  -55.7184,
  -55.6565,
  -55.5929,
  -55.5268,
  -55.4576,
  -55.3851,
  -55.308,
  -55.2261,
  -55.1392,
  -55.0473,
  -54.9497,
  -54.8461,
  -54.7364,
  -54.6203,
  -54.5009,
  -54.3783,
  -54.2534,
  -54.1274,
  -54.0015,
  -53.877,
  -53.7553,
  -53.6368,
  -53.5215,
  -53.4098,
  -53.3021,
  -53.1977,
  -53.0963,
  -52.9978,
  -52.9016,
  -52.808,
  -52.7159,
  -52.6244,
  -52.5328,
  -52.4406,
  -52.3481,
  -52.2558,
  -52.1638,
  -52.0726,
  -51.9827,
  -51.8953,
  -51.8113,
  -51.7305,
  -51.6543,
  -51.583,
  -51.5167,
  -51.4556,
  -51.3985,
  -51.3465,
  -51.2978,
  -51.2525,
  -51.2093,
  -51.1693,
  -51.1309,
  -51.0945,
  -51.0594,
  -51.0254,
  -50.9922,
  -50.9598,
  -50.9283,
  -50.8979,
  -50.869,
  -50.843,
  -50.8216,
  -50.8056,
  -50.7966,
  -50.7956,
  -50.8033,
  -50.8204,
  -50.8467,
  -50.8813,
  -50.923,
  -50.9688,
  -51.0161,
  -51.0622,
  -51.1047,
  -51.142,
  -51.1736,
  -51.2001,
  -51.2229,
  -51.2439,
  -51.2653,
  -51.2892,
  -51.3165,
  -51.3471,
  -51.3802,
  -51.4144,
  -51.4478,
  -51.4776,
  -51.5046,
  -51.527,
  -51.5452,
  -51.5602,
  -51.5735,
  -51.5864,
  -51.5998,
  -51.6141,
  -51.6294,
  -51.6455,
  -51.6625,
  -51.6811,
  -51.7016,
  -51.725,
  -51.7523,
  -40.6581,
  -40.8296,
  -40.9946,
  -41.1664,
  -41.329,
  -41.4951,
  -41.6776,
  -41.8519,
  -42.0217,
  -42.2132,
  -42.406,
  -42.5998,
  -42.7924,
  -42.9874,
  -43.1801,
  -43.3857,
  -43.593,
  -43.8022,
  -44.0152,
  -44.2334,
  -44.4578,
  -44.6871,
  -44.919,
  -45.1521,
  -45.3846,
  -45.617,
  -45.8485,
  -46.0781,
  -46.3061,
  -46.5308,
  -46.7508,
  -46.9656,
  -47.1748,
  -47.378,
  -47.5752,
  -47.7657,
  -47.9479,
  -48.1211,
  -48.2861,
  -48.4422,
  -48.593,
  -48.7365,
  -48.8735,
  -49.0042,
  -49.1287,
  -49.2479,
  -49.3629,
  -49.4762,
  -49.5892,
  -49.7032,
  -49.8179,
  -49.934,
  -50.0516,
  -50.1702,
  -50.2894,
  -50.4074,
  -50.5268,
  -50.6466,
  -50.7672,
  -50.8891,
  -51.0125,
  -51.1372,
  -51.2627,
  -51.3885,
  -51.5142,
  -51.6391,
  -51.763,
  -51.8869,
  -52.0121,
  -52.1401,
  -52.2716,
  -52.4077,
  -52.5478,
  -52.694,
  -52.845,
  -53.0011,
  -53.1617,
  -53.3263,
  -53.4947,
  -53.667,
  -53.8433,
  -54.0237,
  -54.2091,
  -54.3989,
  -54.593,
  -54.7925,
  -54.9969,
  -55.2069,
  -55.4214,
  -55.6379,
  -55.8528,
  -56.0641,
  -56.2665,
  -56.4551,
  -56.6255,
  -56.7736,
  -56.8968,
  -56.9934,
  -57.0638,
  -57.1103,
  -57.1364,
  -57.1462,
  -57.1441,
  -57.1347,
  -57.1228,
  -57.1112,
  -57.1021,
  -57.0963,
  -57.0935,
  -57.0917,
  -57.0915,
  -57.0913,
  -57.09,
  -57.0884,
  -57.0866,
  -57.0855,
  -57.0862,
  -57.0895,
  -57.0966,
  -57.1074,
  -57.1223,
  -57.1417,
  -57.1656,
  -57.1952,
  -57.2312,
  -57.2747,
  -57.3273,
  -57.3894,
  -57.4613,
  -57.5412,
  -57.6294,
  -57.7227,
  -57.8181,
  -57.9127,
  -58.0036,
  -58.0873,
  -58.1614,
  -58.2238,
  -58.2742,
  -58.3118,
  -58.3365,
  -58.348,
  -58.3463,
  -58.3316,
  -58.3043,
  -58.2641,
  -58.2119,
  -58.1482,
  -58.0732,
  -57.9876,
  -57.8918,
  -57.7857,
  -57.6728,
  -57.5526,
  -57.4268,
  -57.2974,
  -57.1665,
  -57.0375,
  -56.9122,
  -56.7922,
  -56.6787,
  -56.5721,
  -56.4742,
  -56.3843,
  -56.3025,
  -56.2278,
  -56.1595,
  -56.0979,
  -56.0417,
  -55.9908,
  -55.9449,
  -55.9035,
  -55.8672,
  -55.8352,
  -55.8083,
  -55.7851,
  -55.7682,
  -55.7575,
  -55.7517,
  -55.7503,
  -55.7522,
  -55.7559,
  -55.7604,
  -55.7639,
  -55.7636,
  -55.7571,
  -55.7429,
  -55.7195,
  -55.687,
  -55.6466,
  -55.5997,
  -55.5481,
  -55.4939,
  -55.438,
  -55.3815,
  -55.325,
  -55.2684,
  -55.2122,
  -55.1556,
  -55.0983,
  -55.0395,
  -54.9777,
  -54.9146,
  -54.8479,
  -54.7769,
  -54.701,
  -54.6199,
  -54.5334,
  -54.4409,
  -54.3425,
  -54.2381,
  -54.1284,
  -54.0146,
  -53.8977,
  -53.779,
  -53.6593,
  -53.54,
  -53.4221,
  -53.3066,
  -53.1942,
  -53.0846,
  -52.9777,
  -52.8743,
  -52.7734,
  -52.6747,
  -52.5781,
  -52.483,
  -52.3898,
  -52.2976,
  -52.2057,
  -52.1138,
  -52.0216,
  -51.9286,
  -51.8368,
  -51.7455,
  -51.6551,
  -51.5661,
  -51.4793,
  -51.3949,
  -51.314,
  -51.2367,
  -51.1642,
  -51.0968,
  -51.0344,
  -50.9773,
  -50.9251,
  -50.8774,
  -50.8336,
  -50.792,
  -50.7532,
  -50.7157,
  -50.6793,
  -50.6434,
  -50.6076,
  -50.5719,
  -50.5365,
  -50.5021,
  -50.4694,
  -50.4391,
  -50.413,
  -50.3921,
  -50.3776,
  -50.3712,
  -50.373,
  -50.3838,
  -50.4037,
  -50.4328,
  -50.4698,
  -50.5129,
  -50.559,
  -50.6069,
  -50.6532,
  -50.6957,
  -50.7331,
  -50.7646,
  -50.7913,
  -50.8146,
  -50.8367,
  -50.8597,
  -50.8861,
  -50.9169,
  -50.9522,
  -50.9907,
  -51.0308,
  -51.0706,
  -51.1078,
  -51.1409,
  -51.169,
  -51.1923,
  -51.2121,
  -51.2299,
  -51.247,
  -51.2647,
  -51.2834,
  -51.3033,
  -51.3242,
  -51.3462,
  -51.3694,
  -51.394,
  -51.4212,
  -51.4518,
  -40.3926,
  -40.5596,
  -40.7307,
  -40.8948,
  -41.0507,
  -41.2171,
  -41.3853,
  -41.5449,
  -41.699,
  -41.8866,
  -42.0884,
  -42.2784,
  -42.4626,
  -42.6543,
  -42.8456,
  -43.0411,
  -43.2473,
  -43.4511,
  -43.6564,
  -43.8649,
  -44.0792,
  -44.2965,
  -44.5164,
  -44.7373,
  -44.9586,
  -45.1798,
  -45.4005,
  -45.6204,
  -45.8391,
  -46.0549,
  -46.2664,
  -46.4729,
  -46.6743,
  -46.8702,
  -47.06,
  -47.2445,
  -47.4217,
  -47.5911,
  -47.7529,
  -47.9074,
  -48.0562,
  -48.1988,
  -48.3352,
  -48.466,
  -48.5912,
  -48.7112,
  -48.8277,
  -48.9425,
  -49.0575,
  -49.1722,
  -49.2889,
  -49.4072,
  -49.5264,
  -49.6465,
  -49.7666,
  -49.8867,
  -50.007,
  -50.1286,
  -50.2514,
  -50.376,
  -50.5026,
  -50.631,
  -50.761,
  -50.8919,
  -51.0228,
  -51.1537,
  -51.2828,
  -51.4128,
  -51.5451,
  -51.6802,
  -51.8198,
  -51.9638,
  -52.1127,
  -52.2665,
  -52.4247,
  -52.5877,
  -52.7552,
  -52.9271,
  -53.1029,
  -53.2828,
  -53.4672,
  -53.6564,
  -53.8505,
  -54.0496,
  -54.2523,
  -54.4609,
  -54.675,
  -54.8931,
  -55.114,
  -55.3356,
  -55.5542,
  -55.7658,
  -55.966,
  -56.1499,
  -56.3131,
  -56.452,
  -56.5644,
  -56.6496,
  -56.708,
  -56.7426,
  -56.7567,
  -56.7553,
  -56.7421,
  -56.7238,
  -56.7039,
  -56.6849,
  -56.6693,
  -56.6578,
  -56.6501,
  -56.6448,
  -56.6408,
  -56.6374,
  -56.6335,
  -56.6295,
  -56.6257,
  -56.6226,
  -56.6213,
  -56.6228,
  -56.6276,
  -56.6361,
  -56.6483,
  -56.665,
  -56.6855,
  -56.7125,
  -56.7466,
  -56.7886,
  -56.8399,
  -56.9009,
  -56.9717,
  -57.0511,
  -57.1374,
  -57.2283,
  -57.3207,
  -57.4118,
  -57.4979,
  -57.5768,
  -57.6456,
  -57.7029,
  -57.7482,
  -57.7806,
  -57.8005,
  -57.8073,
  -57.801,
  -57.781,
  -57.7497,
  -57.706,
  -57.6512,
  -57.5854,
  -57.5093,
  -57.4236,
  -57.3288,
  -57.2255,
  -57.1144,
  -56.9965,
  -56.8725,
  -56.7447,
  -56.6151,
  -56.4867,
  -56.3618,
  -56.2417,
  -56.1285,
  -56.0226,
  -55.9252,
  -55.8361,
  -55.7549,
  -55.6813,
  -55.6135,
  -55.5531,
  -55.4986,
  -55.4492,
  -55.4051,
  -55.3655,
  -55.3305,
  -55.2998,
  -55.2734,
  -55.2516,
  -55.2345,
  -55.2225,
  -55.2146,
  -55.2097,
  -55.2074,
  -55.2061,
  -55.205,
  -55.2029,
  -55.1973,
  -55.187,
  -55.1695,
  -55.1444,
  -55.1113,
  -55.071,
  -55.025,
  -54.9735,
  -54.9207,
  -54.8666,
  -54.8121,
  -54.7579,
  -54.7044,
  -54.6512,
  -54.5983,
  -54.5448,
  -54.4905,
  -54.4346,
  -54.3766,
  -54.3154,
  -54.2498,
  -54.1794,
  -54.1036,
  -54.0222,
  -53.9348,
  -53.8412,
  -53.7421,
  -53.638,
  -53.53,
  -53.4191,
  -53.3067,
  -53.1939,
  -53.0818,
  -52.9709,
  -52.8622,
  -52.7561,
  -52.6519,
  -52.5507,
  -52.4518,
  -52.355,
  -52.2594,
  -52.1649,
  -52.0714,
  -51.9784,
  -51.8858,
  -51.7935,
  -51.7013,
  -51.6092,
  -51.5175,
  -51.4265,
  -51.3361,
  -51.2468,
  -51.1588,
  -51.0726,
  -50.9886,
  -50.9071,
  -50.8293,
  -50.7556,
  -50.6866,
  -50.6228,
  -50.5645,
  -50.5118,
  -50.4639,
  -50.42,
  -50.3787,
  -50.3391,
  -50.3006,
  -50.2622,
  -50.2231,
  -50.1837,
  -50.144,
  -50.1034,
  -50.0651,
  -50.0295,
  -49.9977,
  -49.9714,
  -49.9515,
  -49.9394,
  -49.936,
  -49.9417,
  -49.9565,
  -49.9805,
  -50.013,
  -50.053,
  -50.0984,
  -50.1468,
  -50.1954,
  -50.2419,
  -50.2844,
  -50.3214,
  -50.3529,
  -50.3798,
  -50.4039,
  -50.4272,
  -50.4521,
  -50.4808,
  -50.5153,
  -50.5548,
  -50.5986,
  -50.6445,
  -50.6904,
  -50.7341,
  -50.7736,
  -50.808,
  -50.837,
  -50.8617,
  -50.8843,
  -50.9058,
  -50.928,
  -50.9513,
  -50.9759,
  -51.0018,
  -51.0287,
  -51.057,
  -51.087,
  -51.1195,
  -51.1548,
  -40.1485,
  -40.3053,
  -40.4683,
  -40.6315,
  -40.7938,
  -40.9451,
  -41.0957,
  -41.2573,
  -41.4118,
  -41.5851,
  -41.7829,
  -41.9705,
  -42.1551,
  -42.342,
  -42.5308,
  -42.7196,
  -42.9164,
  -43.1164,
  -43.3153,
  -43.5172,
  -43.7207,
  -43.9271,
  -44.1342,
  -44.3429,
  -44.552,
  -44.762,
  -44.972,
  -45.1819,
  -45.3904,
  -45.5974,
  -45.8004,
  -45.9989,
  -46.1924,
  -46.3811,
  -46.5655,
  -46.7446,
  -46.9168,
  -47.0825,
  -47.2408,
  -47.3932,
  -47.5396,
  -47.6807,
  -47.8168,
  -47.9479,
  -48.0726,
  -48.194,
  -48.3121,
  -48.4288,
  -48.5454,
  -48.6627,
  -48.7807,
  -48.9001,
  -49.0201,
  -49.1406,
  -49.2605,
  -49.3807,
  -49.5015,
  -49.6238,
  -49.7482,
  -49.8748,
  -50.0029,
  -50.1345,
  -50.2678,
  -50.403,
  -50.5391,
  -50.6748,
  -50.8105,
  -50.9468,
  -51.0849,
  -51.2267,
  -51.3727,
  -51.5238,
  -51.679,
  -51.8391,
  -52.0031,
  -52.1716,
  -52.3445,
  -52.5211,
  -52.703,
  -52.8892,
  -53.0808,
  -53.2776,
  -53.4804,
  -53.6882,
  -53.9017,
  -54.1208,
  -54.3445,
  -54.5716,
  -54.8,
  -55.0269,
  -55.2484,
  -55.4604,
  -55.6585,
  -55.8374,
  -55.9936,
  -56.1226,
  -56.2246,
  -56.2983,
  -56.3449,
  -56.3675,
  -56.3703,
  -56.3585,
  -56.3369,
  -56.3101,
  -56.2827,
  -56.2571,
  -56.2352,
  -56.2186,
  -56.2059,
  -56.196,
  -56.1878,
  -56.1806,
  -56.1735,
  -56.1664,
  -56.1598,
  -56.1533,
  -56.1497,
  -56.1488,
  -56.1514,
  -56.1575,
  -56.1675,
  -56.1819,
  -56.2013,
  -56.2266,
  -56.2588,
  -56.2995,
  -56.3495,
  -56.4093,
  -56.4783,
  -56.5557,
  -56.6394,
  -56.7269,
  -56.8153,
  -56.9014,
  -56.9827,
  -57.0549,
  -57.1182,
  -57.1702,
  -57.2104,
  -57.2382,
  -57.254,
  -57.2571,
  -57.2474,
  -57.2247,
  -57.19,
  -57.1441,
  -57.087,
  -57.02,
  -56.9436,
  -56.8588,
  -56.7658,
  -56.6648,
  -56.5565,
  -56.4415,
  -56.3206,
  -56.1956,
  -56.0685,
  -55.9421,
  -55.8174,
  -55.699,
  -55.5873,
  -55.4827,
  -55.3864,
  -55.2984,
  -55.2184,
  -55.146,
  -55.0802,
  -55.0207,
  -54.9672,
  -54.919,
  -54.8762,
  -54.8376,
  -54.8033,
  -54.7734,
  -54.7474,
  -54.7257,
  -54.708,
  -54.6941,
  -54.6837,
  -54.6754,
  -54.6687,
  -54.6624,
  -54.6547,
  -54.6469,
  -54.6365,
  -54.6218,
  -54.6014,
  -54.5745,
  -54.5411,
  -54.5016,
  -54.4569,
  -54.4081,
  -54.357,
  -54.305,
  -54.2532,
  -54.2015,
  -54.1505,
  -54.1,
  -54.0501,
  -54,
  -53.9492,
  -53.897,
  -53.843,
  -53.7862,
  -53.7255,
  -53.6601,
  -53.589,
  -53.5122,
  -53.4298,
  -53.3413,
  -53.2467,
  -53.1483,
  -53.0464,
  -52.9422,
  -52.8369,
  -52.7315,
  -52.627,
  -52.5237,
  -52.4223,
  -52.3232,
  -52.2266,
  -52.1317,
  -52.0377,
  -51.945,
  -51.8527,
  -51.7608,
  -51.6684,
  -51.5756,
  -51.4828,
  -51.39,
  -51.2975,
  -51.2053,
  -51.1142,
  -51.0238,
  -50.9345,
  -50.8464,
  -50.7595,
  -50.6739,
  -50.5903,
  -50.509,
  -50.4307,
  -50.3558,
  -50.2845,
  -50.2192,
  -50.1595,
  -50.1055,
  -50.0563,
  -50.0112,
  -49.9687,
  -49.9269,
  -49.8852,
  -49.8428,
  -49.7988,
  -49.7536,
  -49.7081,
  -49.6632,
  -49.6204,
  -49.5811,
  -49.5478,
  -49.5214,
  -49.5031,
  -49.4939,
  -49.4945,
  -49.5049,
  -49.5246,
  -49.5535,
  -49.5903,
  -49.6336,
  -49.6821,
  -49.7317,
  -49.7816,
  -49.8282,
  -49.8703,
  -49.907,
  -49.9385,
  -49.9656,
  -49.9905,
  -50.0152,
  -50.042,
  -50.0734,
  -50.111,
  -50.1549,
  -50.2025,
  -50.2536,
  -50.3055,
  -50.3555,
  -50.4018,
  -50.4426,
  -50.4778,
  -50.5084,
  -50.536,
  -50.5624,
  -50.5892,
  -50.617,
  -50.6462,
  -50.6771,
  -50.7096,
  -50.7442,
  -50.781,
  -50.8208,
  -50.8646,
  -39.9103,
  -40.0672,
  -40.2302,
  -40.3947,
  -40.5683,
  -40.7236,
  -40.8701,
  -41.0062,
  -41.148,
  -41.3148,
  -41.4914,
  -41.6808,
  -41.8637,
  -42.0479,
  -42.2341,
  -42.4195,
  -42.6049,
  -42.7964,
  -42.9901,
  -43.1855,
  -43.38,
  -43.5749,
  -43.771,
  -43.9673,
  -44.1654,
  -44.3644,
  -44.5646,
  -44.7648,
  -44.9646,
  -45.1631,
  -45.358,
  -45.5484,
  -45.7345,
  -45.9164,
  -46.0947,
  -46.2678,
  -46.4352,
  -46.597,
  -46.7511,
  -46.901,
  -47.0458,
  -47.1855,
  -47.321,
  -47.4524,
  -47.5791,
  -47.7019,
  -47.8219,
  -47.9403,
  -48.0584,
  -48.1768,
  -48.2958,
  -48.4158,
  -48.5359,
  -48.6555,
  -48.7738,
  -48.8933,
  -49.0137,
  -49.136,
  -49.261,
  -49.3888,
  -49.5194,
  -49.6533,
  -49.7895,
  -49.928,
  -50.068,
  -50.2082,
  -50.3488,
  -50.4902,
  -50.6337,
  -50.7803,
  -50.9321,
  -51.0876,
  -51.248,
  -51.4126,
  -51.5812,
  -51.7545,
  -51.9317,
  -52.1133,
  -52.3,
  -52.4917,
  -52.689,
  -52.8927,
  -53.1032,
  -53.3204,
  -53.5441,
  -53.7737,
  -54.0079,
  -54.2446,
  -54.4808,
  -54.7118,
  -54.9362,
  -55.1483,
  -55.3435,
  -55.5173,
  -55.6662,
  -55.7869,
  -55.8782,
  -55.9403,
  -55.9751,
  -55.9859,
  -55.9775,
  -55.9555,
  -55.9249,
  -55.8904,
  -55.8561,
  -55.8246,
  -55.7976,
  -55.7758,
  -55.7573,
  -55.7429,
  -55.7306,
  -55.7196,
  -55.7087,
  -55.6982,
  -55.6883,
  -55.68,
  -55.6738,
  -55.6707,
  -55.6708,
  -55.6749,
  -55.6831,
  -55.6957,
  -55.7134,
  -55.7372,
  -55.7681,
  -55.8076,
  -55.8563,
  -55.9145,
  -55.9808,
  -56.0555,
  -56.1356,
  -56.2186,
  -56.3019,
  -56.3824,
  -56.4576,
  -56.525,
  -56.5824,
  -56.6289,
  -56.6642,
  -56.6882,
  -56.7006,
  -56.7007,
  -56.6882,
  -56.6631,
  -56.626,
  -56.5777,
  -56.5194,
  -56.4518,
  -56.3755,
  -56.2921,
  -56.2005,
  -56.1027,
  -55.9977,
  -55.8859,
  -55.7689,
  -55.6478,
  -55.5249,
  -55.4015,
  -55.2806,
  -55.1649,
  -55.0557,
  -54.9537,
  -54.8592,
  -54.7723,
  -54.6939,
  -54.6225,
  -54.5577,
  -54.4989,
  -54.4457,
  -54.3984,
  -54.356,
  -54.3181,
  -54.2842,
  -54.2531,
  -54.2274,
  -54.2051,
  -54.1864,
  -54.1706,
  -54.1571,
  -54.1456,
  -54.1348,
  -54.1239,
  -54.1123,
  -54.0992,
  -54.0843,
  -54.0661,
  -54.0436,
  -54.0155,
  -53.9819,
  -53.9432,
  -53.9002,
  -53.8537,
  -53.8051,
  -53.7552,
  -53.7059,
  -53.6567,
  -53.6084,
  -53.5596,
  -53.5116,
  -53.4636,
  -53.4144,
  -53.3652,
  -53.3141,
  -53.2604,
  -53.2036,
  -53.1422,
  -53.0756,
  -53.0033,
  -52.9255,
  -52.8427,
  -52.755,
  -52.6631,
  -52.5678,
  -52.4706,
  -52.3732,
  -52.2756,
  -52.1792,
  -52.0842,
  -51.9905,
  -51.8989,
  -51.8089,
  -51.7201,
  -51.6316,
  -51.5427,
  -51.4539,
  -51.3641,
  -51.273,
  -51.1807,
  -51.0872,
  -50.9938,
  -50.9003,
  -50.8082,
  -50.7174,
  -50.6279,
  -50.5397,
  -50.4527,
  -50.3668,
  -50.2822,
  -50.1988,
  -50.1177,
  -50.039,
  -49.9638,
  -49.8923,
  -49.8255,
  -49.7643,
  -49.7084,
  -49.6574,
  -49.6101,
  -49.5646,
  -49.5191,
  -49.4721,
  -49.4235,
  -49.3731,
  -49.3211,
  -49.2689,
  -49.2178,
  -49.1699,
  -49.127,
  -49.0916,
  -49.0652,
  -49.0492,
  -49.0434,
  -49.0488,
  -49.0642,
  -49.0897,
  -49.124,
  -49.1656,
  -49.2121,
  -49.263,
  -49.3148,
  -49.3651,
  -49.4121,
  -49.4536,
  -49.4899,
  -49.521,
  -49.5486,
  -49.5743,
  -49.6006,
  -49.63,
  -49.6643,
  -49.7049,
  -49.7526,
  -49.8056,
  -49.8618,
  -49.9193,
  -49.9754,
  -50.0279,
  -50.0752,
  -50.1169,
  -50.1536,
  -50.187,
  -50.2187,
  -50.2502,
  -50.2826,
  -50.317,
  -50.3535,
  -50.3924,
  -50.4342,
  -50.4791,
  -50.5277,
  -50.5816,
  -39.721,
  -39.8871,
  -40.0418,
  -40.1939,
  -40.3587,
  -40.5116,
  -40.6471,
  -40.7892,
  -40.9361,
  -41.0893,
  -41.2347,
  -41.3991,
  -41.583,
  -41.769,
  -41.9515,
  -42.1311,
  -42.3115,
  -42.4907,
  -42.6762,
  -42.8653,
  -43.0534,
  -43.2394,
  -43.4254,
  -43.6125,
  -43.8006,
  -43.99,
  -44.1809,
  -44.3719,
  -44.5626,
  -44.7524,
  -44.9393,
  -45.1222,
  -45.3012,
  -45.4758,
  -45.648,
  -45.8162,
  -45.9794,
  -46.137,
  -46.2893,
  -46.4367,
  -46.5793,
  -46.7179,
  -46.8529,
  -46.9844,
  -47.112,
  -47.2365,
  -47.3582,
  -47.4784,
  -47.5977,
  -47.7157,
  -47.8351,
  -47.9549,
  -48.0745,
  -48.193,
  -48.311,
  -48.4292,
  -48.5486,
  -48.6702,
  -48.795,
  -48.9232,
  -49.0547,
  -49.1895,
  -49.3281,
  -49.469,
  -49.6117,
  -49.7544,
  -49.8987,
  -50.044,
  -50.1919,
  -50.3433,
  -50.4987,
  -50.6585,
  -50.8229,
  -50.9914,
  -51.1634,
  -51.3398,
  -51.5203,
  -51.7055,
  -51.8958,
  -52.0915,
  -52.2939,
  -52.5036,
  -52.7217,
  -52.9468,
  -53.181,
  -53.422,
  -53.6673,
  -53.9134,
  -54.1568,
  -54.3941,
  -54.621,
  -54.8324,
  -55.0241,
  -55.1919,
  -55.3328,
  -55.4436,
  -55.5238,
  -55.5741,
  -55.5967,
  -55.5956,
  -55.5758,
  -55.5427,
  -55.5035,
  -55.4618,
  -55.4214,
  -55.3844,
  -55.3531,
  -55.3269,
  -55.3051,
  -55.2865,
  -55.2702,
  -55.2553,
  -55.2407,
  -55.2267,
  -55.2136,
  -55.2022,
  -55.1934,
  -55.1879,
  -55.1861,
  -55.1884,
  -55.1952,
  -55.2056,
  -55.2222,
  -55.245,
  -55.275,
  -55.3135,
  -55.3609,
  -55.4173,
  -55.4821,
  -55.5535,
  -55.6293,
  -55.7072,
  -55.7844,
  -55.8583,
  -55.9269,
  -55.988,
  -56.0396,
  -56.0808,
  -56.1111,
  -56.1313,
  -56.1407,
  -56.1384,
  -56.1226,
  -56.0959,
  -56.0572,
  -56.0077,
  -55.9482,
  -55.8806,
  -55.8055,
  -55.7237,
  -55.6356,
  -55.5408,
  -55.4396,
  -55.3319,
  -55.2193,
  -55.1033,
  -54.9846,
  -54.8659,
  -54.7494,
  -54.6377,
  -54.5319,
  -54.4328,
  -54.3411,
  -54.2568,
  -54.1798,
  -54.1085,
  -54.0442,
  -53.9861,
  -53.9333,
  -53.8862,
  -53.844,
  -53.8058,
  -53.7719,
  -53.7417,
  -53.7152,
  -53.6919,
  -53.6714,
  -53.6536,
  -53.6376,
  -53.623,
  -53.6086,
  -53.5936,
  -53.5778,
  -53.5609,
  -53.5423,
  -53.5213,
  -53.4969,
  -53.4687,
  -53.4356,
  -53.3984,
  -53.3567,
  -53.3128,
  -53.2668,
  -53.2196,
  -53.1722,
  -53.125,
  -53.078,
  -53.031,
  -52.984,
  -52.9372,
  -52.8901,
  -52.8423,
  -52.7933,
  -52.7421,
  -52.688,
  -52.6299,
  -52.567,
  -52.4993,
  -52.4267,
  -52.3496,
  -52.2682,
  -52.1831,
  -52.0954,
  -52.0059,
  -51.9164,
  -51.8271,
  -51.7389,
  -51.6522,
  -51.5665,
  -51.4813,
  -51.398,
  -51.315,
  -51.2317,
  -51.1471,
  -51.0612,
  -50.9733,
  -50.8833,
  -50.7915,
  -50.6982,
  -50.6045,
  -50.5116,
  -50.4198,
  -50.3294,
  -50.241,
  -50.1539,
  -50.0679,
  -49.9828,
  -49.8989,
  -49.8164,
  -49.7356,
  -49.6571,
  -49.581,
  -49.5087,
  -49.4407,
  -49.3776,
  -49.3196,
  -49.266,
  -49.215,
  -49.1652,
  -49.1147,
  -49.0618,
  -49.0056,
  -48.9473,
  -48.8867,
  -48.8271,
  -48.7697,
  -48.7169,
  -48.6708,
  -48.6338,
  -48.6078,
  -48.5942,
  -48.5922,
  -48.6023,
  -48.6232,
  -48.6543,
  -48.6941,
  -48.7408,
  -48.7923,
  -48.8459,
  -48.8995,
  -48.9503,
  -48.9968,
  -49.0381,
  -49.0739,
  -49.1051,
  -49.1327,
  -49.1595,
  -49.1871,
  -49.2188,
  -49.256,
  -49.2997,
  -49.3509,
  -49.4081,
  -49.4692,
  -49.5319,
  -49.5935,
  -49.6518,
  -49.7055,
  -49.7535,
  -49.7967,
  -49.8361,
  -49.8735,
  -49.9103,
  -49.9482,
  -49.9882,
  -50.0311,
  -50.0774,
  -50.1264,
  -50.1804,
  -50.2395,
  -50.305,
  -39.568,
  -39.7228,
  -39.8745,
  -40.0195,
  -40.1716,
  -40.3077,
  -40.4499,
  -40.5889,
  -40.7316,
  -40.8694,
  -41.0012,
  -41.1364,
  -41.3106,
  -41.4958,
  -41.6772,
  -41.849,
  -42.0258,
  -42.2018,
  -42.3769,
  -42.5607,
  -42.7417,
  -42.9218,
  -43.0988,
  -43.2774,
  -43.4569,
  -43.6381,
  -43.82,
  -44.0015,
  -44.1838,
  -44.3652,
  -44.5445,
  -44.7207,
  -44.8935,
  -45.0633,
  -45.2301,
  -45.3934,
  -45.5523,
  -45.7064,
  -45.8559,
  -46.0006,
  -46.1417,
  -46.2791,
  -46.4136,
  -46.5441,
  -46.6725,
  -46.798,
  -46.9213,
  -47.0426,
  -47.1626,
  -47.282,
  -47.4012,
  -47.5204,
  -47.6389,
  -47.7559,
  -47.8725,
  -47.9891,
  -48.1071,
  -48.2279,
  -48.3519,
  -48.4786,
  -48.6102,
  -48.7456,
  -48.8847,
  -49.027,
  -49.1716,
  -49.3174,
  -49.4641,
  -49.6126,
  -49.7633,
  -49.9174,
  -50.0757,
  -50.2384,
  -50.4053,
  -50.5759,
  -50.7502,
  -50.9288,
  -51.1106,
  -51.2982,
  -51.4913,
  -51.6905,
  -51.8972,
  -52.1128,
  -52.338,
  -52.5731,
  -52.8177,
  -53.0696,
  -53.3253,
  -53.5808,
  -53.8317,
  -54.0737,
  -54.3024,
  -54.5125,
  -54.7001,
  -54.8616,
  -54.9926,
  -55.0929,
  -55.1613,
  -55.199,
  -55.2091,
  -55.1955,
  -55.1644,
  -55.1221,
  -55.074,
  -55.0253,
  -54.9794,
  -54.9377,
  -54.9023,
  -54.8724,
  -54.8471,
  -54.8249,
  -54.805,
  -54.7865,
  -54.7684,
  -54.7511,
  -54.7339,
  -54.7198,
  -54.7085,
  -54.7008,
  -54.6974,
  -54.6986,
  -54.7042,
  -54.7149,
  -54.731,
  -54.7533,
  -54.7825,
  -54.8201,
  -54.8661,
  -54.9205,
  -54.9822,
  -55.0497,
  -55.1206,
  -55.1926,
  -55.2632,
  -55.3302,
  -55.3909,
  -55.4451,
  -55.4905,
  -55.5265,
  -55.5528,
  -55.5694,
  -55.576,
  -55.5715,
  -55.5552,
  -55.527,
  -55.4872,
  -55.4369,
  -55.3772,
  -55.3098,
  -55.2358,
  -55.1559,
  -55.0706,
  -54.9794,
  -54.8824,
  -54.7795,
  -54.6718,
  -54.5609,
  -54.4471,
  -54.334,
  -54.2228,
  -54.1155,
  -54.0139,
  -53.9188,
  -53.8305,
  -53.7488,
  -53.6734,
  -53.6043,
  -53.5409,
  -53.4833,
  -53.4306,
  -53.3832,
  -53.3406,
  -53.3022,
  -53.268,
  -53.2372,
  -53.2096,
  -53.1849,
  -53.1628,
  -53.143,
  -53.1245,
  -53.1069,
  -53.0893,
  -53.0701,
  -53.0512,
  -53.0313,
  -53.0099,
  -52.9873,
  -52.9621,
  -52.9342,
  -52.9026,
  -52.8675,
  -52.8293,
  -52.7883,
  -52.7453,
  -52.7008,
  -52.6555,
  -52.6099,
  -52.5638,
  -52.5175,
  -52.4709,
  -52.4241,
  -52.3773,
  -52.3302,
  -52.2824,
  -52.2326,
  -52.1802,
  -52.1248,
  -52.0657,
  -52.0027,
  -51.9344,
  -51.8631,
  -51.7881,
  -51.7102,
  -51.6304,
  -51.5492,
  -51.4676,
  -51.3866,
  -51.3065,
  -51.2276,
  -51.1496,
  -51.0723,
  -50.9953,
  -50.9178,
  -50.8393,
  -50.7585,
  -50.675,
  -50.5892,
  -50.5004,
  -50.4093,
  -50.3163,
  -50.2228,
  -50.1298,
  -50.0387,
  -49.9492,
  -49.8616,
  -49.7755,
  -49.6906,
  -49.6066,
  -49.5235,
  -49.4418,
  -49.3615,
  -49.282,
  -49.2059,
  -49.1328,
  -49.0633,
  -48.9982,
  -48.9375,
  -48.8806,
  -48.8252,
  -48.7702,
  -48.7129,
  -48.6529,
  -48.5889,
  -48.5225,
  -48.4552,
  -48.3891,
  -48.3261,
  -48.2694,
  -48.2213,
  -48.1839,
  -48.159,
  -48.1477,
  -48.1498,
  -48.1643,
  -48.19,
  -48.2262,
  -48.2707,
  -48.3215,
  -48.3763,
  -48.4324,
  -48.487,
  -48.5381,
  -48.5842,
  -48.6249,
  -48.66,
  -48.691,
  -48.7188,
  -48.7462,
  -48.7756,
  -48.8091,
  -48.8489,
  -48.8947,
  -48.9493,
  -49.0105,
  -49.0762,
  -49.1434,
  -49.2101,
  -49.2738,
  -49.3333,
  -49.3876,
  -49.4373,
  -49.483,
  -49.5264,
  -49.5692,
  -49.6133,
  -49.6598,
  -49.7102,
  -49.7648,
  -49.824,
  -49.8886,
  -49.9594,
  -50.0382,
  -39.4245,
  -39.5698,
  -39.716,
  -39.8575,
  -39.9977,
  -40.1215,
  -40.2648,
  -40.3959,
  -40.5331,
  -40.6603,
  -40.7833,
  -40.9093,
  -41.0672,
  -41.2356,
  -41.4158,
  -41.5723,
  -41.7479,
  -41.9253,
  -42.0983,
  -42.2723,
  -42.4475,
  -42.6219,
  -42.791,
  -42.9607,
  -43.1328,
  -43.3061,
  -43.4806,
  -43.6552,
  -43.8297,
  -44.0034,
  -44.176,
  -44.3457,
  -44.5129,
  -44.6777,
  -44.8399,
  -44.9987,
  -45.1538,
  -45.3037,
  -45.4506,
  -45.5933,
  -45.7326,
  -45.8693,
  -46.003,
  -46.1344,
  -46.263,
  -46.389,
  -46.5129,
  -46.6346,
  -46.7547,
  -46.874,
  -46.9926,
  -47.1107,
  -47.2276,
  -47.3434,
  -47.4573,
  -47.5724,
  -47.6892,
  -47.8088,
  -47.9317,
  -48.0585,
  -48.1894,
  -48.3244,
  -48.4636,
  -48.6059,
  -48.7509,
  -48.8976,
  -49.0459,
  -49.1959,
  -49.3482,
  -49.5038,
  -49.6625,
  -49.8265,
  -49.9945,
  -50.1663,
  -50.342,
  -50.5217,
  -50.7063,
  -50.8956,
  -51.0909,
  -51.293,
  -51.5036,
  -51.7246,
  -51.9567,
  -52.2006,
  -52.455,
  -52.7171,
  -52.9827,
  -53.247,
  -53.5037,
  -53.7499,
  -53.9796,
  -54.188,
  -54.3712,
  -54.5256,
  -54.6483,
  -54.7375,
  -54.7935,
  -54.8181,
  -54.8147,
  -54.7883,
  -54.7453,
  -54.6925,
  -54.6359,
  -54.5799,
  -54.5285,
  -54.4831,
  -54.4444,
  -54.4104,
  -54.382,
  -54.3569,
  -54.3341,
  -54.3125,
  -54.2914,
  -54.2713,
  -54.2525,
  -54.236,
  -54.2225,
  -54.2132,
  -54.2085,
  -54.2087,
  -54.214,
  -54.2245,
  -54.2403,
  -54.2621,
  -54.2909,
  -54.3273,
  -54.3717,
  -54.4225,
  -54.4808,
  -54.5438,
  -54.6094,
  -54.6751,
  -54.7389,
  -54.7986,
  -54.8531,
  -54.9004,
  -54.9397,
  -54.9706,
  -54.9928,
  -55.0062,
  -55.0101,
  -55.0036,
  -54.9857,
  -54.9564,
  -54.916,
  -54.8654,
  -54.8059,
  -54.7392,
  -54.6657,
  -54.5883,
  -54.506,
  -54.4187,
  -54.326,
  -54.2282,
  -54.1262,
  -54.0213,
  -53.9147,
  -53.8077,
  -53.7024,
  -53.6007,
  -53.5039,
  -53.4132,
  -53.3281,
  -53.2491,
  -53.176,
  -53.1082,
  -53.0457,
  -52.9881,
  -52.9357,
  -52.8881,
  -52.845,
  -52.8062,
  -52.77,
  -52.7383,
  -52.7096,
  -52.6836,
  -52.6599,
  -52.6378,
  -52.617,
  -52.5969,
  -52.5769,
  -52.5563,
  -52.5349,
  -52.5128,
  -52.4901,
  -52.4667,
  -52.4419,
  -52.4148,
  -52.3854,
  -52.353,
  -52.3178,
  -52.28,
  -52.2399,
  -52.198,
  -52.1549,
  -52.1107,
  -52.0656,
  -52.0195,
  -51.9716,
  -51.9246,
  -51.8776,
  -51.8307,
  -51.7831,
  -51.7342,
  -51.6837,
  -51.6307,
  -51.575,
  -51.5161,
  -51.4538,
  -51.3886,
  -51.3205,
  -51.2498,
  -51.1773,
  -51.1041,
  -51.0305,
  -50.9574,
  -50.8848,
  -50.813,
  -50.7418,
  -50.6708,
  -50.5994,
  -50.5266,
  -50.4518,
  -50.3743,
  -50.2934,
  -50.2092,
  -50.1219,
  -50.0317,
  -49.9386,
  -49.8458,
  -49.7537,
  -49.6636,
  -49.5753,
  -49.4889,
  -49.4041,
  -49.3204,
  -49.2375,
  -49.1554,
  -49.0744,
  -48.9949,
  -48.9168,
  -48.8405,
  -48.7665,
  -48.6958,
  -48.6285,
  -48.5646,
  -48.5031,
  -48.4425,
  -48.381,
  -48.3169,
  -48.249,
  -48.1777,
  -48.1038,
  -48.0297,
  -47.9582,
  -47.8916,
  -47.8326,
  -47.784,
  -47.7476,
  -47.7249,
  -47.7165,
  -47.7223,
  -47.7409,
  -47.7709,
  -47.8096,
  -47.8576,
  -47.9113,
  -47.9681,
  -48.0254,
  -48.0805,
  -48.1312,
  -48.1763,
  -48.2158,
  -48.2502,
  -48.2807,
  -48.3085,
  -48.3364,
  -48.3667,
  -48.402,
  -48.4438,
  -48.4934,
  -48.5511,
  -48.6159,
  -48.6856,
  -48.7574,
  -48.8289,
  -48.898,
  -48.9629,
  -49.0231,
  -49.0788,
  -49.131,
  -49.1808,
  -49.2304,
  -49.2812,
  -49.3353,
  -49.3942,
  -49.4583,
  -49.5281,
  -49.6042,
  -49.6878,
  -49.781,
  -39.2916,
  -39.4302,
  -39.5675,
  -39.7039,
  -39.8268,
  -39.9537,
  -40.0898,
  -40.2133,
  -40.3423,
  -40.4604,
  -40.5847,
  -40.7022,
  -40.8449,
  -41.0073,
  -41.1688,
  -41.3102,
  -41.4782,
  -41.6572,
  -41.8325,
  -42.0037,
  -42.1716,
  -42.3377,
  -42.5014,
  -42.664,
  -42.8287,
  -42.9957,
  -43.1633,
  -43.3311,
  -43.499,
  -43.666,
  -43.8324,
  -43.9971,
  -44.1585,
  -44.3186,
  -44.4765,
  -44.6315,
  -44.783,
  -44.9308,
  -45.075,
  -45.2162,
  -45.3541,
  -45.4895,
  -45.6226,
  -45.7533,
  -45.8818,
  -46.0077,
  -46.1314,
  -46.2525,
  -46.3712,
  -46.4898,
  -46.6074,
  -46.7241,
  -46.8395,
  -46.9538,
  -47.0674,
  -47.1812,
  -47.2967,
  -47.4149,
  -47.5365,
  -47.6621,
  -47.7919,
  -47.926,
  -48.0639,
  -48.2054,
  -48.3485,
  -48.4952,
  -48.6432,
  -48.7937,
  -48.9462,
  -49.1023,
  -49.2625,
  -49.4265,
  -49.5947,
  -49.7669,
  -49.943,
  -50.1234,
  -50.3086,
  -50.4991,
  -50.6962,
  -50.9009,
  -51.1151,
  -51.3409,
  -51.5785,
  -51.8301,
  -52.0932,
  -52.3644,
  -52.6388,
  -52.9108,
  -53.1745,
  -53.4244,
  -53.655,
  -53.8615,
  -54.0399,
  -54.187,
  -54.3,
  -54.3776,
  -54.4205,
  -54.4312,
  -54.4137,
  -54.3737,
  -54.3171,
  -54.2537,
  -54.1882,
  -54.1255,
  -54.0689,
  -54.0201,
  -53.9783,
  -53.9432,
  -53.9126,
  -53.8852,
  -53.8599,
  -53.8357,
  -53.8122,
  -53.7898,
  -53.7693,
  -53.751,
  -53.7362,
  -53.7256,
  -53.7202,
  -53.7199,
  -53.724,
  -53.7345,
  -53.7503,
  -53.7721,
  -53.8002,
  -53.8353,
  -53.8775,
  -53.9265,
  -53.9808,
  -54.0389,
  -54.0987,
  -54.1579,
  -54.2146,
  -54.2673,
  -54.3145,
  -54.3551,
  -54.3887,
  -54.4147,
  -54.433,
  -54.4432,
  -54.4445,
  -54.4347,
  -54.4154,
  -54.3851,
  -54.3446,
  -54.2942,
  -54.2354,
  -54.1699,
  -54.0993,
  -54.0247,
  -53.9458,
  -53.8622,
  -53.7743,
  -53.6822,
  -53.5864,
  -53.488,
  -53.3879,
  -53.2878,
  -53.1892,
  -53.093,
  -53.0013,
  -52.9142,
  -52.8327,
  -52.7553,
  -52.6842,
  -52.6178,
  -52.5561,
  -52.4991,
  -52.4468,
  -52.3993,
  -52.3559,
  -52.3162,
  -52.2805,
  -52.2476,
  -52.2178,
  -52.1903,
  -52.1647,
  -52.1408,
  -52.1179,
  -52.0957,
  -52.0736,
  -52.0511,
  -52.0282,
  -52.0049,
  -51.9817,
  -51.9583,
  -51.9344,
  -51.9098,
  -51.8828,
  -51.8524,
  -51.8204,
  -51.7858,
  -51.7487,
  -51.7097,
  -51.669,
  -51.6264,
  -51.5821,
  -51.5364,
  -51.4896,
  -51.4425,
  -51.3954,
  -51.3484,
  -51.3013,
  -51.2533,
  -51.2043,
  -51.1535,
  -51.1006,
  -51.0458,
  -50.9885,
  -50.9289,
  -50.8671,
  -50.803,
  -50.7377,
  -50.6717,
  -50.6054,
  -50.5392,
  -50.4732,
  -50.4065,
  -50.3409,
  -50.2751,
  -50.2081,
  -50.1391,
  -50.0674,
  -49.9926,
  -49.914,
  -49.8315,
  -49.7456,
  -49.6569,
  -49.5664,
  -49.4755,
  -49.3849,
  -49.2963,
  -49.21,
  -49.1253,
  -49.0422,
  -48.9599,
  -48.8782,
  -48.7972,
  -48.7172,
  -48.6385,
  -48.5609,
  -48.4844,
  -48.4095,
  -48.337,
  -48.2671,
  -48.1997,
  -48.1332,
  -48.0667,
  -47.9982,
  -47.9268,
  -47.8516,
  -47.772,
  -47.6921,
  -47.6132,
  -47.5384,
  -47.4704,
  -47.4116,
  -47.3645,
  -47.331,
  -47.3116,
  -47.3068,
  -47.3159,
  -47.3378,
  -47.3708,
  -47.4131,
  -47.4626,
  -47.5175,
  -47.5744,
  -47.6314,
  -47.6855,
  -47.7347,
  -47.7786,
  -47.8167,
  -47.8499,
  -47.8795,
  -47.9069,
  -47.9349,
  -47.9656,
  -48.0017,
  -48.045,
  -48.0969,
  -48.1574,
  -48.2255,
  -48.2991,
  -48.3755,
  -48.4517,
  -48.5256,
  -48.5955,
  -48.6613,
  -48.7229,
  -48.7812,
  -48.8376,
  -48.8942,
  -48.9529,
  -49.0146,
  -49.083,
  -49.1577,
  -49.2391,
  -49.3278,
  -49.4253,
  -49.5333,
  -39.1563,
  -39.2953,
  -39.428,
  -39.5552,
  -39.6809,
  -39.8078,
  -39.9275,
  -40.04,
  -40.1633,
  -40.2774,
  -40.3816,
  -40.4932,
  -40.619,
  -40.7813,
  -40.9347,
  -41.0613,
  -41.2261,
  -41.4023,
  -41.5747,
  -41.7418,
  -41.9066,
  -42.0675,
  -42.2262,
  -42.384,
  -42.5434,
  -42.7037,
  -42.8653,
  -43.0266,
  -43.1891,
  -43.3508,
  -43.5122,
  -43.6719,
  -43.8301,
  -43.9865,
  -44.1408,
  -44.2928,
  -44.441,
  -44.5861,
  -44.7283,
  -44.8674,
  -45.0037,
  -45.1383,
  -45.2694,
  -45.3991,
  -45.5266,
  -45.6516,
  -45.7742,
  -45.8942,
  -46.0125,
  -46.13,
  -46.2465,
  -46.3616,
  -46.4757,
  -46.5886,
  -46.7011,
  -46.8139,
  -46.9281,
  -47.0447,
  -47.1638,
  -47.2876,
  -47.4157,
  -47.5483,
  -47.6847,
  -47.8237,
  -47.9663,
  -48.1114,
  -48.2581,
  -48.4081,
  -48.5601,
  -48.7164,
  -48.8758,
  -49.0388,
  -49.2069,
  -49.379,
  -49.5548,
  -49.7353,
  -49.9198,
  -50.111,
  -50.3094,
  -50.5161,
  -50.7336,
  -50.9639,
  -51.2079,
  -51.4661,
  -51.7363,
  -52.0148,
  -52.2962,
  -52.5746,
  -52.8434,
  -53.0962,
  -53.3273,
  -53.5316,
  -53.7055,
  -53.8448,
  -53.947,
  -54.0125,
  -54.0416,
  -54.0379,
  -54.0056,
  -53.9516,
  -53.8833,
  -53.8087,
  -53.7341,
  -53.6649,
  -53.6036,
  -53.5514,
  -53.5074,
  -53.4705,
  -53.4384,
  -53.4093,
  -53.3822,
  -53.3561,
  -53.3308,
  -53.306,
  -53.2842,
  -53.2651,
  -53.2496,
  -53.2387,
  -53.2328,
  -53.2329,
  -53.2379,
  -53.2486,
  -53.2644,
  -53.286,
  -53.3133,
  -53.3468,
  -53.3865,
  -53.4319,
  -53.4818,
  -53.5347,
  -53.5885,
  -53.6412,
  -53.691,
  -53.7357,
  -53.776,
  -53.8104,
  -53.8385,
  -53.8601,
  -53.8743,
  -53.8814,
  -53.8802,
  -53.8691,
  -53.8487,
  -53.8176,
  -53.7769,
  -53.7274,
  -53.6698,
  -53.6065,
  -53.5382,
  -53.4663,
  -53.3909,
  -53.3115,
  -53.2289,
  -53.1423,
  -53.0531,
  -52.9603,
  -52.8674,
  -52.7747,
  -52.6825,
  -52.5915,
  -52.5044,
  -52.4212,
  -52.3428,
  -52.2688,
  -52.1989,
  -52.1338,
  -52.0731,
  -52.017,
  -51.9651,
  -51.9173,
  -51.8734,
  -51.8335,
  -51.7971,
  -51.763,
  -51.7318,
  -51.7031,
  -51.6761,
  -51.6506,
  -51.6259,
  -51.6019,
  -51.577,
  -51.5532,
  -51.5294,
  -51.5057,
  -51.4827,
  -51.4602,
  -51.4384,
  -51.416,
  -51.3915,
  -51.3652,
  -51.3366,
  -51.3055,
  -51.272,
  -51.2357,
  -51.1973,
  -51.1567,
  -51.114,
  -51.0695,
  -51.0234,
  -50.9765,
  -50.93,
  -50.8836,
  -50.8374,
  -50.7907,
  -50.743,
  -50.6944,
  -50.6445,
  -50.5924,
  -50.5394,
  -50.4847,
  -50.4284,
  -50.3704,
  -50.3114,
  -50.2514,
  -50.1914,
  -50.1309,
  -50.0704,
  -50.0097,
  -49.9483,
  -49.8864,
  -49.8229,
  -49.7568,
  -49.6877,
  -49.6147,
  -49.5381,
  -49.4574,
  -49.3734,
  -49.287,
  -49.1991,
  -49.1107,
  -49.0228,
  -48.9365,
  -48.8527,
  -48.7705,
  -48.6891,
  -48.6087,
  -48.5287,
  -48.4491,
  -48.3691,
  -48.2907,
  -48.2136,
  -48.1369,
  -48.0612,
  -47.9871,
  -47.9145,
  -47.8425,
  -47.7708,
  -47.698,
  -47.6224,
  -47.5434,
  -47.4612,
  -47.377,
  -47.2931,
  -47.2114,
  -47.136,
  -47.0693,
  -47.0133,
  -46.9702,
  -46.9411,
  -46.9264,
  -46.9255,
  -46.938,
  -46.9623,
  -46.9969,
  -47.04,
  -47.0894,
  -47.1433,
  -47.1987,
  -47.2533,
  -47.3053,
  -47.352,
  -47.3935,
  -47.4299,
  -47.4615,
  -47.4898,
  -47.5166,
  -47.544,
  -47.5737,
  -47.6099,
  -47.6542,
  -47.7077,
  -47.7703,
  -47.8415,
  -47.9187,
  -47.9993,
  -48.0801,
  -48.1586,
  -48.2335,
  -48.3044,
  -48.3716,
  -48.436,
  -48.4991,
  -48.5632,
  -48.6303,
  -48.7025,
  -48.7812,
  -48.8673,
  -48.9612,
  -49.0635,
  -49.1757,
  -49.2992,
  -39.0445,
  -39.1529,
  -39.2819,
  -39.4139,
  -39.5428,
  -39.6629,
  -39.7744,
  -39.8882,
  -39.9941,
  -40.0941,
  -40.1962,
  -40.3049,
  -40.4293,
  -40.5755,
  -40.714,
  -40.8366,
  -41.0026,
  -41.1655,
  -41.3295,
  -41.4909,
  -41.649,
  -41.8052,
  -41.9604,
  -42.1177,
  -42.274,
  -42.4296,
  -42.5846,
  -42.742,
  -42.9001,
  -43.0579,
  -43.2153,
  -43.3714,
  -43.526,
  -43.6791,
  -43.8308,
  -43.9797,
  -44.1256,
  -44.2677,
  -44.4078,
  -44.545,
  -44.68,
  -44.8129,
  -44.9435,
  -45.0719,
  -45.198,
  -45.3215,
  -45.4421,
  -45.5606,
  -45.6773,
  -45.7934,
  -45.9082,
  -46.0221,
  -46.1349,
  -46.2459,
  -46.3572,
  -46.4689,
  -46.5817,
  -46.6964,
  -46.8143,
  -46.9358,
  -47.0615,
  -47.1915,
  -47.3252,
  -47.4626,
  -47.6022,
  -47.7441,
  -47.8894,
  -48.038,
  -48.1889,
  -48.3439,
  -48.5014,
  -48.6642,
  -48.8317,
  -49.0026,
  -49.1784,
  -49.3586,
  -49.5441,
  -49.7358,
  -49.9351,
  -50.1437,
  -50.3635,
  -50.5973,
  -50.8456,
  -51.109,
  -51.3843,
  -51.668,
  -51.9548,
  -52.2369,
  -52.5093,
  -52.7643,
  -52.9954,
  -53.1973,
  -53.3661,
  -53.4979,
  -53.5908,
  -53.6438,
  -53.659,
  -53.6403,
  -53.5929,
  -53.5243,
  -53.4431,
  -53.3573,
  -53.2739,
  -53.1979,
  -53.1323,
  -53.0771,
  -53.0302,
  -52.9921,
  -52.959,
  -52.9289,
  -52.9006,
  -52.8732,
  -52.8468,
  -52.8222,
  -52.8,
  -52.7809,
  -52.7655,
  -52.7549,
  -52.7497,
  -52.7502,
  -52.7556,
  -52.7668,
  -52.7828,
  -52.8037,
  -52.8297,
  -52.861,
  -52.8967,
  -52.9381,
  -52.9831,
  -53.0305,
  -53.0783,
  -53.1246,
  -53.1679,
  -53.2071,
  -53.2412,
  -53.2699,
  -53.2928,
  -53.31,
  -53.3209,
  -53.3243,
  -53.3204,
  -53.3077,
  -53.2857,
  -53.2548,
  -53.2146,
  -53.1661,
  -53.1109,
  -53.0494,
  -52.9841,
  -52.915,
  -52.8426,
  -52.7678,
  -52.69,
  -52.6097,
  -52.5266,
  -52.442,
  -52.3561,
  -52.2698,
  -52.1837,
  -52.099,
  -52.0159,
  -51.9359,
  -51.8598,
  -51.7876,
  -51.7192,
  -51.655,
  -51.5953,
  -51.5399,
  -51.4885,
  -51.4409,
  -51.3969,
  -51.3556,
  -51.3183,
  -51.2838,
  -51.2515,
  -51.2216,
  -51.1935,
  -51.1666,
  -51.1405,
  -51.1149,
  -51.0895,
  -51.0649,
  -51.0408,
  -51.0172,
  -50.9949,
  -50.9738,
  -50.9539,
  -50.9336,
  -50.9123,
  -50.8895,
  -50.8644,
  -50.8365,
  -50.8062,
  -50.7731,
  -50.7372,
  -50.6988,
  -50.6584,
  -50.6147,
  -50.5707,
  -50.5257,
  -50.4805,
  -50.4358,
  -50.3911,
  -50.3462,
  -50.3006,
  -50.2542,
  -50.2071,
  -50.159,
  -50.11,
  -50.0594,
  -50.0076,
  -49.9546,
  -49.9003,
  -49.8453,
  -49.79,
  -49.7338,
  -49.6775,
  -49.6203,
  -49.5624,
  -49.5033,
  -49.4422,
  -49.3783,
  -49.3112,
  -49.2401,
  -49.1653,
  -49.0869,
  -49.0054,
  -48.9209,
  -48.8362,
  -48.7514,
  -48.6669,
  -48.5839,
  -48.5031,
  -48.4238,
  -48.345,
  -48.2665,
  -48.1884,
  -48.1103,
  -48.0324,
  -47.9547,
  -47.8776,
  -47.8008,
  -47.7242,
  -47.6482,
  -47.5724,
  -47.4961,
  -47.4188,
  -47.3393,
  -47.2567,
  -47.1708,
  -47.0829,
  -46.9949,
  -46.9087,
  -46.8269,
  -46.7537,
  -46.6905,
  -46.6398,
  -46.6026,
  -46.5796,
  -46.5703,
  -46.5736,
  -46.5892,
  -46.6143,
  -46.6494,
  -46.6918,
  -46.7395,
  -46.7908,
  -46.843,
  -46.8943,
  -46.9421,
  -46.9859,
  -47.0244,
  -47.0581,
  -47.0877,
  -47.1144,
  -47.1398,
  -47.1664,
  -47.1965,
  -47.2328,
  -47.2777,
  -47.3323,
  -47.3968,
  -47.4703,
  -47.5506,
  -47.6348,
  -47.7193,
  -47.8021,
  -47.8816,
  -47.9577,
  -48.0301,
  -48.1009,
  -48.171,
  -48.2431,
  -48.3191,
  -48.4015,
  -48.4912,
  -48.5896,
  -48.6968,
  -48.8138,
  -48.9411,
  -49.0803,
  -38.9287,
  -39.0391,
  -39.148,
  -39.2756,
  -39.4082,
  -39.5241,
  -39.6347,
  -39.7383,
  -39.8327,
  -39.9236,
  -40.0323,
  -40.1472,
  -40.2612,
  -40.388,
  -40.5065,
  -40.6343,
  -40.7757,
  -40.9332,
  -41.0909,
  -41.2459,
  -41.3968,
  -41.5546,
  -41.7083,
  -41.8658,
  -42.021,
  -42.1726,
  -42.3246,
  -42.4769,
  -42.6302,
  -42.7849,
  -42.9394,
  -43.0915,
  -43.243,
  -43.3936,
  -43.5429,
  -43.6902,
  -43.8341,
  -43.9751,
  -44.1135,
  -44.2494,
  -44.3828,
  -44.514,
  -44.6429,
  -44.7695,
  -44.8936,
  -45.0148,
  -45.1332,
  -45.2485,
  -45.3636,
  -45.4777,
  -45.591,
  -45.7037,
  -45.8155,
  -45.9265,
  -46.037,
  -46.1472,
  -46.2579,
  -46.3704,
  -46.4856,
  -46.6042,
  -46.7268,
  -46.8536,
  -46.9841,
  -47.1176,
  -47.2531,
  -47.393,
  -47.5359,
  -47.6822,
  -47.832,
  -47.9857,
  -48.143,
  -48.3053,
  -48.4719,
  -48.6427,
  -48.8175,
  -48.9976,
  -49.183,
  -49.374,
  -49.5738,
  -49.7838,
  -50.0058,
  -50.2408,
  -50.4922,
  -50.7584,
  -51.0369,
  -51.3238,
  -51.6137,
  -51.8998,
  -52.1743,
  -52.4303,
  -52.6606,
  -52.8596,
  -53.0228,
  -53.1465,
  -53.2291,
  -53.2698,
  -53.271,
  -53.2372,
  -53.1744,
  -53.0904,
  -52.9959,
  -52.8992,
  -52.8071,
  -52.7248,
  -52.655,
  -52.597,
  -52.5496,
  -52.5106,
  -52.4768,
  -52.4462,
  -52.4174,
  -52.3895,
  -52.3627,
  -52.3378,
  -52.3157,
  -52.2973,
  -52.2829,
  -52.2735,
  -52.2695,
  -52.2699,
  -52.2767,
  -52.2884,
  -52.3042,
  -52.3242,
  -52.3487,
  -52.3774,
  -52.4105,
  -52.4476,
  -52.4878,
  -52.5295,
  -52.5714,
  -52.6116,
  -52.6487,
  -52.6818,
  -52.7103,
  -52.7337,
  -52.7522,
  -52.7651,
  -52.7724,
  -52.7729,
  -52.7655,
  -52.7512,
  -52.7285,
  -52.6975,
  -52.6584,
  -52.6121,
  -52.5595,
  -52.5016,
  -52.4396,
  -52.3743,
  -52.3061,
  -52.2353,
  -52.1621,
  -52.0871,
  -52.0104,
  -51.9322,
  -51.853,
  -51.773,
  -51.6927,
  -51.6128,
  -51.5341,
  -51.4571,
  -51.3817,
  -51.3107,
  -51.2434,
  -51.1806,
  -51.1217,
  -51.0667,
  -51.0159,
  -50.9684,
  -50.9249,
  -50.8843,
  -50.8464,
  -50.8113,
  -50.7784,
  -50.7478,
  -50.7188,
  -50.6907,
  -50.6634,
  -50.6367,
  -50.6107,
  -50.5855,
  -50.5613,
  -50.5381,
  -50.5167,
  -50.497,
  -50.4788,
  -50.4599,
  -50.4415,
  -50.4217,
  -50.4,
  -50.3755,
  -50.348,
  -50.3177,
  -50.2849,
  -50.2495,
  -50.2119,
  -50.1721,
  -50.131,
  -50.0889,
  -50.0469,
  -50.005,
  -49.9627,
  -49.9203,
  -49.8771,
  -49.8337,
  -49.7893,
  -49.7442,
  -49.6982,
  -49.651,
  -49.6028,
  -49.5533,
  -49.5025,
  -49.451,
  -49.3987,
  -49.346,
  -49.2913,
  -49.2369,
  -49.1813,
  -49.1242,
  -49.0653,
  -49.0033,
  -48.9378,
  -48.8688,
  -48.796,
  -48.7203,
  -48.642,
  -48.562,
  -48.4813,
  -48.4007,
  -48.3207,
  -48.2416,
  -48.164,
  -48.088,
  -48.012,
  -47.936,
  -47.86,
  -47.7834,
  -47.7066,
  -47.6296,
  -47.5527,
  -47.4757,
  -47.3981,
  -47.3201,
  -47.2412,
  -47.1607,
  -47.0778,
  -46.9916,
  -46.9027,
  -46.8101,
  -46.7179,
  -46.6274,
  -46.5411,
  -46.4617,
  -46.3927,
  -46.3355,
  -46.2917,
  -46.2619,
  -46.2456,
  -46.2417,
  -46.2498,
  -46.268,
  -46.2949,
  -46.3294,
  -46.3701,
  -46.4151,
  -46.4627,
  -46.5108,
  -46.5575,
  -46.6011,
  -46.6409,
  -46.6759,
  -46.7066,
  -46.7337,
  -46.7588,
  -46.7828,
  -46.8084,
  -46.8381,
  -46.8745,
  -46.9197,
  -46.9752,
  -47.0411,
  -47.1161,
  -47.1982,
  -47.2847,
  -47.3724,
  -47.4587,
  -47.5426,
  -47.6231,
  -47.7009,
  -47.7778,
  -47.8545,
  -47.9354,
  -48.0209,
  -48.1138,
  -48.2155,
  -48.3267,
  -48.4481,
  -48.5798,
  -48.7226,
  -48.8776,
  -38.8133,
  -38.9238,
  -39.0305,
  -39.1605,
  -39.2835,
  -39.3967,
  -39.4997,
  -39.5917,
  -39.6792,
  -39.7831,
  -39.8891,
  -39.9909,
  -40.0937,
  -40.2125,
  -40.3202,
  -40.429,
  -40.561,
  -40.7054,
  -40.8589,
  -41.0035,
  -41.1571,
  -41.3153,
  -41.4708,
  -41.626,
  -41.7815,
  -41.9321,
  -42.079,
  -42.2284,
  -42.3775,
  -42.5281,
  -42.6806,
  -42.8308,
  -42.9806,
  -43.1293,
  -43.2771,
  -43.4232,
  -43.566,
  -43.7061,
  -43.8432,
  -43.9775,
  -44.1096,
  -44.2383,
  -44.3652,
  -44.4895,
  -44.6111,
  -44.7296,
  -44.8451,
  -44.9587,
  -45.0716,
  -45.1837,
  -45.2955,
  -45.4069,
  -45.5181,
  -45.6282,
  -45.7375,
  -45.8462,
  -45.9547,
  -46.0644,
  -46.1753,
  -46.2906,
  -46.4093,
  -46.5325,
  -46.6592,
  -46.7891,
  -46.9224,
  -47.0593,
  -47.1997,
  -47.344,
  -47.4925,
  -47.6449,
  -47.8015,
  -47.9628,
  -48.1287,
  -48.2991,
  -48.4739,
  -48.6521,
  -48.8367,
  -49.0277,
  -49.2279,
  -49.4382,
  -49.661,
  -49.8979,
  -50.1504,
  -50.4174,
  -50.6967,
  -50.9847,
  -51.2755,
  -51.5622,
  -51.8375,
  -52.0929,
  -52.3214,
  -52.5166,
  -52.674,
  -52.7885,
  -52.8606,
  -52.8888,
  -52.8757,
  -52.8267,
  -52.7487,
  -52.6511,
  -52.5438,
  -52.4365,
  -52.3361,
  -52.2481,
  -52.1744,
  -52.1138,
  -52.0653,
  -52.0254,
  -51.9917,
  -51.9608,
  -51.9319,
  -51.9039,
  -51.8762,
  -51.8513,
  -51.8299,
  -51.8126,
  -51.7998,
  -51.7922,
  -51.7903,
  -51.7937,
  -51.802,
  -51.8144,
  -51.8302,
  -51.8493,
  -51.8718,
  -51.8978,
  -51.9273,
  -51.96,
  -51.9951,
  -52.0315,
  -52.0677,
  -52.1021,
  -52.1325,
  -52.1602,
  -52.1837,
  -52.2025,
  -52.2166,
  -52.2258,
  -52.2299,
  -52.228,
  -52.2196,
  -52.2041,
  -52.1812,
  -52.1507,
  -52.1133,
  -52.0697,
  -52.0201,
  -51.9651,
  -51.9068,
  -51.8451,
  -51.7806,
  -51.7139,
  -51.6452,
  -51.5753,
  -51.503,
  -51.4307,
  -51.3574,
  -51.2829,
  -51.2079,
  -51.1323,
  -51.0572,
  -50.9828,
  -50.9101,
  -50.8402,
  -50.7739,
  -50.7118,
  -50.6537,
  -50.5995,
  -50.5492,
  -50.5022,
  -50.4587,
  -50.4181,
  -50.3801,
  -50.3445,
  -50.3112,
  -50.2802,
  -50.2508,
  -50.2222,
  -50.1932,
  -50.1658,
  -50.1394,
  -50.1141,
  -50.09,
  -50.0675,
  -50.0468,
  -50.0282,
  -50.0114,
  -49.9954,
  -49.9794,
  -49.9623,
  -49.9433,
  -49.9218,
  -49.8973,
  -49.87,
  -49.8401,
  -49.808,
  -49.7738,
  -49.7377,
  -49.7004,
  -49.6626,
  -49.6247,
  -49.5868,
  -49.5483,
  -49.5093,
  -49.4694,
  -49.428,
  -49.3866,
  -49.344,
  -49.3004,
  -49.2558,
  -49.21,
  -49.163,
  -49.1147,
  -49.0655,
  -49.0153,
  -48.9648,
  -48.9132,
  -48.8607,
  -48.807,
  -48.7516,
  -48.6941,
  -48.6339,
  -48.5704,
  -48.5037,
  -48.4334,
  -48.3609,
  -48.2865,
  -48.2108,
  -48.1348,
  -48.0591,
  -47.984,
  -47.9093,
  -47.8354,
  -47.7626,
  -47.6898,
  -47.6164,
  -47.5426,
  -47.4667,
  -47.3913,
  -47.3151,
  -47.2384,
  -47.1614,
  -47.083,
  -47.0032,
  -46.9214,
  -46.8368,
  -46.7485,
  -46.6566,
  -46.5617,
  -46.4655,
  -46.3704,
  -46.2791,
  -46.1948,
  -46.1198,
  -46.0563,
  -46.0065,
  -45.9708,
  -45.9488,
  -45.9393,
  -45.9411,
  -45.9531,
  -45.9733,
  -46.0005,
  -46.0338,
  -46.0718,
  -46.1133,
  -46.1568,
  -46.2004,
  -46.2426,
  -46.2819,
  -46.3173,
  -46.3486,
  -46.3765,
  -46.4013,
  -46.4245,
  -46.4468,
  -46.4722,
  -46.502,
  -46.5389,
  -46.5847,
  -46.6405,
  -46.7068,
  -46.7824,
  -46.8651,
  -46.9526,
  -47.0421,
  -47.131,
  -47.218,
  -47.3026,
  -47.3865,
  -47.4701,
  -47.5552,
  -47.6448,
  -47.7407,
  -47.8449,
  -47.959,
  -48.0836,
  -48.2192,
  -48.3661,
  -48.5242,
  -48.6936,
  -38.712,
  -38.8179,
  -38.9283,
  -39.045,
  -39.1669,
  -39.2749,
  -39.3638,
  -39.4641,
  -39.5593,
  -39.6549,
  -39.7531,
  -39.8461,
  -39.9498,
  -40.0519,
  -40.1529,
  -40.2528,
  -40.3745,
  -40.5151,
  -40.6478,
  -40.774,
  -40.9366,
  -41.0942,
  -41.2484,
  -41.4034,
  -41.5563,
  -41.7033,
  -41.8492,
  -41.9955,
  -42.143,
  -42.2907,
  -42.4391,
  -42.5877,
  -42.7349,
  -42.8827,
  -43.0295,
  -43.1746,
  -43.3157,
  -43.455,
  -43.5912,
  -43.7244,
  -43.8557,
  -43.9841,
  -44.1093,
  -44.2316,
  -44.3506,
  -44.4663,
  -44.579,
  -44.69,
  -44.8004,
  -44.9104,
  -45.0203,
  -45.1305,
  -45.2395,
  -45.3486,
  -45.4563,
  -45.563,
  -45.6691,
  -45.7758,
  -45.8842,
  -45.9954,
  -46.1101,
  -46.2286,
  -46.351,
  -46.4771,
  -46.6072,
  -46.7415,
  -46.8799,
  -47.0229,
  -47.1702,
  -47.3204,
  -47.476,
  -47.6363,
  -47.8014,
  -47.9712,
  -48.1454,
  -48.3238,
  -48.508,
  -48.6991,
  -48.8988,
  -49.1086,
  -49.3311,
  -49.5677,
  -49.8191,
  -50.0847,
  -50.3629,
  -50.6497,
  -50.9385,
  -51.224,
  -51.4976,
  -51.7507,
  -51.9758,
  -52.166,
  -52.3165,
  -52.4233,
  -52.4847,
  -52.5007,
  -52.4739,
  -52.4098,
  -52.3171,
  -52.2058,
  -52.0863,
  -51.9688,
  -51.8609,
  -51.7673,
  -51.6897,
  -51.6262,
  -51.5763,
  -51.5363,
  -51.5024,
  -51.4715,
  -51.4422,
  -51.4148,
  -51.3883,
  -51.3641,
  -51.3434,
  -51.3275,
  -51.3169,
  -51.312,
  -51.3129,
  -51.3189,
  -51.3293,
  -51.3429,
  -51.3592,
  -51.3777,
  -51.3984,
  -51.4204,
  -51.4461,
  -51.4746,
  -51.5048,
  -51.5361,
  -51.5669,
  -51.5961,
  -51.6225,
  -51.6453,
  -51.664,
  -51.6785,
  -51.6888,
  -51.6948,
  -51.6961,
  -51.692,
  -51.682,
  -51.6659,
  -51.6433,
  -51.6142,
  -51.5786,
  -51.5372,
  -51.49,
  -51.4391,
  -51.3843,
  -51.3259,
  -51.2649,
  -51.202,
  -51.1377,
  -51.0724,
  -51.0058,
  -50.9383,
  -50.87,
  -50.8004,
  -50.7297,
  -50.6579,
  -50.5857,
  -50.5137,
  -50.4429,
  -50.3743,
  -50.3088,
  -50.2471,
  -50.1897,
  -50.1362,
  -50.0865,
  -50.04,
  -49.9958,
  -49.9553,
  -49.9174,
  -49.8819,
  -49.8485,
  -49.8173,
  -49.788,
  -49.7593,
  -49.7316,
  -49.7038,
  -49.6775,
  -49.6525,
  -49.6288,
  -49.6069,
  -49.5871,
  -49.5694,
  -49.5535,
  -49.539,
  -49.5246,
  -49.5094,
  -49.4928,
  -49.4737,
  -49.4519,
  -49.4276,
  -49.4007,
  -49.3709,
  -49.3402,
  -49.3083,
  -49.2756,
  -49.2426,
  -49.2095,
  -49.1765,
  -49.1427,
  -49.108,
  -49.0719,
  -49.0347,
  -48.9962,
  -48.9561,
  -48.9146,
  -48.8717,
  -48.8276,
  -48.7822,
  -48.7356,
  -48.688,
  -48.6393,
  -48.5902,
  -48.5405,
  -48.4897,
  -48.4379,
  -48.3841,
  -48.3284,
  -48.2702,
  -48.2092,
  -48.1452,
  -48.0784,
  -48.0086,
  -47.9386,
  -47.8676,
  -47.7966,
  -47.7261,
  -47.6562,
  -47.5864,
  -47.5168,
  -47.4475,
  -47.3777,
  -47.3068,
  -47.2349,
  -47.162,
  -47.0879,
  -47.0125,
  -46.9363,
  -46.8592,
  -46.7805,
  -46.6993,
  -46.6149,
  -46.5268,
  -46.4343,
  -46.338,
  -46.2389,
  -46.1397,
  -46.0429,
  -45.9524,
  -45.8709,
  -45.8008,
  -45.7443,
  -45.7021,
  -45.6743,
  -45.6597,
  -45.6565,
  -45.6632,
  -45.6771,
  -45.6987,
  -45.7256,
  -45.7571,
  -45.7922,
  -45.8303,
  -45.8697,
  -45.909,
  -45.9469,
  -45.9819,
  -46.0133,
  -46.0412,
  -46.0663,
  -46.0893,
  -46.1119,
  -46.1351,
  -46.1608,
  -46.1921,
  -46.2304,
  -46.2769,
  -46.3326,
  -46.3985,
  -46.4738,
  -46.5559,
  -46.6427,
  -46.732,
  -46.8218,
  -46.911,
  -46.9994,
  -47.0884,
  -47.1785,
  -47.2726,
  -47.3714,
  -47.4784,
  -47.5945,
  -47.7214,
  -47.86,
  -48.0105,
  -48.1725,
  -48.3454,
  -48.5278,
  -38.6163,
  -38.715,
  -38.8295,
  -38.9388,
  -39.0579,
  -39.159,
  -39.2386,
  -39.3417,
  -39.4421,
  -39.5373,
  -39.6305,
  -39.7156,
  -39.8126,
  -39.9056,
  -39.9964,
  -40.0978,
  -40.2157,
  -40.3304,
  -40.4698,
  -40.6008,
  -40.739,
  -40.8982,
  -41.0504,
  -41.2006,
  -41.3457,
  -41.4889,
  -41.6342,
  -41.7794,
  -41.9246,
  -42.0698,
  -42.214,
  -42.3594,
  -42.5051,
  -42.6512,
  -42.7974,
  -42.942,
  -43.0837,
  -43.2222,
  -43.3579,
  -43.4906,
  -43.6209,
  -43.7481,
  -43.872,
  -43.9924,
  -44.109,
  -44.2221,
  -44.3317,
  -44.4403,
  -44.5482,
  -44.656,
  -44.7641,
  -44.8726,
  -44.9809,
  -45.0883,
  -45.1941,
  -45.2986,
  -45.4019,
  -45.5052,
  -45.6098,
  -45.7165,
  -45.8266,
  -45.9404,
  -46.0582,
  -46.1796,
  -46.3066,
  -46.4387,
  -46.5758,
  -46.718,
  -46.8647,
  -47.0152,
  -47.17,
  -47.3293,
  -47.4931,
  -47.6619,
  -47.835,
  -48.0129,
  -48.1966,
  -48.3871,
  -48.5859,
  -48.7947,
  -49.0146,
  -49.2489,
  -49.4975,
  -49.76,
  -50.0348,
  -50.3183,
  -50.6049,
  -50.887,
  -51.1567,
  -51.4056,
  -51.6254,
  -51.8092,
  -51.9518,
  -52.0495,
  -52.1,
  -52.1038,
  -52.0635,
  -51.9857,
  -51.8781,
  -51.7538,
  -51.6232,
  -51.4963,
  -51.3812,
  -51.2825,
  -51.2014,
  -51.1362,
  -51.0854,
  -51.0449,
  -51.0103,
  -50.9791,
  -50.9496,
  -50.9224,
  -50.8965,
  -50.8726,
  -50.8531,
  -50.839,
  -50.8311,
  -50.8293,
  -50.8325,
  -50.8418,
  -50.8548,
  -50.8705,
  -50.8878,
  -50.9061,
  -50.9255,
  -50.9464,
  -50.9689,
  -50.9933,
  -51.0192,
  -51.0456,
  -51.0716,
  -51.0961,
  -51.1178,
  -51.1362,
  -51.1507,
  -51.1611,
  -51.1685,
  -51.1717,
  -51.1705,
  -51.1637,
  -51.1527,
  -51.1366,
  -51.1145,
  -51.0864,
  -51.0526,
  -51.0137,
  -50.9707,
  -50.9232,
  -50.8717,
  -50.8168,
  -50.7591,
  -50.7003,
  -50.6399,
  -50.5783,
  -50.516,
  -50.4526,
  -50.3887,
  -50.3231,
  -50.2556,
  -50.1872,
  -50.1175,
  -50.0471,
  -49.978,
  -49.9107,
  -49.846,
  -49.7851,
  -49.7286,
  -49.676,
  -49.6267,
  -49.5809,
  -49.5379,
  -49.4979,
  -49.4603,
  -49.4247,
  -49.3918,
  -49.3609,
  -49.3322,
  -49.3044,
  -49.2769,
  -49.2501,
  -49.2243,
  -49.2001,
  -49.1767,
  -49.1555,
  -49.1366,
  -49.1199,
  -49.1037,
  -49.0901,
  -49.077,
  -49.0632,
  -49.0479,
  -49.0309,
  -49.0115,
  -48.9895,
  -48.9656,
  -48.9399,
  -48.9132,
  -48.8855,
  -48.8573,
  -48.8291,
  -48.8011,
  -48.7733,
  -48.7447,
  -48.7145,
  -48.6826,
  -48.6487,
  -48.6132,
  -48.5754,
  -48.5356,
  -48.4943,
  -48.4514,
  -48.4072,
  -48.3619,
  -48.3155,
  -48.2673,
  -48.2195,
  -48.1716,
  -48.1226,
  -48.0726,
  -48.0209,
  -47.9673,
  -47.9117,
  -47.8537,
  -47.7931,
  -47.7303,
  -47.6658,
  -47.6007,
  -47.535,
  -47.4694,
  -47.4043,
  -47.3397,
  -47.2751,
  -47.2099,
  -47.1439,
  -47.0769,
  -47.0084,
  -46.9385,
  -46.867,
  -46.7941,
  -46.7198,
  -46.6443,
  -46.5676,
  -46.4891,
  -46.4068,
  -46.3207,
  -46.2301,
  -46.1349,
  -46.0345,
  -45.9332,
  -45.8325,
  -45.736,
  -45.6474,
  -45.5696,
  -45.5049,
  -45.4552,
  -45.4202,
  -45.3993,
  -45.3908,
  -45.3928,
  -45.403,
  -45.4199,
  -45.442,
  -45.4682,
  -45.4975,
  -45.5295,
  -45.564,
  -45.5995,
  -45.6349,
  -45.6687,
  -45.6999,
  -45.7279,
  -45.7532,
  -45.7764,
  -45.799,
  -45.8218,
  -45.8464,
  -45.875,
  -45.9097,
  -45.9507,
  -45.9983,
  -46.0534,
  -46.1174,
  -46.19,
  -46.2696,
  -46.3538,
  -46.4412,
  -46.5307,
  -46.6211,
  -46.7128,
  -46.8056,
  -46.9028,
  -47.0052,
  -47.1144,
  -47.2324,
  -47.3611,
  -47.5016,
  -47.6546,
  -47.82,
  -47.9964,
  -48.1823,
  -48.3754,
  -38.5282,
  -38.6265,
  -38.7354,
  -38.8535,
  -38.9599,
  -39.0547,
  -39.1306,
  -39.2204,
  -39.3272,
  -39.423,
  -39.5124,
  -39.5981,
  -39.6846,
  -39.7658,
  -39.8637,
  -39.9568,
  -40.0688,
  -40.1794,
  -40.3037,
  -40.4384,
  -40.5707,
  -40.7195,
  -40.8646,
  -41.0068,
  -41.15,
  -41.2884,
  -41.4297,
  -41.5741,
  -41.7179,
  -41.8617,
  -42.0047,
  -42.1485,
  -42.2923,
  -42.4374,
  -42.5828,
  -42.7268,
  -42.8681,
  -43.0061,
  -43.1409,
  -43.2733,
  -43.4027,
  -43.528,
  -43.6507,
  -43.7695,
  -43.8841,
  -43.9952,
  -44.1036,
  -44.2103,
  -44.3161,
  -44.4215,
  -44.5276,
  -44.6338,
  -44.7397,
  -44.8447,
  -44.9481,
  -45.0498,
  -45.1503,
  -45.2493,
  -45.3501,
  -45.4527,
  -45.558,
  -45.6668,
  -45.7799,
  -45.8981,
  -46.022,
  -46.1522,
  -46.2892,
  -46.4309,
  -46.5777,
  -46.7283,
  -46.8826,
  -47.0403,
  -47.2026,
  -47.3698,
  -47.5405,
  -47.7177,
  -47.9007,
  -48.0903,
  -48.2878,
  -48.4945,
  -48.7124,
  -48.943,
  -49.1873,
  -49.4449,
  -49.7145,
  -49.993,
  -50.2742,
  -50.5507,
  -50.8144,
  -51.0568,
  -51.2695,
  -51.4456,
  -51.5786,
  -51.6666,
  -51.7063,
  -51.6983,
  -51.6453,
  -51.5546,
  -51.4358,
  -51.3,
  -51.1591,
  -51.0237,
  -50.9022,
  -50.7986,
  -50.7135,
  -50.6462,
  -50.5934,
  -50.5511,
  -50.5152,
  -50.4829,
  -50.4529,
  -50.4237,
  -50.3977,
  -50.3745,
  -50.356,
  -50.3437,
  -50.3384,
  -50.3402,
  -50.3485,
  -50.3616,
  -50.3782,
  -50.3965,
  -50.4156,
  -50.4347,
  -50.4537,
  -50.4731,
  -50.4932,
  -50.5146,
  -50.5368,
  -50.5591,
  -50.5807,
  -50.5998,
  -50.6173,
  -50.6312,
  -50.642,
  -50.6492,
  -50.6533,
  -50.6543,
  -50.6513,
  -50.6443,
  -50.6328,
  -50.6165,
  -50.595,
  -50.5686,
  -50.5366,
  -50.5,
  -50.4594,
  -50.4149,
  -50.3665,
  -50.3149,
  -50.2605,
  -50.2046,
  -50.1477,
  -50.0889,
  -50.0301,
  -49.9704,
  -49.9095,
  -49.8471,
  -49.7829,
  -49.717,
  -49.65,
  -49.5828,
  -49.516,
  -49.4503,
  -49.3871,
  -49.3274,
  -49.2716,
  -49.2199,
  -49.1713,
  -49.1259,
  -49.0835,
  -49.0437,
  -49.0064,
  -48.9718,
  -48.9396,
  -48.9097,
  -48.882,
  -48.8544,
  -48.8288,
  -48.8036,
  -48.7792,
  -48.7559,
  -48.7338,
  -48.7142,
  -48.6963,
  -48.6798,
  -48.6656,
  -48.6529,
  -48.6403,
  -48.6272,
  -48.6131,
  -48.597,
  -48.5794,
  -48.5595,
  -48.5381,
  -48.5152,
  -48.4915,
  -48.4676,
  -48.4439,
  -48.4204,
  -48.3973,
  -48.3743,
  -48.3505,
  -48.3251,
  -48.2963,
  -48.2657,
  -48.2326,
  -48.1968,
  -48.1587,
  -48.1185,
  -48.0768,
  -48.0339,
  -47.9897,
  -47.9448,
  -47.8992,
  -47.8533,
  -47.8072,
  -47.7605,
  -47.7129,
  -47.6639,
  -47.6131,
  -47.5605,
  -47.506,
  -47.4495,
  -47.3912,
  -47.3317,
  -47.2717,
  -47.2115,
  -47.1515,
  -47.0918,
  -47.0326,
  -46.9731,
  -46.9121,
  -46.8496,
  -46.7855,
  -46.7185,
  -46.6502,
  -46.5801,
  -46.5081,
  -46.435,
  -46.3606,
  -46.2845,
  -46.2064,
  -46.1244,
  -46.0376,
  -45.9459,
  -45.849,
  -45.7482,
  -45.6462,
  -45.5459,
  -45.4512,
  -45.3658,
  -45.2924,
  -45.2334,
  -45.1895,
  -45.1605,
  -45.1451,
  -45.1411,
  -45.1464,
  -45.1586,
  -45.1761,
  -45.1977,
  -45.2225,
  -45.2494,
  -45.2787,
  -45.3096,
  -45.3415,
  -45.3735,
  -45.4042,
  -45.4324,
  -45.4579,
  -45.4812,
  -45.5041,
  -45.5261,
  -45.5507,
  -45.5781,
  -45.6107,
  -45.6493,
  -45.6931,
  -45.742,
  -45.7971,
  -45.8592,
  -45.9286,
  -46.0037,
  -46.0842,
  -46.1687,
  -46.2569,
  -46.3479,
  -46.4424,
  -46.5414,
  -46.646,
  -46.7575,
  -46.877,
  -47.0066,
  -47.1479,
  -47.302,
  -47.469,
  -47.648,
  -47.8372,
  -48.0334,
  -48.2349,
  -38.4497,
  -38.5491,
  -38.6584,
  -38.7687,
  -38.8697,
  -38.9562,
  -39.0407,
  -39.1188,
  -39.2136,
  -39.3062,
  -39.3979,
  -39.4851,
  -39.5681,
  -39.6478,
  -39.7344,
  -39.8354,
  -39.9369,
  -40.0426,
  -40.1606,
  -40.2812,
  -40.4067,
  -40.5464,
  -40.6866,
  -40.8255,
  -40.9654,
  -41.1033,
  -41.2413,
  -41.3814,
  -41.5255,
  -41.6706,
  -41.8139,
  -41.9556,
  -42.0987,
  -42.2416,
  -42.3856,
  -42.5276,
  -42.6688,
  -42.8054,
  -42.9399,
  -43.0713,
  -43.1997,
  -43.3247,
  -43.4461,
  -43.5631,
  -43.6759,
  -43.7853,
  -43.8922,
  -43.9969,
  -44.1009,
  -44.2046,
  -44.3085,
  -44.4114,
  -44.5147,
  -44.6167,
  -44.7171,
  -44.8161,
  -44.9132,
  -45.0095,
  -45.1062,
  -45.2043,
  -45.3048,
  -45.4088,
  -45.5178,
  -45.6329,
  -45.7543,
  -45.8837,
  -46.0198,
  -46.1618,
  -46.3083,
  -46.4591,
  -46.6125,
  -46.7688,
  -46.9292,
  -47.0939,
  -47.2639,
  -47.4394,
  -47.6209,
  -47.8087,
  -48.0039,
  -48.2077,
  -48.4218,
  -48.6476,
  -48.8863,
  -49.1379,
  -49.4009,
  -49.6711,
  -49.9448,
  -50.2135,
  -50.4691,
  -50.7032,
  -50.9073,
  -51.0746,
  -51.1996,
  -51.278,
  -51.3076,
  -51.2886,
  -51.2246,
  -51.1231,
  -50.9935,
  -50.8478,
  -50.6978,
  -50.5546,
  -50.4271,
  -50.3181,
  -50.2279,
  -50.157,
  -50.101,
  -50.0561,
  -50.0181,
  -49.9839,
  -49.9521,
  -49.9226,
  -49.8957,
  -49.8725,
  -49.8549,
  -49.8442,
  -49.8415,
  -49.8466,
  -49.8591,
  -49.8764,
  -49.8968,
  -49.9188,
  -49.9403,
  -49.9612,
  -49.9803,
  -49.9993,
  -50.0181,
  -50.0371,
  -50.0563,
  -50.0753,
  -50.0933,
  -50.1096,
  -50.1234,
  -50.1339,
  -50.1417,
  -50.1464,
  -50.1479,
  -50.1468,
  -50.1423,
  -50.1344,
  -50.1224,
  -50.1057,
  -50.0841,
  -50.0581,
  -50.0275,
  -49.9913,
  -49.9525,
  -49.9101,
  -49.8646,
  -49.8157,
  -49.7646,
  -49.7116,
  -49.6576,
  -49.6033,
  -49.5479,
  -49.4913,
  -49.4335,
  -49.3739,
  -49.3124,
  -49.2494,
  -49.1849,
  -49.1201,
  -49.0554,
  -48.9923,
  -48.9312,
  -48.8731,
  -48.8186,
  -48.7678,
  -48.719,
  -48.6746,
  -48.6327,
  -48.5933,
  -48.5567,
  -48.5224,
  -48.4912,
  -48.4626,
  -48.4364,
  -48.4117,
  -48.388,
  -48.3652,
  -48.3429,
  -48.3215,
  -48.3017,
  -48.2839,
  -48.2674,
  -48.2524,
  -48.2387,
  -48.2262,
  -48.2139,
  -48.2013,
  -48.1878,
  -48.1728,
  -48.1561,
  -48.1379,
  -48.1174,
  -48.0968,
  -48.0759,
  -48.0551,
  -48.035,
  -48.0155,
  -47.9965,
  -47.9775,
  -47.9578,
  -47.9361,
  -47.912,
  -47.8843,
  -47.8535,
  -47.8195,
  -47.7829,
  -47.7442,
  -47.7038,
  -47.662,
  -47.6192,
  -47.5761,
  -47.5328,
  -47.4894,
  -47.446,
  -47.4022,
  -47.3576,
  -47.3119,
  -47.2644,
  -47.2154,
  -47.1648,
  -47.1116,
  -47.0584,
  -47.0043,
  -46.9497,
  -46.895,
  -46.8408,
  -46.7868,
  -46.7326,
  -46.6778,
  -46.6208,
  -46.5617,
  -46.5001,
  -46.4361,
  -46.3697,
  -46.3008,
  -46.2305,
  -46.1588,
  -46.0857,
  -46.0108,
  -45.9336,
  -45.8528,
  -45.7666,
  -45.6751,
  -45.5783,
  -45.4782,
  -45.3771,
  -45.279,
  -45.1874,
  -45.106,
  -45.0375,
  -44.9836,
  -44.9446,
  -44.9203,
  -44.9084,
  -44.9074,
  -44.9132,
  -44.9253,
  -44.9421,
  -44.9625,
  -44.985,
  -45.0094,
  -45.0358,
  -45.0637,
  -45.0925,
  -45.121,
  -45.1488,
  -45.1746,
  -45.1988,
  -45.2216,
  -45.2449,
  -45.2696,
  -45.2972,
  -45.3285,
  -45.3653,
  -45.4073,
  -45.4537,
  -45.5042,
  -45.5595,
  -45.6199,
  -45.686,
  -45.7573,
  -45.8334,
  -45.9147,
  -46.0013,
  -46.0934,
  -46.1904,
  -46.2951,
  -46.4078,
  -46.5287,
  -46.6584,
  -46.8003,
  -46.9543,
  -47.121,
  -47.3002,
  -47.4904,
  -47.6888,
  -47.8924,
  -48.0973,
  -38.3845,
  -38.4837,
  -38.5863,
  -38.6877,
  -38.7839,
  -38.8731,
  -38.9587,
  -39.0411,
  -39.1264,
  -39.2058,
  -39.2917,
  -39.3799,
  -39.4624,
  -39.5403,
  -39.623,
  -39.7176,
  -39.8153,
  -39.9206,
  -40.0298,
  -40.143,
  -40.2636,
  -40.3936,
  -40.5269,
  -40.661,
  -40.7952,
  -40.9307,
  -41.0675,
  -41.2064,
  -41.3475,
  -41.4937,
  -41.6374,
  -41.7794,
  -41.9219,
  -42.0639,
  -42.2054,
  -42.3468,
  -42.487,
  -42.6228,
  -42.7557,
  -42.8859,
  -43.0135,
  -43.137,
  -43.2567,
  -43.3721,
  -43.4831,
  -43.591,
  -43.6953,
  -43.7988,
  -43.9013,
  -44.003,
  -44.1049,
  -44.2062,
  -44.3065,
  -44.4057,
  -44.5029,
  -44.5981,
  -44.6919,
  -44.7847,
  -44.8772,
  -44.9708,
  -45.0667,
  -45.1665,
  -45.2708,
  -45.383,
  -45.5029,
  -45.6311,
  -45.7672,
  -45.9101,
  -46.0577,
  -46.2083,
  -46.3607,
  -46.5151,
  -46.6727,
  -46.8347,
  -47.0018,
  -47.1748,
  -47.3539,
  -47.5393,
  -47.7316,
  -47.9306,
  -48.1401,
  -48.3601,
  -48.5923,
  -48.8366,
  -49.0919,
  -49.3546,
  -49.6189,
  -49.878,
  -50.1236,
  -50.3476,
  -50.5419,
  -50.7001,
  -50.816,
  -50.8853,
  -50.9057,
  -50.8775,
  -50.8045,
  -50.6931,
  -50.555,
  -50.4013,
  -50.2439,
  -50.0944,
  -49.9607,
  -49.846,
  -49.7516,
  -49.6759,
  -49.6152,
  -49.5658,
  -49.5237,
  -49.486,
  -49.4513,
  -49.4193,
  -49.3905,
  -49.3665,
  -49.3492,
  -49.3401,
  -49.3396,
  -49.3471,
  -49.3628,
  -49.3843,
  -49.4094,
  -49.4351,
  -49.4602,
  -49.4837,
  -49.5054,
  -49.5255,
  -49.5438,
  -49.5615,
  -49.5786,
  -49.595,
  -49.6102,
  -49.6233,
  -49.6337,
  -49.6416,
  -49.6465,
  -49.6489,
  -49.6487,
  -49.6456,
  -49.6389,
  -49.6297,
  -49.6171,
  -49.5997,
  -49.578,
  -49.5519,
  -49.5218,
  -49.4878,
  -49.4498,
  -49.4092,
  -49.3656,
  -49.3194,
  -49.2712,
  -49.221,
  -49.1698,
  -49.118,
  -49.0656,
  -49.0123,
  -48.9573,
  -48.9006,
  -48.8419,
  -48.7816,
  -48.7192,
  -48.6572,
  -48.5954,
  -48.5351,
  -48.4766,
  -48.4209,
  -48.3682,
  -48.3185,
  -48.2717,
  -48.2283,
  -48.187,
  -48.1485,
  -48.1124,
  -48.0792,
  -48.049,
  -48.0219,
  -47.9974,
  -47.9752,
  -47.9542,
  -47.9343,
  -47.915,
  -47.8967,
  -47.8796,
  -47.8639,
  -47.8497,
  -47.8354,
  -47.8228,
  -47.8105,
  -47.7984,
  -47.786,
  -47.7727,
  -47.7582,
  -47.7424,
  -47.7251,
  -47.7069,
  -47.6881,
  -47.6691,
  -47.6507,
  -47.6333,
  -47.6168,
  -47.6008,
  -47.5848,
  -47.5681,
  -47.5492,
  -47.5277,
  -47.5027,
  -47.4738,
  -47.4414,
  -47.4062,
  -47.3688,
  -47.3298,
  -47.2896,
  -47.2488,
  -47.207,
  -47.1665,
  -47.1263,
  -47.0863,
  -47.0462,
  -47.0052,
  -46.9633,
  -46.9201,
  -46.875,
  -46.8286,
  -46.7811,
  -46.7328,
  -46.6841,
  -46.6352,
  -46.5863,
  -46.5378,
  -46.4891,
  -46.44,
  -46.3895,
  -46.3366,
  -46.2803,
  -46.2211,
  -46.1593,
  -46.0946,
  -46.0275,
  -45.9589,
  -45.8888,
  -45.8175,
  -45.7447,
  -45.6691,
  -45.5901,
  -45.5055,
  -45.4145,
  -45.3198,
  -45.2217,
  -45.1234,
  -45.029,
  -44.9418,
  -44.8652,
  -44.8018,
  -44.7525,
  -44.7175,
  -44.6961,
  -44.6862,
  -44.6859,
  -44.6924,
  -44.7033,
  -44.7182,
  -44.7361,
  -44.756,
  -44.778,
  -44.8014,
  -44.8264,
  -44.8522,
  -44.878,
  -44.9035,
  -44.9279,
  -44.9513,
  -44.9747,
  -44.9994,
  -45.0266,
  -45.0577,
  -45.0935,
  -45.1336,
  -45.1787,
  -45.2276,
  -45.2803,
  -45.3359,
  -45.3948,
  -45.4576,
  -45.5254,
  -45.5982,
  -45.6768,
  -45.7632,
  -45.8556,
  -45.9573,
  -46.0681,
  -46.1886,
  -46.3195,
  -46.4613,
  -46.6146,
  -46.7798,
  -46.9572,
  -47.1462,
  -47.3441,
  -47.5478,
  -47.7536,
  -47.9581,
  -38.3265,
  -38.4231,
  -38.5188,
  -38.6142,
  -38.7067,
  -38.7959,
  -38.8796,
  -38.9603,
  -39.0403,
  -39.1206,
  -39.1976,
  -39.2813,
  -39.3628,
  -39.4395,
  -39.5181,
  -39.6094,
  -39.7078,
  -39.8065,
  -39.9109,
  -40.0189,
  -40.1351,
  -40.2573,
  -40.3836,
  -40.5122,
  -40.6426,
  -40.7727,
  -40.9089,
  -41.0466,
  -41.1857,
  -41.3293,
  -41.4757,
  -41.6187,
  -41.762,
  -41.9042,
  -42.0447,
  -42.1829,
  -42.3218,
  -42.4567,
  -42.5881,
  -42.7169,
  -42.8418,
  -42.9638,
  -43.0817,
  -43.1951,
  -43.3046,
  -43.4108,
  -43.5147,
  -43.6171,
  -43.7179,
  -43.8179,
  -43.9176,
  -44.0162,
  -44.1135,
  -44.2095,
  -44.3036,
  -44.3956,
  -44.4848,
  -44.5738,
  -44.6624,
  -44.7517,
  -44.8434,
  -44.9394,
  -45.0417,
  -45.1515,
  -45.2703,
  -45.3979,
  -45.5341,
  -45.6767,
  -45.8242,
  -45.974,
  -46.1249,
  -46.2769,
  -46.4312,
  -46.5887,
  -46.7524,
  -46.9222,
  -47.098,
  -47.2795,
  -47.4679,
  -47.6632,
  -47.8667,
  -48.0806,
  -48.3056,
  -48.5422,
  -48.7885,
  -49.0413,
  -49.2947,
  -49.5422,
  -49.7764,
  -49.9892,
  -50.1734,
  -50.3209,
  -50.4284,
  -50.49,
  -50.503,
  -50.4678,
  -50.3886,
  -50.2727,
  -50.1288,
  -49.9697,
  -49.8072,
  -49.6524,
  -49.5124,
  -49.3907,
  -49.2897,
  -49.2071,
  -49.1396,
  -49.0837,
  -49.0357,
  -48.9923,
  -48.9519,
  -48.9163,
  -48.8847,
  -48.8587,
  -48.8409,
  -48.8324,
  -48.8339,
  -48.8447,
  -48.8635,
  -48.8886,
  -48.9174,
  -48.9478,
  -48.9769,
  -49.0034,
  -49.0279,
  -49.0498,
  -49.0687,
  -49.086,
  -49.1019,
  -49.1156,
  -49.1273,
  -49.138,
  -49.1459,
  -49.1511,
  -49.1538,
  -49.1542,
  -49.1525,
  -49.148,
  -49.1409,
  -49.1305,
  -49.1165,
  -49.0984,
  -49.0761,
  -49.0493,
  -49.019,
  -48.9852,
  -48.9483,
  -48.9084,
  -48.8666,
  -48.8225,
  -48.7768,
  -48.7296,
  -48.6802,
  -48.6311,
  -48.5815,
  -48.5311,
  -48.4793,
  -48.4255,
  -48.3698,
  -48.3126,
  -48.2545,
  -48.1962,
  -48.1381,
  -48.081,
  -48.0256,
  -47.9726,
  -47.9222,
  -47.874,
  -47.8289,
  -47.7861,
  -47.7462,
  -47.7082,
  -47.6731,
  -47.6405,
  -47.6115,
  -47.5862,
  -47.5632,
  -47.5438,
  -47.5261,
  -47.5095,
  -47.4942,
  -47.4796,
  -47.466,
  -47.4535,
  -47.4414,
  -47.4302,
  -47.4191,
  -47.4075,
  -47.3958,
  -47.3833,
  -47.3699,
  -47.3559,
  -47.3404,
  -47.3237,
  -47.3061,
  -47.2884,
  -47.271,
  -47.2542,
  -47.2386,
  -47.2241,
  -47.21,
  -47.1958,
  -47.1809,
  -47.163,
  -47.1431,
  -47.1198,
  -47.0928,
  -47.0618,
  -47.0279,
  -46.9919,
  -46.9544,
  -46.9162,
  -46.8777,
  -46.8394,
  -46.8023,
  -46.7661,
  -46.7302,
  -46.6944,
  -46.658,
  -46.6204,
  -46.5817,
  -46.5413,
  -46.4995,
  -46.4563,
  -46.4129,
  -46.3694,
  -46.3261,
  -46.283,
  -46.2399,
  -46.1965,
  -46.1521,
  -46.1058,
  -46.0564,
  -46.0021,
  -45.9454,
  -45.8858,
  -45.8233,
  -45.7582,
  -45.6916,
  -45.6236,
  -45.5543,
  -45.4841,
  -45.411,
  -45.3342,
  -45.2523,
  -45.165,
  -45.0736,
  -44.9794,
  -44.8855,
  -44.7959,
  -44.7141,
  -44.6429,
  -44.5846,
  -44.5397,
  -44.5077,
  -44.488,
  -44.4782,
  -44.4768,
  -44.4812,
  -44.4897,
  -44.5016,
  -44.5164,
  -44.5337,
  -44.553,
  -44.574,
  -44.5966,
  -44.6198,
  -44.6437,
  -44.6673,
  -44.6907,
  -44.7143,
  -44.7379,
  -44.7647,
  -44.7949,
  -44.8291,
  -44.8686,
  -44.913,
  -44.9606,
  -45.012,
  -45.0657,
  -45.1216,
  -45.179,
  -45.2391,
  -45.3044,
  -45.3756,
  -45.454,
  -45.5413,
  -45.6383,
  -45.7451,
  -45.8643,
  -45.9931,
  -46.1348,
  -46.2882,
  -46.4534,
  -46.6281,
  -46.8137,
  -47.008,
  -47.2088,
  -47.4125,
  -47.6155,
  -47.8144,
  -38.2696,
  -38.3638,
  -38.4541,
  -38.5448,
  -38.6337,
  -38.7192,
  -38.8014,
  -38.8798,
  -38.9574,
  -39.036,
  -39.1124,
  -39.191,
  -39.2724,
  -39.3491,
  -39.4263,
  -39.5107,
  -39.6059,
  -39.7024,
  -39.8035,
  -39.9054,
  -40.0182,
  -40.1354,
  -40.2558,
  -40.379,
  -40.5039,
  -40.6329,
  -40.7666,
  -40.9036,
  -41.0423,
  -41.1832,
  -41.3263,
  -41.4724,
  -41.6167,
  -41.7592,
  -41.8986,
  -42.0346,
  -42.1712,
  -42.3052,
  -42.4347,
  -42.5617,
  -42.6859,
  -42.8061,
  -42.9226,
  -43.0341,
  -43.1418,
  -43.2463,
  -43.3485,
  -43.4493,
  -43.5486,
  -43.647,
  -43.7448,
  -43.84,
  -43.9347,
  -44.0278,
  -44.1186,
  -44.2078,
  -44.2948,
  -44.38,
  -44.4645,
  -44.5498,
  -44.6377,
  -44.7307,
  -44.8307,
  -44.9392,
  -45.0569,
  -45.1838,
  -45.3192,
  -45.4601,
  -45.606,
  -45.7539,
  -45.9024,
  -46.0516,
  -46.2024,
  -46.3571,
  -46.5168,
  -46.6822,
  -46.8536,
  -47.0308,
  -47.2139,
  -47.4037,
  -47.6015,
  -47.8084,
  -48.0256,
  -48.253,
  -48.4891,
  -48.7293,
  -48.9703,
  -49.2051,
  -49.4267,
  -49.6277,
  -49.8013,
  -49.9414,
  -50.0412,
  -50.0968,
  -50.1052,
  -50.0666,
  -49.985,
  -49.8668,
  -49.7213,
  -49.5597,
  -49.3937,
  -49.2342,
  -49.0882,
  -48.9582,
  -48.8479,
  -48.7561,
  -48.6792,
  -48.6138,
  -48.5578,
  -48.5066,
  -48.4609,
  -48.4198,
  -48.3842,
  -48.3552,
  -48.3355,
  -48.3266,
  -48.3286,
  -48.3409,
  -48.3622,
  -48.3903,
  -48.4227,
  -48.4569,
  -48.4901,
  -48.5197,
  -48.5466,
  -48.5703,
  -48.5911,
  -48.6083,
  -48.6232,
  -48.6362,
  -48.6465,
  -48.6548,
  -48.6606,
  -48.6643,
  -48.665,
  -48.6637,
  -48.6606,
  -48.6552,
  -48.6468,
  -48.6352,
  -48.6198,
  -48.6007,
  -48.5774,
  -48.5494,
  -48.5173,
  -48.4831,
  -48.4462,
  -48.4074,
  -48.3669,
  -48.3245,
  -48.281,
  -48.2367,
  -48.1914,
  -48.1452,
  -48.0983,
  -48.0508,
  -48.0021,
  -47.9517,
  -47.8993,
  -47.8457,
  -47.7911,
  -47.7368,
  -47.6828,
  -47.6297,
  -47.5779,
  -47.528,
  -47.4801,
  -47.4331,
  -47.3897,
  -47.3484,
  -47.3093,
  -47.2723,
  -47.2378,
  -47.2063,
  -47.1785,
  -47.155,
  -47.135,
  -47.1188,
  -47.1047,
  -47.0921,
  -47.0807,
  -47.0706,
  -47.0609,
  -47.0519,
  -47.0427,
  -47.0341,
  -47.0246,
  -47.0143,
  -47.0027,
  -46.9906,
  -46.9771,
  -46.963,
  -46.9474,
  -46.9301,
  -46.9132,
  -46.8962,
  -46.8797,
  -46.8641,
  -46.8495,
  -46.8361,
  -46.8229,
  -46.8096,
  -46.7952,
  -46.7793,
  -46.7604,
  -46.7383,
  -46.7126,
  -46.6833,
  -46.651,
  -46.6165,
  -46.5808,
  -46.5445,
  -46.5087,
  -46.4738,
  -46.44,
  -46.408,
  -46.3769,
  -46.346,
  -46.3146,
  -46.2818,
  -46.2478,
  -46.2121,
  -46.174,
  -46.1358,
  -46.097,
  -46.0583,
  -46.0203,
  -45.9825,
  -45.9447,
  -45.9061,
  -45.8659,
  -45.8234,
  -45.7777,
  -45.7277,
  -45.6738,
  -45.6168,
  -45.5568,
  -45.4944,
  -45.43,
  -45.3652,
  -45.299,
  -45.2315,
  -45.161,
  -45.0872,
  -45.0091,
  -44.9254,
  -44.838,
  -44.7489,
  -44.6605,
  -44.5766,
  -44.5007,
  -44.4352,
  -44.3817,
  -44.3404,
  -44.311,
  -44.2918,
  -44.2813,
  -44.2766,
  -44.2782,
  -44.2833,
  -44.2914,
  -44.3028,
  -44.3173,
  -44.3342,
  -44.353,
  -44.3733,
  -44.395,
  -44.4174,
  -44.4401,
  -44.463,
  -44.4872,
  -44.5134,
  -44.5425,
  -44.5754,
  -44.613,
  -44.6553,
  -44.7019,
  -44.7528,
  -44.8061,
  -44.8606,
  -44.9161,
  -44.9729,
  -45.0326,
  -45.097,
  -45.1686,
  -45.2491,
  -45.3401,
  -45.4439,
  -45.5593,
  -45.6885,
  -45.8296,
  -45.9825,
  -46.1458,
  -46.319,
  -46.5006,
  -46.6897,
  -46.8842,
  -47.0819,
  -47.2797,
  -47.4742,
  -47.6635,
  -38.2122,
  -38.3025,
  -38.3908,
  -38.4779,
  -38.5624,
  -38.6472,
  -38.7282,
  -38.8052,
  -38.8796,
  -38.9569,
  -39.0314,
  -39.1094,
  -39.1882,
  -39.2656,
  -39.3422,
  -39.426,
  -39.5127,
  -39.6062,
  -39.7043,
  -39.8044,
  -39.9125,
  -40.0257,
  -40.1421,
  -40.2618,
  -40.3834,
  -40.509,
  -40.6413,
  -40.7761,
  -40.9135,
  -41.0527,
  -41.1937,
  -41.3361,
  -41.4828,
  -41.6255,
  -41.7647,
  -41.9008,
  -42.0354,
  -42.1678,
  -42.2966,
  -42.4228,
  -42.5451,
  -42.6636,
  -42.7778,
  -42.8875,
  -42.9934,
  -43.0952,
  -43.1957,
  -43.2944,
  -43.3921,
  -43.489,
  -43.5847,
  -43.6791,
  -43.7717,
  -43.8624,
  -43.9507,
  -44.0364,
  -44.1201,
  -44.2021,
  -44.2829,
  -44.3645,
  -44.4493,
  -44.539,
  -44.6373,
  -44.7448,
  -44.8616,
  -44.9877,
  -45.1215,
  -45.2612,
  -45.4044,
  -45.5491,
  -45.6941,
  -45.8398,
  -45.9871,
  -46.1376,
  -46.2932,
  -46.4534,
  -46.6191,
  -46.7902,
  -46.9662,
  -47.1503,
  -47.3415,
  -47.5415,
  -47.7504,
  -47.9681,
  -48.1928,
  -48.4208,
  -48.6481,
  -48.8683,
  -49.0762,
  -49.2652,
  -49.429,
  -49.5604,
  -49.6544,
  -49.7059,
  -49.7126,
  -49.674,
  -49.5938,
  -49.4771,
  -49.3338,
  -49.1733,
  -49.0065,
  -48.8437,
  -48.692,
  -48.5543,
  -48.4333,
  -48.3292,
  -48.2398,
  -48.1629,
  -48.0968,
  -48.0361,
  -47.9823,
  -47.9342,
  -47.8932,
  -47.86,
  -47.8376,
  -47.8267,
  -47.8268,
  -47.8395,
  -47.862,
  -47.892,
  -47.9271,
  -47.9644,
  -48.0012,
  -48.0351,
  -48.0653,
  -48.0915,
  -48.1131,
  -48.1307,
  -48.1454,
  -48.1569,
  -48.1656,
  -48.1715,
  -48.1761,
  -48.1787,
  -48.1781,
  -48.1756,
  -48.1713,
  -48.1638,
  -48.1545,
  -48.1416,
  -48.1249,
  -48.1042,
  -48.0793,
  -48.0502,
  -48.0178,
  -47.9828,
  -47.9455,
  -47.907,
  -47.868,
  -47.8275,
  -47.7861,
  -47.7444,
  -47.7021,
  -47.6595,
  -47.6159,
  -47.5716,
  -47.5261,
  -47.4788,
  -47.4303,
  -47.3795,
  -47.3288,
  -47.2787,
  -47.2291,
  -47.1804,
  -47.1326,
  -47.0862,
  -47.0412,
  -46.9976,
  -46.9565,
  -46.9167,
  -46.8785,
  -46.8426,
  -46.8093,
  -46.7786,
  -46.7521,
  -46.7298,
  -46.7121,
  -46.6984,
  -46.6875,
  -46.679,
  -46.6721,
  -46.6659,
  -46.6605,
  -46.6556,
  -46.6492,
  -46.6431,
  -46.6358,
  -46.6271,
  -46.6165,
  -46.6045,
  -46.591,
  -46.5764,
  -46.5608,
  -46.5445,
  -46.5279,
  -46.5119,
  -46.496,
  -46.4811,
  -46.4676,
  -46.4546,
  -46.4417,
  -46.4283,
  -46.414,
  -46.3983,
  -46.3799,
  -46.3586,
  -46.3344,
  -46.3068,
  -46.2763,
  -46.2437,
  -46.2097,
  -46.1747,
  -46.1415,
  -46.1098,
  -46.0801,
  -46.0523,
  -46.0261,
  -46.0003,
  -45.9744,
  -45.9472,
  -45.9183,
  -45.8876,
  -45.8551,
  -45.8213,
  -45.7871,
  -45.7529,
  -45.7194,
  -45.6865,
  -45.6533,
  -45.6192,
  -45.583,
  -45.5441,
  -45.502,
  -45.4557,
  -45.4052,
  -45.3515,
  -45.2947,
  -45.2355,
  -45.1746,
  -45.1127,
  -45.0501,
  -44.9855,
  -44.9182,
  -44.8482,
  -44.7724,
  -44.6928,
  -44.6107,
  -44.5274,
  -44.4455,
  -44.3681,
  -44.2985,
  -44.2387,
  -44.1898,
  -44.1518,
  -44.1237,
  -44.1045,
  -44.0925,
  -44.0859,
  -44.0839,
  -44.0854,
  -44.0899,
  -44.0982,
  -44.1096,
  -44.1242,
  -44.1412,
  -44.1601,
  -44.1807,
  -44.2024,
  -44.2246,
  -44.248,
  -44.2733,
  -44.3013,
  -44.3325,
  -44.3675,
  -44.407,
  -44.4514,
  -44.5002,
  -44.5524,
  -44.607,
  -44.6626,
  -44.719,
  -44.7769,
  -44.838,
  -44.9047,
  -44.9795,
  -45.0643,
  -45.1628,
  -45.2757,
  -45.4028,
  -45.5439,
  -45.6971,
  -45.8607,
  -46.033,
  -46.2119,
  -46.3959,
  -46.5836,
  -46.7725,
  -46.9611,
  -47.1475,
  -47.3284,
  -47.5032,
  -38.1549,
  -38.2435,
  -38.3302,
  -38.4134,
  -38.4959,
  -38.5768,
  -38.6565,
  -38.7342,
  -38.8063,
  -38.8822,
  -38.9564,
  -39.0335,
  -39.1102,
  -39.187,
  -39.2625,
  -39.3454,
  -39.4314,
  -39.5207,
  -39.6158,
  -39.7133,
  -39.8174,
  -39.9257,
  -40.0381,
  -40.1545,
  -40.2742,
  -40.4004,
  -40.5284,
  -40.6614,
  -40.7954,
  -40.9341,
  -41.0743,
  -41.2154,
  -41.3581,
  -41.5025,
  -41.6416,
  -41.778,
  -41.9113,
  -42.0432,
  -42.1715,
  -42.2958,
  -42.4172,
  -42.5345,
  -42.6471,
  -42.7551,
  -42.8593,
  -42.9602,
  -43.0586,
  -43.1548,
  -43.2502,
  -43.3448,
  -43.4384,
  -43.5309,
  -43.622,
  -43.7106,
  -43.7965,
  -43.8797,
  -43.9594,
  -44.038,
  -44.1159,
  -44.1949,
  -44.2775,
  -44.3667,
  -44.4638,
  -44.5701,
  -44.6852,
  -44.8092,
  -44.9406,
  -45.0769,
  -45.2161,
  -45.3564,
  -45.4974,
  -45.6389,
  -45.7816,
  -45.9283,
  -46.0791,
  -46.2337,
  -46.3931,
  -46.5576,
  -46.7281,
  -46.9054,
  -47.09,
  -47.2822,
  -47.4822,
  -47.6891,
  -47.9012,
  -48.1152,
  -48.3273,
  -48.5327,
  -48.7267,
  -48.9032,
  -49.0553,
  -49.1787,
  -49.2673,
  -49.3167,
  -49.3238,
  -49.2887,
  -49.2135,
  -49.1039,
  -48.9668,
  -48.8113,
  -48.647,
  -48.4833,
  -48.3265,
  -48.1801,
  -48.0476,
  -47.9296,
  -47.8257,
  -47.7338,
  -47.6547,
  -47.582,
  -47.5182,
  -47.4615,
  -47.4139,
  -47.3753,
  -47.3491,
  -47.3354,
  -47.3347,
  -47.3464,
  -47.3686,
  -47.3996,
  -47.436,
  -47.4752,
  -47.5142,
  -47.5507,
  -47.5835,
  -47.6113,
  -47.6336,
  -47.6516,
  -47.6655,
  -47.6752,
  -47.6822,
  -47.6871,
  -47.6894,
  -47.691,
  -47.6896,
  -47.6861,
  -47.6809,
  -47.6735,
  -47.6632,
  -47.6498,
  -47.6319,
  -47.6099,
  -47.5839,
  -47.5529,
  -47.5199,
  -47.484,
  -47.4464,
  -47.408,
  -47.3704,
  -47.3317,
  -47.2925,
  -47.2523,
  -47.213,
  -47.1734,
  -47.1335,
  -47.0925,
  -47.0504,
  -47.0068,
  -46.9619,
  -46.916,
  -46.8698,
  -46.8239,
  -46.7789,
  -46.7347,
  -46.6913,
  -46.6488,
  -46.6073,
  -46.5666,
  -46.5278,
  -46.4898,
  -46.4532,
  -46.4184,
  -46.3861,
  -46.3563,
  -46.3311,
  -46.3095,
  -46.2938,
  -46.2828,
  -46.2752,
  -46.2708,
  -46.268,
  -46.2664,
  -46.2649,
  -46.2639,
  -46.2621,
  -46.2589,
  -46.2538,
  -46.2464,
  -46.2365,
  -46.2244,
  -46.2107,
  -46.1957,
  -46.18,
  -46.1637,
  -46.1477,
  -46.1321,
  -46.1174,
  -46.1036,
  -46.0907,
  -46.0782,
  -46.0654,
  -46.0508,
  -46.0362,
  -46.0202,
  -46.0023,
  -45.9818,
  -45.9587,
  -45.9327,
  -45.9041,
  -45.8737,
  -45.8419,
  -45.8104,
  -45.78,
  -45.7518,
  -45.726,
  -45.7026,
  -45.6811,
  -45.6603,
  -45.6397,
  -45.618,
  -45.5944,
  -45.5687,
  -45.5408,
  -45.5118,
  -45.482,
  -45.4522,
  -45.4229,
  -45.3941,
  -45.365,
  -45.3347,
  -45.3024,
  -45.2673,
  -45.2278,
  -45.1858,
  -45.1398,
  -45.0903,
  -45.0378,
  -44.983,
  -44.9262,
  -44.8683,
  -44.8089,
  -44.7476,
  -44.6838,
  -44.6167,
  -44.5458,
  -44.4711,
  -44.3938,
  -44.3164,
  -44.2409,
  -44.1702,
  -44.1065,
  -44.0522,
  -44.0074,
  -43.9722,
  -43.9453,
  -43.9257,
  -43.9116,
  -43.9021,
  -43.8965,
  -43.8943,
  -43.8955,
  -43.9009,
  -43.9095,
  -43.9218,
  -43.9375,
  -43.9558,
  -43.9762,
  -43.9978,
  -44.0204,
  -44.0439,
  -44.0707,
  -44.1002,
  -44.1332,
  -44.1701,
  -44.2111,
  -44.2571,
  -44.3071,
  -44.3606,
  -44.4162,
  -44.4734,
  -44.5315,
  -44.592,
  -44.6572,
  -44.7294,
  -44.8114,
  -44.9062,
  -45.0156,
  -45.1412,
  -45.2818,
  -45.4358,
  -45.6007,
  -45.7734,
  -45.9516,
  -46.1322,
  -46.3137,
  -46.4945,
  -46.6726,
  -46.8474,
  -47.0175,
  -47.1818,
  -47.3394,
  -38.0967,
  -38.1852,
  -38.2705,
  -38.3514,
  -38.4295,
  -38.5068,
  -38.5849,
  -38.6647,
  -38.7397,
  -38.8134,
  -38.8867,
  -38.9633,
  -39.0392,
  -39.1133,
  -39.1903,
  -39.2714,
  -39.3556,
  -39.444,
  -39.536,
  -39.6311,
  -39.7295,
  -39.8325,
  -39.9416,
  -40.0551,
  -40.1737,
  -40.2967,
  -40.4234,
  -40.5547,
  -40.6886,
  -40.8244,
  -40.9639,
  -41.105,
  -41.2461,
  -41.3887,
  -41.527,
  -41.6629,
  -41.7966,
  -41.9286,
  -42.0571,
  -42.1821,
  -42.3036,
  -42.4205,
  -42.5317,
  -42.6382,
  -42.7406,
  -42.8397,
  -42.9357,
  -43.0294,
  -43.1218,
  -43.2138,
  -43.304,
  -43.3947,
  -43.4842,
  -43.5711,
  -43.6555,
  -43.7363,
  -43.814,
  -43.8898,
  -43.9652,
  -44.0422,
  -44.1236,
  -44.2117,
  -44.3081,
  -44.4128,
  -44.5262,
  -44.6473,
  -44.7735,
  -44.9049,
  -45.0386,
  -45.1736,
  -45.3097,
  -45.4475,
  -45.5877,
  -45.7306,
  -45.8763,
  -46.0251,
  -46.1773,
  -46.3343,
  -46.4976,
  -46.6678,
  -46.8453,
  -47.0297,
  -47.2203,
  -47.4154,
  -47.6126,
  -47.8113,
  -48.0074,
  -48.1971,
  -48.3762,
  -48.5394,
  -48.6816,
  -48.7973,
  -48.8812,
  -48.9292,
  -48.9389,
  -48.9096,
  -48.8429,
  -48.7434,
  -48.6161,
  -48.4695,
  -48.3103,
  -48.149,
  -47.9872,
  -47.8319,
  -47.6871,
  -47.5541,
  -47.4339,
  -47.3264,
  -47.2326,
  -47.1476,
  -47.0728,
  -47.0075,
  -46.9519,
  -46.9074,
  -46.8767,
  -46.8597,
  -46.8564,
  -46.8658,
  -46.8865,
  -46.9165,
  -46.9527,
  -46.9922,
  -47.031,
  -47.0688,
  -47.103,
  -47.132,
  -47.155,
  -47.1726,
  -47.1856,
  -47.1948,
  -47.2009,
  -47.2039,
  -47.2046,
  -47.2062,
  -47.2042,
  -47.2005,
  -47.1947,
  -47.1863,
  -47.1751,
  -47.1612,
  -47.1425,
  -47.1192,
  -47.0917,
  -47.058,
  -47.0237,
  -46.9873,
  -46.9495,
  -46.9113,
  -46.875,
  -46.8379,
  -46.8009,
  -46.7642,
  -46.7275,
  -46.6913,
  -46.6547,
  -46.6176,
  -46.5791,
  -46.5391,
  -46.4981,
  -46.4561,
  -46.4141,
  -46.3725,
  -46.3319,
  -46.2924,
  -46.2534,
  -46.2152,
  -46.1763,
  -46.1386,
  -46.1025,
  -46.0664,
  -46.0316,
  -45.9982,
  -45.967,
  -45.9381,
  -45.9142,
  -45.8951,
  -45.8811,
  -45.8723,
  -45.8679,
  -45.8668,
  -45.8679,
  -45.87,
  -45.8725,
  -45.875,
  -45.8764,
  -45.876,
  -45.8731,
  -45.8671,
  -45.8578,
  -45.8458,
  -45.8317,
  -45.8163,
  -45.7994,
  -45.7837,
  -45.7683,
  -45.7539,
  -45.7405,
  -45.728,
  -45.7162,
  -45.7043,
  -45.6919,
  -45.6784,
  -45.6636,
  -45.6477,
  -45.6304,
  -45.6111,
  -45.5894,
  -45.5649,
  -45.5386,
  -45.5104,
  -45.4812,
  -45.4525,
  -45.4251,
  -45.4004,
  -45.3784,
  -45.3594,
  -45.3425,
  -45.3268,
  -45.3115,
  -45.2952,
  -45.277,
  -45.2554,
  -45.2324,
  -45.2076,
  -45.1821,
  -45.1565,
  -45.1312,
  -45.1058,
  -45.0802,
  -45.0534,
  -45.0248,
  -44.9935,
  -44.959,
  -44.9215,
  -44.8805,
  -44.836,
  -44.7888,
  -44.7389,
  -44.687,
  -44.6332,
  -44.5777,
  -44.5197,
  -44.4588,
  -44.3949,
  -44.3277,
  -44.2574,
  -44.1852,
  -44.1134,
  -44.044,
  -43.9796,
  -43.9219,
  -43.8724,
  -43.8314,
  -43.7986,
  -43.7726,
  -43.7514,
  -43.7356,
  -43.7234,
  -43.7149,
  -43.7096,
  -43.708,
  -43.7105,
  -43.7169,
  -43.728,
  -43.7427,
  -43.7607,
  -43.7813,
  -43.8035,
  -43.8276,
  -43.8536,
  -43.8822,
  -43.9135,
  -43.9479,
  -43.986,
  -44.0283,
  -44.075,
  -44.126,
  -44.1804,
  -44.2377,
  -44.2968,
  -44.3589,
  -44.4241,
  -44.4966,
  -44.578,
  -44.6707,
  -44.777,
  -44.8995,
  -45.0396,
  -45.1953,
  -45.3626,
  -45.5377,
  -45.717,
  -45.8968,
  -46.0753,
  -46.2493,
  -46.418,
  -46.5807,
  -46.7374,
  -46.8879,
  -47.0327,
  -47.1698,
  -38.037,
  -38.1253,
  -38.2108,
  -38.2909,
  -38.3681,
  -38.4441,
  -38.5193,
  -38.5972,
  -38.6758,
  -38.7488,
  -38.8199,
  -38.8981,
  -38.972,
  -39.0441,
  -39.1201,
  -39.2019,
  -39.286,
  -39.372,
  -39.4627,
  -39.5576,
  -39.6538,
  -39.7498,
  -39.8529,
  -39.9614,
  -40.0773,
  -40.1977,
  -40.3227,
  -40.4527,
  -40.5855,
  -40.7201,
  -40.8583,
  -40.9986,
  -41.1414,
  -41.283,
  -41.421,
  -41.5572,
  -41.6917,
  -41.8251,
  -41.9546,
  -42.0808,
  -42.2028,
  -42.3195,
  -42.4303,
  -42.5361,
  -42.6361,
  -42.733,
  -42.8263,
  -42.9169,
  -43.006,
  -43.0948,
  -43.183,
  -43.2712,
  -43.3588,
  -43.4442,
  -43.5264,
  -43.6054,
  -43.6811,
  -43.7551,
  -43.8287,
  -43.9044,
  -43.9851,
  -44.0715,
  -44.1665,
  -44.2696,
  -44.3797,
  -44.4975,
  -44.6196,
  -44.7451,
  -44.8727,
  -45.0019,
  -45.1329,
  -45.2667,
  -45.4027,
  -45.541,
  -45.6816,
  -45.8244,
  -45.9698,
  -46.1193,
  -46.2739,
  -46.4366,
  -46.6061,
  -46.7816,
  -46.9615,
  -47.1443,
  -47.3287,
  -47.5122,
  -47.6922,
  -47.8657,
  -48.029,
  -48.1782,
  -48.3083,
  -48.4148,
  -48.4935,
  -48.5401,
  -48.5529,
  -48.5303,
  -48.473,
  -48.3859,
  -48.2712,
  -48.1354,
  -47.9859,
  -47.828,
  -47.6671,
  -47.5064,
  -47.3501,
  -47.2034,
  -47.0673,
  -46.9432,
  -46.8341,
  -46.7355,
  -46.6489,
  -46.574,
  -46.5106,
  -46.4597,
  -46.4244,
  -46.4021,
  -46.3953,
  -46.4018,
  -46.4192,
  -46.4465,
  -46.4802,
  -46.5179,
  -46.5567,
  -46.5936,
  -46.6278,
  -46.6565,
  -46.6794,
  -46.6963,
  -46.7084,
  -46.7166,
  -46.7211,
  -46.7226,
  -46.7221,
  -46.7226,
  -46.7204,
  -46.7162,
  -46.7091,
  -46.7003,
  -46.6887,
  -46.6742,
  -46.655,
  -46.631,
  -46.6022,
  -46.5676,
  -46.5328,
  -46.496,
  -46.4584,
  -46.4208,
  -46.3856,
  -46.3502,
  -46.3155,
  -46.2809,
  -46.2467,
  -46.213,
  -46.1797,
  -46.146,
  -46.1109,
  -46.0744,
  -46.036,
  -45.9981,
  -45.9602,
  -45.9228,
  -45.8866,
  -45.8514,
  -45.8171,
  -45.7833,
  -45.749,
  -45.7144,
  -45.6814,
  -45.6475,
  -45.6147,
  -45.5829,
  -45.5533,
  -45.5249,
  -45.5023,
  -45.4846,
  -45.4721,
  -45.465,
  -45.4634,
  -45.4653,
  -45.4697,
  -45.4752,
  -45.4813,
  -45.4857,
  -45.4903,
  -45.4917,
  -45.4907,
  -45.4855,
  -45.4763,
  -45.4645,
  -45.4502,
  -45.4349,
  -45.4192,
  -45.404,
  -45.39,
  -45.3775,
  -45.3658,
  -45.3552,
  -45.3449,
  -45.3345,
  -45.3231,
  -45.3102,
  -45.296,
  -45.2807,
  -45.2641,
  -45.246,
  -45.2259,
  -45.2036,
  -45.1795,
  -45.1542,
  -45.1269,
  -45.1015,
  -45.0777,
  -45.0566,
  -45.0388,
  -45.0238,
  -45.0115,
  -45.0005,
  -44.9901,
  -44.979,
  -44.966,
  -44.9504,
  -44.9322,
  -44.912,
  -44.8908,
  -44.8691,
  -44.8475,
  -44.8257,
  -44.8033,
  -44.78,
  -44.7547,
  -44.7271,
  -44.6969,
  -44.6642,
  -44.6281,
  -44.589,
  -44.5474,
  -44.503,
  -44.4562,
  -44.4072,
  -44.3556,
  -44.301,
  -44.2416,
  -44.1805,
  -44.1164,
  -44.05,
  -43.9821,
  -43.9153,
  -43.8514,
  -43.7927,
  -43.7408,
  -43.696,
  -43.6588,
  -43.6283,
  -43.6031,
  -43.5825,
  -43.5651,
  -43.5509,
  -43.5395,
  -43.5318,
  -43.5282,
  -43.5287,
  -43.5336,
  -43.5439,
  -43.5585,
  -43.577,
  -43.5985,
  -43.6223,
  -43.6485,
  -43.6765,
  -43.7069,
  -43.7395,
  -43.7744,
  -43.8131,
  -43.8558,
  -43.903,
  -43.9552,
  -44.0108,
  -44.0707,
  -44.1343,
  -44.2014,
  -44.2748,
  -44.3565,
  -44.4501,
  -44.5556,
  -44.6761,
  -44.8139,
  -44.9699,
  -45.1399,
  -45.3185,
  -45.5012,
  -45.6832,
  -45.8609,
  -46.0321,
  -46.1943,
  -46.3476,
  -46.4919,
  -46.6289,
  -46.7586,
  -46.8827,
  -47.0009,
  -37.9775,
  -38.0652,
  -38.1529,
  -38.2331,
  -38.3089,
  -38.3839,
  -38.4571,
  -38.5329,
  -38.6098,
  -38.6871,
  -38.7575,
  -38.8311,
  -38.9027,
  -38.977,
  -39.0549,
  -39.137,
  -39.2214,
  -39.3077,
  -39.3965,
  -39.4874,
  -39.5766,
  -39.6703,
  -39.7687,
  -39.8721,
  -39.9834,
  -40.1031,
  -40.2257,
  -40.3542,
  -40.4871,
  -40.621,
  -40.7576,
  -40.8976,
  -41.0416,
  -41.1867,
  -41.3244,
  -41.4598,
  -41.5951,
  -41.7306,
  -41.8617,
  -41.9885,
  -42.112,
  -42.2294,
  -42.3409,
  -42.4462,
  -42.5463,
  -42.6411,
  -42.7316,
  -42.8189,
  -42.9041,
  -42.9889,
  -43.0741,
  -43.1599,
  -43.2451,
  -43.3288,
  -43.4093,
  -43.4853,
  -43.5591,
  -43.6317,
  -43.7044,
  -43.7794,
  -43.8596,
  -43.946,
  -44.0398,
  -44.1402,
  -44.247,
  -44.3599,
  -44.4764,
  -44.5958,
  -44.7167,
  -44.8401,
  -44.9659,
  -45.0949,
  -45.2258,
  -45.3595,
  -45.4947,
  -45.6307,
  -45.7689,
  -45.9111,
  -46.0588,
  -46.2133,
  -46.374,
  -46.5398,
  -46.7086,
  -46.879,
  -47.0492,
  -47.2171,
  -47.3809,
  -47.5375,
  -47.6846,
  -47.8176,
  -47.9339,
  -48.0294,
  -48.1013,
  -48.1456,
  -48.1608,
  -48.1453,
  -48.1,
  -48.0259,
  -47.9253,
  -47.8034,
  -47.6653,
  -47.5148,
  -47.356,
  -47.1917,
  -47.0275,
  -46.8694,
  -46.7196,
  -46.5798,
  -46.4557,
  -46.3438,
  -46.2455,
  -46.1613,
  -46.0911,
  -46.0341,
  -45.9936,
  -45.9685,
  -45.9573,
  -45.959,
  -45.972,
  -45.9946,
  -46.0244,
  -46.0587,
  -46.0943,
  -46.1287,
  -46.1608,
  -46.1884,
  -46.2103,
  -46.2265,
  -46.2366,
  -46.2432,
  -46.2464,
  -46.2469,
  -46.2454,
  -46.2456,
  -46.2423,
  -46.238,
  -46.2316,
  -46.2229,
  -46.2109,
  -46.1957,
  -46.1758,
  -46.151,
  -46.1212,
  -46.0853,
  -46.0493,
  -46.0122,
  -45.9747,
  -45.9379,
  -45.904,
  -45.8702,
  -45.8357,
  -45.8033,
  -45.7716,
  -45.7401,
  -45.7091,
  -45.678,
  -45.6457,
  -45.6126,
  -45.5788,
  -45.5446,
  -45.5106,
  -45.4774,
  -45.4455,
  -45.4147,
  -45.3846,
  -45.3548,
  -45.3246,
  -45.2938,
  -45.2637,
  -45.2328,
  -45.2019,
  -45.172,
  -45.1435,
  -45.1168,
  -45.0944,
  -45.0772,
  -45.0657,
  -45.0598,
  -45.0603,
  -45.0644,
  -45.0716,
  -45.0805,
  -45.0897,
  -45.0972,
  -45.1041,
  -45.1077,
  -45.108,
  -45.1028,
  -45.0945,
  -45.083,
  -45.0684,
  -45.0526,
  -45.0375,
  -45.0241,
  -45.0115,
  -45.0012,
  -44.9922,
  -44.9842,
  -44.976,
  -44.9677,
  -44.9571,
  -44.9462,
  -44.9332,
  -44.9191,
  -44.9039,
  -44.8872,
  -44.8689,
  -44.8491,
  -44.8278,
  -44.8054,
  -44.7829,
  -44.7612,
  -44.7413,
  -44.7243,
  -44.7104,
  -44.6995,
  -44.6914,
  -44.6851,
  -44.6796,
  -44.6733,
  -44.6651,
  -44.6544,
  -44.6416,
  -44.6262,
  -44.6091,
  -44.5914,
  -44.5733,
  -44.5549,
  -44.5359,
  -44.5154,
  -44.4925,
  -44.4686,
  -44.4423,
  -44.4138,
  -44.3825,
  -44.3487,
  -44.3126,
  -44.2739,
  -44.2326,
  -44.1879,
  -44.14,
  -44.0887,
  -44.0339,
  -43.9752,
  -43.9134,
  -43.8498,
  -43.7855,
  -43.7231,
  -43.6644,
  -43.6111,
  -43.5644,
  -43.5242,
  -43.4903,
  -43.462,
  -43.4381,
  -43.4172,
  -43.399,
  -43.3833,
  -43.3704,
  -43.361,
  -43.3558,
  -43.3552,
  -43.3599,
  -43.3701,
  -43.3849,
  -43.4038,
  -43.4277,
  -43.4524,
  -43.4809,
  -43.5112,
  -43.5435,
  -43.5771,
  -43.6127,
  -43.6514,
  -43.6943,
  -43.7423,
  -43.7954,
  -43.8543,
  -43.9186,
  -43.9875,
  -44.0635,
  -44.1481,
  -44.243,
  -44.3496,
  -44.4693,
  -44.6057,
  -44.7607,
  -44.9317,
  -45.1139,
  -45.3008,
  -45.4872,
  -45.6675,
  -45.8384,
  -45.9982,
  -46.1454,
  -46.2806,
  -46.4051,
  -46.5211,
  -46.6303,
  -46.734,
  -46.8322,
  -37.919,
  -38.0087,
  -38.0956,
  -38.1743,
  -38.2526,
  -38.3279,
  -38.4018,
  -38.4757,
  -38.5498,
  -38.6265,
  -38.6943,
  -38.7642,
  -38.8377,
  -38.9132,
  -38.9925,
  -39.0743,
  -39.1583,
  -39.2439,
  -39.3299,
  -39.4177,
  -39.5045,
  -39.5935,
  -39.687,
  -39.7875,
  -39.8957,
  -40.0121,
  -40.1366,
  -40.2642,
  -40.3947,
  -40.5281,
  -40.6649,
  -40.8034,
  -40.947,
  -41.0915,
  -41.2317,
  -41.3695,
  -41.5054,
  -41.6429,
  -41.7767,
  -41.9068,
  -42.0319,
  -42.1508,
  -42.263,
  -42.3688,
  -42.4685,
  -42.5618,
  -42.6497,
  -42.7335,
  -42.8155,
  -42.8955,
  -42.9776,
  -43.0604,
  -43.1433,
  -43.2248,
  -43.3031,
  -43.3779,
  -43.4499,
  -43.5207,
  -43.5927,
  -43.6673,
  -43.747,
  -43.8325,
  -43.9241,
  -44.022,
  -44.1255,
  -44.2329,
  -44.3425,
  -44.4554,
  -44.5702,
  -44.6874,
  -44.8077,
  -44.9317,
  -45.0581,
  -45.1865,
  -45.3156,
  -45.4451,
  -45.576,
  -45.7104,
  -45.8501,
  -45.9959,
  -46.1473,
  -46.3027,
  -46.4602,
  -46.6169,
  -46.7728,
  -46.9254,
  -47.0725,
  -47.2124,
  -47.3415,
  -47.4591,
  -47.5603,
  -47.6426,
  -47.7056,
  -47.7465,
  -47.7621,
  -47.7526,
  -47.717,
  -47.6557,
  -47.5697,
  -47.4623,
  -47.3369,
  -47.1955,
  -47.0408,
  -46.8756,
  -46.708,
  -46.5422,
  -46.3809,
  -46.2306,
  -46.0964,
  -45.9731,
  -45.8654,
  -45.7736,
  -45.6982,
  -45.6372,
  -45.5928,
  -45.563,
  -45.5458,
  -45.5414,
  -45.5479,
  -45.5638,
  -45.5889,
  -45.6167,
  -45.6475,
  -45.6769,
  -45.7057,
  -45.7307,
  -45.751,
  -45.7663,
  -45.7766,
  -45.782,
  -45.7845,
  -45.7841,
  -45.7825,
  -45.7826,
  -45.7791,
  -45.7746,
  -45.7679,
  -45.7589,
  -45.7458,
  -45.7295,
  -45.7083,
  -45.6821,
  -45.65,
  -45.6115,
  -45.5743,
  -45.5361,
  -45.4986,
  -45.4622,
  -45.4299,
  -45.3969,
  -45.3648,
  -45.3338,
  -45.3036,
  -45.2734,
  -45.2439,
  -45.2143,
  -45.1845,
  -45.1542,
  -45.1242,
  -45.0935,
  -45.0635,
  -45.0346,
  -45.0072,
  -44.9805,
  -44.9549,
  -44.9284,
  -44.9025,
  -44.8762,
  -44.8507,
  -44.8225,
  -44.7944,
  -44.7668,
  -44.74,
  -44.7129,
  -44.692,
  -44.6756,
  -44.6648,
  -44.6602,
  -44.6635,
  -44.6697,
  -44.6794,
  -44.6912,
  -44.7033,
  -44.7132,
  -44.7213,
  -44.7257,
  -44.7269,
  -44.7223,
  -44.7127,
  -44.7005,
  -44.6863,
  -44.6707,
  -44.6564,
  -44.6436,
  -44.6332,
  -44.6252,
  -44.6192,
  -44.6145,
  -44.6102,
  -44.6043,
  -44.5973,
  -44.5887,
  -44.5782,
  -44.566,
  -44.552,
  -44.5373,
  -44.5213,
  -44.5045,
  -44.4864,
  -44.4676,
  -44.4491,
  -44.4317,
  -44.4161,
  -44.4034,
  -44.3937,
  -44.387,
  -44.3831,
  -44.3811,
  -44.3798,
  -44.3772,
  -44.3744,
  -44.3687,
  -44.3611,
  -44.3507,
  -44.3382,
  -44.3243,
  -44.3098,
  -44.2948,
  -44.2787,
  -44.2612,
  -44.2421,
  -44.2212,
  -44.1985,
  -44.1737,
  -44.1465,
  -44.1174,
  -44.0864,
  -44.0527,
  -44.0163,
  -43.9763,
  -43.9323,
  -43.8839,
  -43.8315,
  -43.7747,
  -43.7146,
  -43.6533,
  -43.5921,
  -43.5339,
  -43.4802,
  -43.432,
  -43.3901,
  -43.354,
  -43.3237,
  -43.2966,
  -43.2738,
  -43.2532,
  -43.2348,
  -43.2185,
  -43.2051,
  -43.1952,
  -43.1897,
  -43.1894,
  -43.195,
  -43.2062,
  -43.2224,
  -43.243,
  -43.2682,
  -43.2971,
  -43.3279,
  -43.3604,
  -43.3937,
  -43.4279,
  -43.4645,
  -43.5039,
  -43.5476,
  -43.5968,
  -43.653,
  -43.7165,
  -43.7866,
  -43.8642,
  -43.9505,
  -44.0471,
  -44.1553,
  -44.276,
  -44.4117,
  -44.5657,
  -44.7358,
  -44.9191,
  -45.1093,
  -45.3002,
  -45.4858,
  -45.66,
  -45.8205,
  -45.9652,
  -46.0949,
  -46.2107,
  -46.3155,
  -46.4116,
  -46.5003,
  -46.5848,
  -46.6647,
  -37.8658,
  -37.9548,
  -38.0402,
  -38.1211,
  -38.2003,
  -38.2766,
  -38.3521,
  -38.4244,
  -38.4962,
  -38.5689,
  -38.6349,
  -38.7041,
  -38.777,
  -38.8507,
  -38.9303,
  -39.0128,
  -39.0957,
  -39.1788,
  -39.2653,
  -39.3522,
  -39.4373,
  -39.5216,
  -39.6122,
  -39.7097,
  -39.8149,
  -39.9284,
  -40.0504,
  -40.1792,
  -40.3093,
  -40.4416,
  -40.5767,
  -40.7146,
  -40.8539,
  -40.9997,
  -41.1429,
  -41.2848,
  -41.4247,
  -41.5638,
  -41.7004,
  -41.8328,
  -41.9601,
  -42.0807,
  -42.1946,
  -42.3014,
  -42.4001,
  -42.4926,
  -42.5786,
  -42.66,
  -42.7386,
  -42.8168,
  -42.8955,
  -42.9758,
  -43.056,
  -43.1348,
  -43.2102,
  -43.2824,
  -43.3524,
  -43.4217,
  -43.4924,
  -43.5662,
  -43.6437,
  -43.7277,
  -43.817,
  -43.9118,
  -44.0113,
  -44.1137,
  -44.2188,
  -44.3254,
  -44.4342,
  -44.5455,
  -44.6602,
  -44.778,
  -44.8982,
  -45.0199,
  -45.1423,
  -45.2653,
  -45.3891,
  -45.5149,
  -45.6465,
  -45.7835,
  -45.9249,
  -46.0694,
  -46.215,
  -46.3599,
  -46.5017,
  -46.6386,
  -46.7694,
  -46.8911,
  -47.0026,
  -47.1011,
  -47.1853,
  -47.2534,
  -47.3057,
  -47.34,
  -47.3548,
  -47.3479,
  -47.32,
  -47.2699,
  -47.1971,
  -47.1038,
  -46.991,
  -46.86,
  -46.7134,
  -46.5526,
  -46.3854,
  -46.2155,
  -46.0473,
  -45.8886,
  -45.7453,
  -45.6139,
  -45.4984,
  -45.4016,
  -45.3227,
  -45.2592,
  -45.2114,
  -45.1766,
  -45.153,
  -45.1406,
  -45.1382,
  -45.1456,
  -45.1625,
  -45.186,
  -45.2119,
  -45.2358,
  -45.2602,
  -45.2821,
  -45.3003,
  -45.3146,
  -45.3235,
  -45.3287,
  -45.3303,
  -45.3291,
  -45.3271,
  -45.327,
  -45.324,
  -45.3176,
  -45.31,
  -45.3001,
  -45.2865,
  -45.2691,
  -45.2468,
  -45.2185,
  -45.1862,
  -45.147,
  -45.1103,
  -45.0727,
  -45.0345,
  -44.9983,
  -44.9666,
  -44.9337,
  -44.9024,
  -44.8718,
  -44.8425,
  -44.8123,
  -44.7832,
  -44.7544,
  -44.7253,
  -44.6973,
  -44.6706,
  -44.6437,
  -44.6178,
  -44.5928,
  -44.5695,
  -44.5469,
  -44.5255,
  -44.5043,
  -44.4825,
  -44.4598,
  -44.438,
  -44.4135,
  -44.3885,
  -44.3635,
  -44.3391,
  -44.3136,
  -44.2937,
  -44.2778,
  -44.2672,
  -44.2629,
  -44.267,
  -44.2742,
  -44.2853,
  -44.2974,
  -44.3108,
  -44.3219,
  -44.3312,
  -44.3371,
  -44.3381,
  -44.3346,
  -44.3259,
  -44.3144,
  -44.3014,
  -44.2877,
  -44.2752,
  -44.2655,
  -44.2579,
  -44.2532,
  -44.2506,
  -44.2497,
  -44.2492,
  -44.2476,
  -44.2438,
  -44.2381,
  -44.2304,
  -44.2204,
  -44.2094,
  -44.1968,
  -44.1835,
  -44.1699,
  -44.1558,
  -44.1406,
  -44.1265,
  -44.1135,
  -44.1028,
  -44.0945,
  -44.0893,
  -44.0867,
  -44.0865,
  -44.0886,
  -44.0917,
  -44.0949,
  -44.0969,
  -44.0962,
  -44.0939,
  -44.0884,
  -44.0807,
  -44.071,
  -44.06,
  -44.0482,
  -44.035,
  -44.0202,
  -44.0034,
  -43.9848,
  -43.9644,
  -43.9421,
  -43.9181,
  -43.8924,
  -43.8651,
  -43.8357,
  -43.8036,
  -43.7678,
  -43.7277,
  -43.682,
  -43.6323,
  -43.5779,
  -43.5207,
  -43.4621,
  -43.4041,
  -43.3496,
  -43.3004,
  -43.2572,
  -43.2198,
  -43.188,
  -43.161,
  -43.1376,
  -43.1164,
  -43.0968,
  -43.0785,
  -43.0624,
  -43.049,
  -43.0395,
  -43.0348,
  -43.0357,
  -43.0431,
  -43.0561,
  -43.0743,
  -43.0975,
  -43.1246,
  -43.1556,
  -43.1876,
  -43.2223,
  -43.2571,
  -43.2927,
  -43.3306,
  -43.3711,
  -43.416,
  -43.4681,
  -43.528,
  -43.5985,
  -43.6774,
  -43.7657,
  -43.8629,
  -43.9722,
  -44.0941,
  -44.2305,
  -44.3836,
  -44.5516,
  -44.733,
  -44.9239,
  -45.1176,
  -45.3071,
  -45.486,
  -45.65,
  -45.7963,
  -45.9246,
  -46.0361,
  -46.1334,
  -46.2197,
  -46.2979,
  -46.3702,
  -46.4372,
  -46.5004,
  -37.8233,
  -37.9113,
  -37.9962,
  -38.0773,
  -38.1568,
  -38.234,
  -38.3085,
  -38.3794,
  -38.4494,
  -38.5185,
  -38.5803,
  -38.6479,
  -38.7189,
  -38.7919,
  -38.8711,
  -38.952,
  -39.0333,
  -39.1153,
  -39.1999,
  -39.286,
  -39.3711,
  -39.4529,
  -39.5439,
  -39.6395,
  -39.7429,
  -39.8536,
  -39.9723,
  -40.0965,
  -40.2266,
  -40.3604,
  -40.4972,
  -40.6347,
  -40.7737,
  -40.9161,
  -41.0636,
  -41.208,
  -41.3508,
  -41.4925,
  -41.6302,
  -41.7651,
  -41.8942,
  -42.0167,
  -42.1325,
  -42.2405,
  -42.341,
  -42.4336,
  -42.5193,
  -42.5994,
  -42.6764,
  -42.7521,
  -42.8287,
  -42.9061,
  -42.9834,
  -43.0588,
  -43.1301,
  -43.1991,
  -43.2662,
  -43.3336,
  -43.4022,
  -43.4741,
  -43.5503,
  -43.6317,
  -43.7185,
  -43.8099,
  -43.9054,
  -44.0036,
  -44.1035,
  -44.2047,
  -44.3075,
  -44.413,
  -44.5214,
  -44.6316,
  -44.7448,
  -44.8594,
  -44.9743,
  -45.09,
  -45.2066,
  -45.3259,
  -45.4492,
  -45.5769,
  -45.7081,
  -45.8415,
  -45.9752,
  -46.107,
  -46.2346,
  -46.3559,
  -46.4695,
  -46.5732,
  -46.6649,
  -46.7427,
  -46.8085,
  -46.861,
  -46.9005,
  -46.9269,
  -46.9386,
  -46.9346,
  -46.9128,
  -46.8715,
  -46.8093,
  -46.7278,
  -46.6265,
  -46.5057,
  -46.3674,
  -46.2121,
  -46.0476,
  -45.8782,
  -45.709,
  -45.5455,
  -45.3977,
  -45.2604,
  -45.1397,
  -45.0372,
  -44.9517,
  -44.8872,
  -44.8386,
  -44.8009,
  -44.7717,
  -44.752,
  -44.7411,
  -44.739,
  -44.7463,
  -44.7627,
  -44.7796,
  -44.7982,
  -44.8171,
  -44.8362,
  -44.8532,
  -44.8659,
  -44.8747,
  -44.8791,
  -44.8813,
  -44.8803,
  -44.8784,
  -44.8788,
  -44.8762,
  -44.8716,
  -44.8644,
  -44.8531,
  -44.8367,
  -44.8176,
  -44.7926,
  -44.7622,
  -44.7304,
  -44.6909,
  -44.6547,
  -44.6174,
  -44.579,
  -44.5425,
  -44.5117,
  -44.4781,
  -44.4468,
  -44.4159,
  -44.386,
  -44.3536,
  -44.3224,
  -44.2925,
  -44.2649,
  -44.241,
  -44.2183,
  -44.1962,
  -44.1749,
  -44.1548,
  -44.1355,
  -44.1167,
  -44.0992,
  -44.0822,
  -44.0656,
  -44.0472,
  -44.0293,
  -44.0083,
  -43.9868,
  -43.9649,
  -43.9434,
  -43.919,
  -43.9006,
  -43.8858,
  -43.8759,
  -43.8718,
  -43.876,
  -43.8831,
  -43.8947,
  -43.9081,
  -43.9216,
  -43.9325,
  -43.9422,
  -43.9486,
  -43.9506,
  -43.9482,
  -43.9413,
  -43.9316,
  -43.9202,
  -43.9087,
  -43.8987,
  -43.8921,
  -43.8882,
  -43.8873,
  -43.8891,
  -43.8924,
  -43.8963,
  -43.8976,
  -43.8979,
  -43.8957,
  -43.8911,
  -43.8843,
  -43.876,
  -43.8666,
  -43.8568,
  -43.847,
  -43.8373,
  -43.8275,
  -43.8185,
  -43.8105,
  -43.8046,
  -43.8011,
  -43.8001,
  -43.8018,
  -43.8057,
  -43.812,
  -43.8193,
  -43.8269,
  -43.8334,
  -43.8378,
  -43.84,
  -43.8394,
  -43.8361,
  -43.8305,
  -43.8231,
  -43.8143,
  -43.8039,
  -43.7902,
  -43.7753,
  -43.7584,
  -43.7395,
  -43.7186,
  -43.6964,
  -43.6729,
  -43.6482,
  -43.6219,
  -43.593,
  -43.5608,
  -43.5245,
  -43.4834,
  -43.4371,
  -43.3865,
  -43.3323,
  -43.277,
  -43.2229,
  -43.1727,
  -43.1277,
  -43.0891,
  -43.0564,
  -43.0288,
  -43.0051,
  -42.9845,
  -42.9651,
  -42.9467,
  -42.9294,
  -42.9138,
  -42.9013,
  -42.8928,
  -42.8896,
  -42.893,
  -42.903,
  -42.9187,
  -42.9392,
  -42.9625,
  -42.9925,
  -43.0255,
  -43.0601,
  -43.0967,
  -43.135,
  -43.1729,
  -43.2115,
  -43.2542,
  -43.3026,
  -43.3567,
  -43.4149,
  -43.5023,
  -43.5939,
  -43.6922,
  -43.8029,
  -43.9279,
  -44.065,
  -44.2164,
  -44.3817,
  -44.5596,
  -44.7471,
  -44.9395,
  -45.1304,
  -45.3128,
  -45.4809,
  -45.6308,
  -45.7614,
  -45.8729,
  -45.9674,
  -46.0479,
  -46.118,
  -46.1806,
  -46.2379,
  -46.2899,
  -46.338,
  -37.7943,
  -37.8797,
  -37.9646,
  -38.0445,
  -38.1235,
  -38.1994,
  -38.273,
  -38.3411,
  -38.4089,
  -38.4692,
  -38.5313,
  -38.5961,
  -38.6644,
  -38.736,
  -38.8128,
  -38.8927,
  -38.9726,
  -39.0521,
  -39.1336,
  -39.2167,
  -39.3021,
  -39.3892,
  -39.4781,
  -39.5749,
  -39.6781,
  -39.7887,
  -39.9062,
  -40.0298,
  -40.1574,
  -40.2888,
  -40.423,
  -40.5596,
  -40.7016,
  -40.8452,
  -40.9927,
  -41.1391,
  -41.2842,
  -41.427,
  -41.5679,
  -41.7044,
  -41.8351,
  -41.9597,
  -42.0768,
  -42.1867,
  -42.2893,
  -42.3831,
  -42.4694,
  -42.5497,
  -42.6263,
  -42.7,
  -42.7749,
  -42.8498,
  -42.924,
  -42.9954,
  -43.0638,
  -43.1288,
  -43.1926,
  -43.2568,
  -43.3228,
  -43.392,
  -43.4652,
  -43.5437,
  -43.627,
  -43.715,
  -43.8069,
  -43.8998,
  -43.9949,
  -44.0911,
  -44.1886,
  -44.2879,
  -44.3897,
  -44.4934,
  -44.5986,
  -44.7054,
  -44.8127,
  -44.9208,
  -45.03,
  -45.1418,
  -45.2568,
  -45.375,
  -45.4958,
  -45.6176,
  -45.7379,
  -45.8564,
  -45.9698,
  -46.0759,
  -46.1725,
  -46.2575,
  -46.3295,
  -46.3883,
  -46.4347,
  -46.47,
  -46.4958,
  -46.5125,
  -46.5198,
  -46.5151,
  -46.4972,
  -46.4614,
  -46.4074,
  -46.3353,
  -46.2443,
  -46.1316,
  -46.0014,
  -45.8533,
  -45.6954,
  -45.5307,
  -45.364,
  -45.2019,
  -45.0543,
  -44.9143,
  -44.7881,
  -44.6776,
  -44.5955,
  -44.5304,
  -44.4807,
  -44.441,
  -44.4083,
  -44.3831,
  -44.3638,
  -44.3529,
  -44.3483,
  -44.3511,
  -44.3574,
  -44.3654,
  -44.3761,
  -44.3943,
  -44.4116,
  -44.4228,
  -44.4337,
  -44.4404,
  -44.4456,
  -44.4445,
  -44.4421,
  -44.443,
  -44.4411,
  -44.437,
  -44.4288,
  -44.4163,
  -44.3994,
  -44.3786,
  -44.3516,
  -44.3192,
  -44.2862,
  -44.2471,
  -44.2111,
  -44.1745,
  -44.1353,
  -44.0974,
  -44.0666,
  -44.0332,
  -43.9996,
  -43.9671,
  -43.9349,
  -43.9011,
  -43.8678,
  -43.8383,
  -43.8131,
  -43.7914,
  -43.7727,
  -43.7544,
  -43.7368,
  -43.7212,
  -43.7062,
  -43.6915,
  -43.6773,
  -43.6652,
  -43.6534,
  -43.64,
  -43.6259,
  -43.6092,
  -43.5913,
  -43.5723,
  -43.5532,
  -43.5323,
  -43.5159,
  -43.5038,
  -43.4956,
  -43.4924,
  -43.4964,
  -43.5027,
  -43.5145,
  -43.5272,
  -43.5384,
  -43.5476,
  -43.557,
  -43.5636,
  -43.5669,
  -43.5665,
  -43.5627,
  -43.5545,
  -43.546,
  -43.5376,
  -43.5308,
  -43.5279,
  -43.5283,
  -43.5317,
  -43.5379,
  -43.5458,
  -43.554,
  -43.5609,
  -43.5655,
  -43.5672,
  -43.566,
  -43.5625,
  -43.5572,
  -43.5514,
  -43.5452,
  -43.5397,
  -43.5346,
  -43.5303,
  -43.5266,
  -43.5241,
  -43.523,
  -43.5244,
  -43.5277,
  -43.5336,
  -43.5413,
  -43.5509,
  -43.561,
  -43.5725,
  -43.5831,
  -43.5917,
  -43.5979,
  -43.6017,
  -43.6025,
  -43.6009,
  -43.597,
  -43.5912,
  -43.5833,
  -43.5729,
  -43.5597,
  -43.5437,
  -43.5255,
  -43.5052,
  -43.4838,
  -43.4613,
  -43.4379,
  -43.4137,
  -43.3876,
  -43.3587,
  -43.3262,
  -43.289,
  -43.2466,
  -43.2002,
  -43.15,
  -43.0991,
  -43.0495,
  -43.0037,
  -42.9628,
  -42.929,
  -42.9008,
  -42.8773,
  -42.856,
  -42.8382,
  -42.8203,
  -42.8031,
  -42.7872,
  -42.773,
  -42.7622,
  -42.7552,
  -42.7539,
  -42.7595,
  -42.7724,
  -42.7909,
  -42.8132,
  -42.8394,
  -42.8715,
  -42.9077,
  -42.9396,
  -42.9838,
  -43.0277,
  -43.0708,
  -43.1129,
  -43.16,
  -43.2142,
  -43.2719,
  -43.3294,
  -43.4377,
  -43.5414,
  -43.6549,
  -43.7784,
  -43.914,
  -44.0632,
  -44.2249,
  -44.3985,
  -44.5814,
  -44.7692,
  -44.9571,
  -45.139,
  -45.3088,
  -45.4617,
  -45.5952,
  -45.7089,
  -45.8044,
  -45.8841,
  -45.9501,
  -46.0076,
  -46.0583,
  -46.1034,
  -46.1436,
  -46.1793,
  -37.7812,
  -37.8641,
  -37.9467,
  -38.0245,
  -38.1041,
  -38.178,
  -38.2469,
  -38.3129,
  -38.3728,
  -38.4307,
  -38.4898,
  -38.5513,
  -38.6157,
  -38.6841,
  -38.7564,
  -38.8332,
  -38.9093,
  -38.9857,
  -39.0703,
  -39.153,
  -39.2366,
  -39.3247,
  -39.4165,
  -39.511,
  -39.6139,
  -39.726,
  -39.8457,
  -39.9706,
  -40.0995,
  -40.2316,
  -40.365,
  -40.5001,
  -40.6403,
  -40.7837,
  -40.9333,
  -41.0796,
  -41.2266,
  -41.3708,
  -41.5115,
  -41.6494,
  -41.782,
  -41.9091,
  -42.0285,
  -42.1392,
  -42.2435,
  -42.3395,
  -42.4272,
  -42.5085,
  -42.5856,
  -42.6604,
  -42.7341,
  -42.807,
  -42.8779,
  -42.9455,
  -43.0097,
  -43.0708,
  -43.1307,
  -43.1916,
  -43.254,
  -43.3188,
  -43.3881,
  -43.4628,
  -43.5424,
  -43.6262,
  -43.7139,
  -43.8036,
  -43.8944,
  -43.9856,
  -44.0778,
  -44.1711,
  -44.2658,
  -44.3619,
  -44.4589,
  -44.5575,
  -44.657,
  -44.7574,
  -44.8578,
  -44.9612,
  -45.0676,
  -45.176,
  -45.2862,
  -45.3963,
  -45.5055,
  -45.6107,
  -45.7099,
  -45.8008,
  -45.8805,
  -45.9469,
  -45.9999,
  -46.0393,
  -46.0675,
  -46.0857,
  -46.0987,
  -46.1043,
  -46.1045,
  -46.0979,
  -46.0796,
  -46.0479,
  -45.9989,
  -45.9333,
  -45.8494,
  -45.7451,
  -45.6227,
  -45.4822,
  -45.332,
  -45.1737,
  -45.0129,
  -44.8555,
  -44.7118,
  -44.5733,
  -44.4448,
  -44.333,
  -44.2477,
  -44.1807,
  -44.1285,
  -44.0874,
  -44.053,
  -44.0254,
  -44.0015,
  -43.9844,
  -43.9731,
  -43.9673,
  -43.965,
  -43.962,
  -43.9645,
  -43.9729,
  -43.9842,
  -43.9947,
  -44.0045,
  -44.0114,
  -44.0188,
  -44.0186,
  -44.0161,
  -44.0177,
  -44.013,
  -44.0063,
  -43.9987,
  -43.9881,
  -43.9707,
  -43.9492,
  -43.9218,
  -43.8899,
  -43.8558,
  -43.8157,
  -43.779,
  -43.7421,
  -43.7046,
  -43.6681,
  -43.6353,
  -43.5988,
  -43.5609,
  -43.5249,
  -43.4924,
  -43.4582,
  -43.4265,
  -43.3981,
  -43.3745,
  -43.3547,
  -43.3384,
  -43.3219,
  -43.3069,
  -43.2956,
  -43.2844,
  -43.2752,
  -43.267,
  -43.2604,
  -43.2537,
  -43.2445,
  -43.234,
  -43.2209,
  -43.2058,
  -43.1894,
  -43.1735,
  -43.1556,
  -43.1427,
  -43.1327,
  -43.1277,
  -43.1261,
  -43.1302,
  -43.1363,
  -43.1453,
  -43.1555,
  -43.1636,
  -43.1687,
  -43.1757,
  -43.1813,
  -43.1857,
  -43.1898,
  -43.1917,
  -43.1888,
  -43.1846,
  -43.1804,
  -43.1783,
  -43.1799,
  -43.1843,
  -43.1929,
  -43.2043,
  -43.2165,
  -43.2288,
  -43.2403,
  -43.2491,
  -43.2547,
  -43.2572,
  -43.2569,
  -43.255,
  -43.2526,
  -43.251,
  -43.2501,
  -43.2488,
  -43.2497,
  -43.2513,
  -43.254,
  -43.2579,
  -43.2638,
  -43.2714,
  -43.281,
  -43.2922,
  -43.3054,
  -43.3195,
  -43.3336,
  -43.3472,
  -43.3592,
  -43.369,
  -43.3764,
  -43.381,
  -43.3828,
  -43.3823,
  -43.3798,
  -43.3749,
  -43.3665,
  -43.3547,
  -43.3398,
  -43.322,
  -43.3017,
  -43.2805,
  -43.2581,
  -43.2352,
  -43.2126,
  -43.1886,
  -43.1615,
  -43.1326,
  -43.0997,
  -43.0617,
  -43.0212,
  -42.9758,
  -42.9295,
  -42.8854,
  -42.8447,
  -42.8084,
  -42.7791,
  -42.7546,
  -42.7352,
  -42.7191,
  -42.7035,
  -42.684,
  -42.6667,
  -42.6536,
  -42.6441,
  -42.6366,
  -42.6317,
  -42.6319,
  -42.6386,
  -42.6529,
  -42.673,
  -42.697,
  -42.7267,
  -42.7577,
  -42.8036,
  -42.8439,
  -42.894,
  -42.9418,
  -42.9906,
  -43.038,
  -43.0917,
  -43.1543,
  -43.225,
  -43.3078,
  -43.4132,
  -43.5253,
  -43.6474,
  -43.7802,
  -43.9256,
  -44.082,
  -44.2495,
  -44.4254,
  -44.6068,
  -44.7884,
  -44.966,
  -45.134,
  -45.2877,
  -45.4231,
  -45.5395,
  -45.6371,
  -45.7185,
  -45.7857,
  -45.8422,
  -45.8904,
  -45.9324,
  -45.9688,
  -46.0003,
  -46.027,
  -37.7886,
  -37.8681,
  -37.9491,
  -38.0256,
  -38.0989,
  -38.1683,
  -38.2324,
  -38.2933,
  -38.3486,
  -38.4037,
  -38.4593,
  -38.5164,
  -38.5778,
  -38.6404,
  -38.7098,
  -38.7814,
  -38.8548,
  -38.9305,
  -39.0122,
  -39.0951,
  -39.1782,
  -39.2619,
  -39.3501,
  -39.4485,
  -39.553,
  -39.665,
  -39.789,
  -39.9178,
  -40.0497,
  -40.1822,
  -40.3183,
  -40.454,
  -40.5931,
  -40.7343,
  -40.8823,
  -41.0317,
  -41.1782,
  -41.3209,
  -41.4627,
  -41.5998,
  -41.7351,
  -41.8636,
  -41.9854,
  -42.0996,
  -42.2058,
  -42.3037,
  -42.393,
  -42.4759,
  -42.5542,
  -42.6294,
  -42.7027,
  -42.7737,
  -42.8418,
  -42.9059,
  -42.9649,
  -43.0221,
  -43.0785,
  -43.1355,
  -43.1943,
  -43.2559,
  -43.321,
  -43.391,
  -43.4658,
  -43.5454,
  -43.6284,
  -43.7137,
  -43.8001,
  -43.8866,
  -43.9732,
  -44.0601,
  -44.1468,
  -44.2351,
  -44.324,
  -44.4141,
  -44.5054,
  -44.5976,
  -44.6912,
  -44.7861,
  -44.8835,
  -44.9819,
  -45.081,
  -45.1797,
  -45.2763,
  -45.3687,
  -45.454,
  -45.53,
  -45.5939,
  -45.643,
  -45.6768,
  -45.6987,
  -45.709,
  -45.7127,
  -45.713,
  -45.7099,
  -45.7034,
  -45.6927,
  -45.6728,
  -45.6416,
  -45.5961,
  -45.5341,
  -45.4545,
  -45.3551,
  -45.2389,
  -45.1051,
  -44.9624,
  -44.8116,
  -44.6587,
  -44.5079,
  -44.371,
  -44.2391,
  -44.1158,
  -43.9983,
  -43.9104,
  -43.8422,
  -43.7901,
  -43.7464,
  -43.7096,
  -43.6772,
  -43.648,
  -43.6253,
  -43.6095,
  -43.5972,
  -43.5887,
  -43.5795,
  -43.5768,
  -43.578,
  -43.5807,
  -43.5864,
  -43.5933,
  -43.5978,
  -43.6025,
  -43.6041,
  -43.6019,
  -43.599,
  -43.5922,
  -43.583,
  -43.5744,
  -43.5654,
  -43.5484,
  -43.5263,
  -43.498,
  -43.4649,
  -43.4268,
  -43.3921,
  -43.3543,
  -43.3189,
  -43.2844,
  -43.2494,
  -43.2167,
  -43.1785,
  -43.1363,
  -43.0988,
  -43.0629,
  -43.0278,
  -42.9975,
  -42.9705,
  -42.9486,
  -42.9303,
  -42.9162,
  -42.9024,
  -42.8913,
  -42.8826,
  -42.878,
  -42.8744,
  -42.8718,
  -42.8683,
  -42.8651,
  -42.859,
  -42.8506,
  -42.8412,
  -42.8291,
  -42.8146,
  -42.8004,
  -42.789,
  -42.7791,
  -42.7717,
  -42.7679,
  -42.7693,
  -42.7739,
  -42.7782,
  -42.7867,
  -42.7939,
  -42.7987,
  -42.797,
  -42.8026,
  -42.8064,
  -42.8096,
  -42.8143,
  -42.8223,
  -42.8276,
  -42.8307,
  -42.8342,
  -42.8394,
  -42.8471,
  -42.8579,
  -42.8722,
  -42.8887,
  -42.9059,
  -42.9226,
  -42.9382,
  -42.9516,
  -42.9612,
  -42.9674,
  -42.9701,
  -42.9715,
  -42.9732,
  -42.9752,
  -42.9788,
  -42.9832,
  -42.9897,
  -42.9962,
  -43.0037,
  -43.0123,
  -43.0222,
  -43.0337,
  -43.0466,
  -43.0608,
  -43.0769,
  -43.0932,
  -43.1095,
  -43.1253,
  -43.1392,
  -43.1515,
  -43.1617,
  -43.17,
  -43.1755,
  -43.1784,
  -43.1792,
  -43.1758,
  -43.17,
  -43.16,
  -43.1461,
  -43.129,
  -43.1084,
  -43.0871,
  -43.0648,
  -43.0424,
  -43.0208,
  -42.9997,
  -42.977,
  -42.9526,
  -42.9246,
  -42.8928,
  -42.8585,
  -42.8191,
  -42.7787,
  -42.7399,
  -42.7045,
  -42.6713,
  -42.6459,
  -42.6254,
  -42.6099,
  -42.5967,
  -42.5825,
  -42.5623,
  -42.5357,
  -42.5275,
  -42.5296,
  -42.5258,
  -42.5232,
  -42.5224,
  -42.5258,
  -42.5351,
  -42.561,
  -42.5889,
  -42.6212,
  -42.6592,
  -42.718,
  -42.7725,
  -42.8245,
  -42.8802,
  -42.9333,
  -42.9876,
  -43.0492,
  -43.1213,
  -43.2077,
  -43.3056,
  -43.4161,
  -43.5375,
  -43.668,
  -43.8078,
  -43.9579,
  -44.1171,
  -44.2844,
  -44.4567,
  -44.6302,
  -44.8004,
  -44.9629,
  -45.1132,
  -45.2483,
  -45.3654,
  -45.4649,
  -45.5484,
  -45.6179,
  -45.6759,
  -45.7255,
  -45.7682,
  -45.805,
  -45.8364,
  -45.8621,
  -45.8826,
  -37.8194,
  -37.896,
  -37.9726,
  -38.046,
  -38.1145,
  -38.1774,
  -38.2363,
  -38.2902,
  -38.3389,
  -38.3887,
  -38.4392,
  -38.4914,
  -38.5478,
  -38.607,
  -38.6701,
  -38.7372,
  -38.8099,
  -38.8812,
  -38.958,
  -39.0405,
  -39.1226,
  -39.2065,
  -39.2959,
  -39.3938,
  -39.5,
  -39.6137,
  -39.7357,
  -39.8672,
  -40.0024,
  -40.1377,
  -40.2739,
  -40.4146,
  -40.5544,
  -40.6968,
  -40.8442,
  -40.9918,
  -41.1375,
  -41.2805,
  -41.422,
  -41.5607,
  -41.6963,
  -41.827,
  -41.9506,
  -42.0669,
  -42.1747,
  -42.2738,
  -42.3647,
  -42.4489,
  -42.5274,
  -42.6032,
  -42.6763,
  -42.7462,
  -42.8117,
  -42.8728,
  -42.9296,
  -42.9833,
  -43.0359,
  -43.089,
  -43.1438,
  -43.2013,
  -43.2619,
  -43.3267,
  -43.396,
  -43.4704,
  -43.5469,
  -43.6278,
  -43.7095,
  -43.7908,
  -43.8719,
  -43.9525,
  -44.033,
  -44.1136,
  -44.1942,
  -44.2759,
  -44.359,
  -44.4427,
  -44.528,
  -44.6143,
  -44.7018,
  -44.7904,
  -44.8787,
  -44.9661,
  -45.05,
  -45.1299,
  -45.202,
  -45.2636,
  -45.3127,
  -45.3467,
  -45.3655,
  -45.3712,
  -45.3685,
  -45.3596,
  -45.3485,
  -45.3369,
  -45.324,
  -45.3083,
  -45.2861,
  -45.2537,
  -45.2084,
  -45.1474,
  -45.0678,
  -44.971,
  -44.8589,
  -44.7299,
  -44.5946,
  -44.4529,
  -44.3093,
  -44.1697,
  -44.0433,
  -43.923,
  -43.8078,
  -43.6964,
  -43.5998,
  -43.5286,
  -43.4722,
  -43.4256,
  -43.3854,
  -43.3484,
  -43.3136,
  -43.2854,
  -43.2595,
  -43.2397,
  -43.2256,
  -43.2129,
  -43.2017,
  -43.1961,
  -43.1943,
  -43.1943,
  -43.1957,
  -43.1955,
  -43.1966,
  -43.1973,
  -43.1948,
  -43.1909,
  -43.1824,
  -43.1718,
  -43.1615,
  -43.1557,
  -43.1396,
  -43.115,
  -43.0835,
  -43.0459,
  -43.0114,
  -42.9748,
  -42.9396,
  -42.9063,
  -42.873,
  -42.84,
  -42.809,
  -42.7728,
  -42.7329,
  -42.6909,
  -42.6507,
  -42.6124,
  -42.5807,
  -42.5533,
  -42.531,
  -42.5154,
  -42.5034,
  -42.4914,
  -42.4818,
  -42.4792,
  -42.4802,
  -42.4828,
  -42.487,
  -42.489,
  -42.4888,
  -42.486,
  -42.4813,
  -42.4761,
  -42.4684,
  -42.4562,
  -42.4453,
  -42.4364,
  -42.4279,
  -42.4225,
  -42.421,
  -42.4214,
  -42.4273,
  -42.4316,
  -42.438,
  -42.4428,
  -42.4463,
  -42.4438,
  -42.4497,
  -42.4541,
  -42.4586,
  -42.4651,
  -42.4761,
  -42.4847,
  -42.4948,
  -42.506,
  -42.5189,
  -42.5337,
  -42.5504,
  -42.5706,
  -42.5925,
  -42.6148,
  -42.6362,
  -42.6569,
  -42.6739,
  -42.6874,
  -42.6969,
  -42.704,
  -42.7105,
  -42.7154,
  -42.7217,
  -42.729,
  -42.7383,
  -42.7484,
  -42.7599,
  -42.7719,
  -42.7849,
  -42.7983,
  -42.813,
  -42.8286,
  -42.8454,
  -42.862,
  -42.8798,
  -42.8975,
  -42.9143,
  -42.9296,
  -42.9438,
  -42.9564,
  -42.9679,
  -42.9768,
  -42.9837,
  -42.9879,
  -42.9892,
  -42.986,
  -42.9783,
  -42.9659,
  -42.9497,
  -42.929,
  -42.9073,
  -42.8844,
  -42.862,
  -42.8406,
  -42.8208,
  -42.801,
  -42.7807,
  -42.7577,
  -42.7315,
  -42.7046,
  -42.6711,
  -42.6368,
  -42.6043,
  -42.5761,
  -42.5484,
  -42.5288,
  -42.5122,
  -42.501,
  -42.4918,
  -42.481,
  -42.4662,
  -42.4508,
  -42.4403,
  -42.4371,
  -42.4338,
  -42.4317,
  -42.4283,
  -42.4181,
  -42.431,
  -42.4688,
  -42.499,
  -42.5457,
  -42.6073,
  -42.6684,
  -42.7264,
  -42.7843,
  -42.846,
  -42.9031,
  -42.9654,
  -43.0369,
  -43.1184,
  -43.2179,
  -43.3272,
  -43.4472,
  -43.5762,
  -43.7123,
  -43.8556,
  -44.0056,
  -44.1619,
  -44.3225,
  -44.485,
  -44.6451,
  -44.7988,
  -44.9425,
  -45.0733,
  -45.189,
  -45.2884,
  -45.3729,
  -45.4448,
  -45.5053,
  -45.5579,
  -45.6035,
  -45.6441,
  -45.6791,
  -45.7083,
  -45.7312,
  -45.7483,
  -37.8659,
  -37.9418,
  -38.0158,
  -38.0859,
  -38.1493,
  -38.2058,
  -38.2584,
  -38.3036,
  -38.346,
  -38.3887,
  -38.4339,
  -38.4798,
  -38.5287,
  -38.5825,
  -38.6402,
  -38.7026,
  -38.7683,
  -38.8373,
  -38.911,
  -38.99,
  -39.0725,
  -39.1576,
  -39.2472,
  -39.3464,
  -39.4544,
  -39.5686,
  -39.6932,
  -39.8234,
  -39.9586,
  -40.0925,
  -40.2295,
  -40.3703,
  -40.5195,
  -40.6671,
  -40.8123,
  -40.9598,
  -41.1042,
  -41.2483,
  -41.3911,
  -41.5309,
  -41.668,
  -41.7994,
  -41.9232,
  -42.0401,
  -42.1483,
  -42.2477,
  -42.3392,
  -42.424,
  -42.5044,
  -42.5809,
  -42.6536,
  -42.7224,
  -42.7863,
  -42.8454,
  -42.8994,
  -42.9501,
  -42.9994,
  -43.0488,
  -43.0996,
  -43.1518,
  -43.208,
  -43.2675,
  -43.3311,
  -43.399,
  -43.471,
  -43.5457,
  -43.6226,
  -43.698,
  -43.7731,
  -43.8477,
  -43.9213,
  -43.9946,
  -44.0678,
  -44.1412,
  -44.2158,
  -44.2909,
  -44.3662,
  -44.4436,
  -44.5215,
  -44.5997,
  -44.6776,
  -44.7543,
  -44.8282,
  -44.8962,
  -44.956,
  -45.0049,
  -45.0405,
  -45.0613,
  -45.068,
  -45.0619,
  -45.0473,
  -45.0288,
  -45.0097,
  -44.9913,
  -44.9722,
  -44.9521,
  -44.9264,
  -44.8916,
  -44.8445,
  -44.7822,
  -44.7028,
  -44.6065,
  -44.4951,
  -44.3703,
  -44.2389,
  -44.1062,
  -43.9724,
  -43.8446,
  -43.7295,
  -43.6194,
  -43.5147,
  -43.4115,
  -43.3186,
  -43.2382,
  -43.177,
  -43.1253,
  -43.0803,
  -43.0382,
  -42.9951,
  -42.9608,
  -42.93,
  -42.9035,
  -42.8835,
  -42.866,
  -42.8504,
  -42.8361,
  -42.826,
  -42.8168,
  -42.8117,
  -42.8028,
  -42.8014,
  -42.8002,
  -42.7962,
  -42.789,
  -42.7792,
  -42.7672,
  -42.7552,
  -42.7463,
  -42.7367,
  -42.7108,
  -42.6716,
  -42.6379,
  -42.6043,
  -42.5682,
  -42.5364,
  -42.5042,
  -42.4726,
  -42.4369,
  -42.4036,
  -42.3693,
  -42.337,
  -42.2914,
  -42.2519,
  -42.2132,
  -42.1816,
  -42.1525,
  -42.1315,
  -42.1124,
  -42.0965,
  -42.0902,
  -42.0898,
  -42.0896,
  -42.0926,
  -42.0985,
  -42.1094,
  -42.1165,
  -42.1177,
  -42.1194,
  -42.1195,
  -42.1206,
  -42.1192,
  -42.113,
  -42.1038,
  -42.0942,
  -42.0875,
  -42.084,
  -42.0844,
  -42.0842,
  -42.0888,
  -42.0938,
  -42.0994,
  -42.1044,
  -42.1085,
  -42.1073,
  -42.1151,
  -42.1196,
  -42.1268,
  -42.1361,
  -42.1525,
  -42.1651,
  -42.1785,
  -42.1961,
  -42.2144,
  -42.2355,
  -42.2591,
  -42.2857,
  -42.3144,
  -42.3427,
  -42.3696,
  -42.395,
  -42.4171,
  -42.4348,
  -42.4488,
  -42.4607,
  -42.4711,
  -42.4809,
  -42.4887,
  -42.4994,
  -42.5117,
  -42.5262,
  -42.5414,
  -42.557,
  -42.5733,
  -42.59,
  -42.6074,
  -42.6253,
  -42.6439,
  -42.6625,
  -42.6808,
  -42.6989,
  -42.7162,
  -42.7329,
  -42.7489,
  -42.7638,
  -42.7778,
  -42.7904,
  -42.8014,
  -42.8097,
  -42.8151,
  -42.8152,
  -42.8099,
  -42.7996,
  -42.7848,
  -42.7645,
  -42.743,
  -42.7198,
  -42.6971,
  -42.6764,
  -42.6559,
  -42.6391,
  -42.6229,
  -42.6056,
  -42.5857,
  -42.5667,
  -42.5396,
  -42.5109,
  -42.485,
  -42.4633,
  -42.4412,
  -42.4271,
  -42.4177,
  -42.4116,
  -42.4058,
  -42.4009,
  -42.3921,
  -42.3817,
  -42.3724,
  -42.3663,
  -42.364,
  -42.3624,
  -42.3515,
  -42.3448,
  -42.3855,
  -42.4342,
  -42.475,
  -42.5228,
  -42.5834,
  -42.6476,
  -42.7139,
  -42.7751,
  -42.8364,
  -42.901,
  -42.9728,
  -43.0555,
  -43.1506,
  -43.2579,
  -43.3765,
  -43.5031,
  -43.6372,
  -43.7753,
  -43.9172,
  -44.0623,
  -44.2099,
  -44.3585,
  -44.5054,
  -44.6475,
  -44.7812,
  -44.904,
  -45.0145,
  -45.1121,
  -45.1961,
  -45.269,
  -45.3329,
  -45.3896,
  -45.4396,
  -45.4848,
  -45.5254,
  -45.5613,
  -45.5902,
  -45.6125,
  -45.628,
  -37.9226,
  -37.996,
  -38.0672,
  -38.1345,
  -38.1952,
  -38.2482,
  -38.2957,
  -38.3344,
  -38.3688,
  -38.4056,
  -38.4427,
  -38.481,
  -38.5236,
  -38.5707,
  -38.6226,
  -38.6783,
  -38.7382,
  -38.8021,
  -38.8701,
  -38.945,
  -39.0243,
  -39.1097,
  -39.2011,
  -39.3033,
  -39.4142,
  -39.5346,
  -39.6634,
  -39.7941,
  -39.9276,
  -40.0611,
  -40.197,
  -40.3362,
  -40.4855,
  -40.6401,
  -40.7878,
  -40.9354,
  -41.0819,
  -41.2262,
  -41.37,
  -41.5114,
  -41.6489,
  -41.78,
  -41.9044,
  -42.0205,
  -42.1276,
  -42.2258,
  -42.3169,
  -42.402,
  -42.4823,
  -42.5588,
  -42.6309,
  -42.6986,
  -42.7611,
  -42.8173,
  -42.8695,
  -42.9173,
  -42.9639,
  -43.0099,
  -43.0571,
  -43.1063,
  -43.158,
  -43.2126,
  -43.2704,
  -43.3323,
  -43.3978,
  -43.4662,
  -43.5364,
  -43.6064,
  -43.6751,
  -43.7438,
  -43.8101,
  -43.8764,
  -43.9423,
  -44.0079,
  -44.0737,
  -44.1399,
  -44.2072,
  -44.2752,
  -44.3435,
  -44.4115,
  -44.4792,
  -44.5457,
  -44.6089,
  -44.6659,
  -44.7148,
  -44.7528,
  -44.7774,
  -44.787,
  -44.7841,
  -44.77,
  -44.7475,
  -44.7222,
  -44.6978,
  -44.6745,
  -44.6522,
  -44.6284,
  -44.5996,
  -44.5614,
  -44.5117,
  -44.4471,
  -44.366,
  -44.2686,
  -44.157,
  -44.0334,
  -43.9068,
  -43.779,
  -43.6544,
  -43.5368,
  -43.4303,
  -43.3301,
  -43.2365,
  -43.1463,
  -43.0618,
  -42.9854,
  -42.9188,
  -42.8608,
  -42.8038,
  -42.7527,
  -42.7035,
  -42.6617,
  -42.6221,
  -42.5873,
  -42.5613,
  -42.5413,
  -42.5177,
  -42.4935,
  -42.4724,
  -42.4549,
  -42.4418,
  -42.4292,
  -42.4224,
  -42.4174,
  -42.4084,
  -42.398,
  -42.3896,
  -42.3777,
  -42.3663,
  -42.3495,
  -42.3371,
  -42.32,
  -42.2795,
  -42.2464,
  -42.2139,
  -42.1773,
  -42.1458,
  -42.1145,
  -42.0813,
  -42.0448,
  -42.0118,
  -41.9762,
  -41.9509,
  -41.9045,
  -41.8659,
  -41.8302,
  -41.8004,
  -41.7756,
  -41.7533,
  -41.729,
  -41.7134,
  -41.7049,
  -41.7021,
  -41.7065,
  -41.7148,
  -41.7246,
  -41.7386,
  -41.7513,
  -41.7562,
  -41.7626,
  -41.7685,
  -41.7761,
  -41.7819,
  -41.7811,
  -41.7733,
  -41.7673,
  -41.7614,
  -41.7592,
  -41.7589,
  -41.7589,
  -41.7629,
  -41.7687,
  -41.7763,
  -41.7841,
  -41.7921,
  -41.7926,
  -41.8007,
  -41.8093,
  -41.8197,
  -41.8311,
  -41.8506,
  -41.8661,
  -41.8828,
  -41.9022,
  -41.9242,
  -41.9499,
  -41.9795,
  -42.0128,
  -42.0484,
  -42.0828,
  -42.1174,
  -42.1502,
  -42.1783,
  -42.2018,
  -42.2202,
  -42.2381,
  -42.2552,
  -42.2701,
  -42.2816,
  -42.2949,
  -42.3097,
  -42.3257,
  -42.3434,
  -42.3621,
  -42.3811,
  -42.4004,
  -42.4202,
  -42.4396,
  -42.4586,
  -42.4771,
  -42.4956,
  -42.5137,
  -42.5317,
  -42.549,
  -42.5664,
  -42.5838,
  -42.6011,
  -42.6177,
  -42.6316,
  -42.6443,
  -42.6545,
  -42.6584,
  -42.6565,
  -42.6486,
  -42.6355,
  -42.6167,
  -42.5963,
  -42.5744,
  -42.5527,
  -42.5331,
  -42.5149,
  -42.5016,
  -42.4889,
  -42.475,
  -42.4604,
  -42.4482,
  -42.4294,
  -42.4057,
  -42.3858,
  -42.37,
  -42.3532,
  -42.3437,
  -42.339,
  -42.3366,
  -42.335,
  -42.334,
  -42.3285,
  -42.3206,
  -42.3144,
  -42.3108,
  -42.3095,
  -42.3111,
  -42.301,
  -42.3211,
  -42.3722,
  -42.4174,
  -42.4654,
  -42.5207,
  -42.584,
  -42.6506,
  -42.7173,
  -42.7844,
  -42.8536,
  -42.9278,
  -43.0104,
  -43.1042,
  -43.2088,
  -43.325,
  -43.4503,
  -43.5822,
  -43.7177,
  -43.8543,
  -43.9907,
  -44.1264,
  -44.2605,
  -44.392,
  -44.5188,
  -44.639,
  -44.7504,
  -44.8519,
  -44.943,
  -45.025,
  -45.0979,
  -45.1633,
  -45.2228,
  -45.278,
  -45.329,
  -45.3759,
  -45.4188,
  -45.4558,
  -45.4858,
  -45.5079,
  -45.5222,
  -37.9843,
  -38.0562,
  -38.1239,
  -38.1888,
  -38.247,
  -38.2967,
  -38.3398,
  -38.3759,
  -38.4081,
  -38.4393,
  -38.468,
  -38.4962,
  -38.5298,
  -38.5689,
  -38.6129,
  -38.661,
  -38.7136,
  -38.7713,
  -38.8328,
  -38.9018,
  -38.9774,
  -39.0611,
  -39.1548,
  -39.2645,
  -39.3848,
  -39.5104,
  -39.6408,
  -39.7728,
  -39.9054,
  -40.0392,
  -40.1751,
  -40.313,
  -40.4595,
  -40.6186,
  -40.7705,
  -40.9188,
  -41.068,
  -41.2161,
  -41.3613,
  -41.5032,
  -41.64,
  -41.7696,
  -41.8921,
  -42.0057,
  -42.1099,
  -42.206,
  -42.2955,
  -42.3789,
  -42.4587,
  -42.5346,
  -42.6059,
  -42.6723,
  -42.7333,
  -42.789,
  -42.8394,
  -42.8855,
  -42.9293,
  -42.9723,
  -43.016,
  -43.0612,
  -43.1083,
  -43.1576,
  -43.2098,
  -43.2654,
  -43.3235,
  -43.3852,
  -43.4482,
  -43.5116,
  -43.5747,
  -43.6375,
  -43.6987,
  -43.7589,
  -43.818,
  -43.8763,
  -43.9338,
  -43.9914,
  -44.0493,
  -44.1082,
  -44.1667,
  -44.2249,
  -44.2825,
  -44.3377,
  -44.3907,
  -44.4377,
  -44.4773,
  -44.5056,
  -44.5211,
  -44.5237,
  -44.515,
  -44.4955,
  -44.4689,
  -44.4361,
  -44.4123,
  -44.3867,
  -44.3618,
  -44.3361,
  -44.3046,
  -44.2643,
  -44.2121,
  -44.1438,
  -44.0597,
  -43.9613,
  -43.8481,
  -43.7232,
  -43.5976,
  -43.4736,
  -43.3568,
  -43.2473,
  -43.1484,
  -43.0544,
  -42.9681,
  -42.8848,
  -42.8053,
  -42.7332,
  -42.6675,
  -42.6068,
  -42.5505,
  -42.4958,
  -42.4422,
  -42.3946,
  -42.3469,
  -42.3025,
  -42.2667,
  -42.2301,
  -42.199,
  -42.1733,
  -42.1425,
  -42.116,
  -42.0954,
  -42.0756,
  -42.0582,
  -42.051,
  -42.0349,
  -42.0255,
  -42.0172,
  -42.0075,
  -41.9967,
  -41.9773,
  -41.9594,
  -41.9492,
  -41.9066,
  -41.8714,
  -41.8373,
  -41.8008,
  -41.7682,
  -41.7372,
  -41.7036,
  -41.6695,
  -41.6361,
  -41.6016,
  -41.5784,
  -41.5461,
  -41.5003,
  -41.4669,
  -41.4401,
  -41.4182,
  -41.3967,
  -41.3699,
  -41.3499,
  -41.3466,
  -41.3376,
  -41.3437,
  -41.3543,
  -41.3666,
  -41.3817,
  -41.3992,
  -41.4097,
  -41.4194,
  -41.4276,
  -41.4411,
  -41.4538,
  -41.4602,
  -41.4591,
  -41.4552,
  -41.4522,
  -41.4513,
  -41.4512,
  -41.4518,
  -41.4532,
  -41.4601,
  -41.4701,
  -41.4835,
  -41.4936,
  -41.4966,
  -41.5069,
  -41.518,
  -41.5285,
  -41.5389,
  -41.5597,
  -41.5774,
  -41.5974,
  -41.6199,
  -41.6457,
  -41.6744,
  -41.7094,
  -41.752,
  -41.7932,
  -41.8362,
  -41.8777,
  -41.919,
  -41.9552,
  -41.9858,
  -42.0107,
  -42.0366,
  -42.0615,
  -42.0813,
  -42.0975,
  -42.1126,
  -42.1291,
  -42.1466,
  -42.1651,
  -42.1855,
  -42.2065,
  -42.2281,
  -42.2496,
  -42.2696,
  -42.2877,
  -42.3058,
  -42.3231,
  -42.3418,
  -42.3609,
  -42.3795,
  -42.3983,
  -42.4184,
  -42.4391,
  -42.4598,
  -42.4794,
  -42.4969,
  -42.5121,
  -42.5204,
  -42.5221,
  -42.5169,
  -42.5062,
  -42.4898,
  -42.4722,
  -42.4534,
  -42.434,
  -42.4172,
  -42.4011,
  -42.3904,
  -42.3802,
  -42.3671,
  -42.3543,
  -42.3496,
  -42.337,
  -42.323,
  -42.3088,
  -42.2959,
  -42.2831,
  -42.2762,
  -42.2754,
  -42.2763,
  -42.2769,
  -42.278,
  -42.2739,
  -42.2666,
  -42.2658,
  -42.2684,
  -42.2714,
  -42.2853,
  -42.3014,
  -42.3338,
  -42.3756,
  -42.423,
  -42.4783,
  -42.5391,
  -42.6054,
  -42.6746,
  -42.7479,
  -42.8225,
  -42.9022,
  -42.987,
  -43.0799,
  -43.1834,
  -43.296,
  -43.418,
  -43.5465,
  -43.6787,
  -43.812,
  -43.943,
  -44.0702,
  -44.1929,
  -44.3104,
  -44.4216,
  -44.5256,
  -44.6216,
  -44.7101,
  -44.7905,
  -44.8643,
  -44.9338,
  -44.9995,
  -45.0613,
  -45.1209,
  -45.1778,
  -45.2314,
  -45.2812,
  -45.3258,
  -45.3639,
  -45.394,
  -45.4154,
  -45.428,
  -38.0488,
  -38.1184,
  -38.1859,
  -38.2489,
  -38.3046,
  -38.3524,
  -38.3922,
  -38.4252,
  -38.4532,
  -38.4791,
  -38.5018,
  -38.5193,
  -38.5409,
  -38.5698,
  -38.6074,
  -38.6482,
  -38.696,
  -38.7468,
  -38.8022,
  -38.8668,
  -38.9389,
  -39.0215,
  -39.1182,
  -39.2339,
  -39.3595,
  -39.4902,
  -39.6239,
  -39.7563,
  -39.8889,
  -40.0222,
  -40.1603,
  -40.2986,
  -40.4465,
  -40.6048,
  -40.7607,
  -40.9123,
  -41.0642,
  -41.215,
  -41.362,
  -41.5022,
  -41.6375,
  -41.7655,
  -41.8833,
  -41.9928,
  -42.0936,
  -42.187,
  -42.2745,
  -42.3575,
  -42.4359,
  -42.5106,
  -42.5804,
  -42.6449,
  -42.7042,
  -42.758,
  -42.8062,
  -42.8501,
  -42.8911,
  -42.9309,
  -42.9701,
  -43.0116,
  -43.0543,
  -43.0989,
  -43.1461,
  -43.1961,
  -43.2486,
  -43.3033,
  -43.3595,
  -43.4164,
  -43.4739,
  -43.5309,
  -43.5869,
  -43.6412,
  -43.6939,
  -43.7452,
  -43.7947,
  -43.8426,
  -43.8915,
  -43.9409,
  -43.9898,
  -44.0382,
  -44.0855,
  -44.1315,
  -44.1743,
  -44.212,
  -44.2426,
  -44.2628,
  -44.2716,
  -44.2685,
  -44.2555,
  -44.2329,
  -44.2042,
  -44.1745,
  -44.1457,
  -44.1185,
  -44.0918,
  -44.0652,
  -44.0317,
  -43.9904,
  -43.9384,
  -43.8696,
  -43.7839,
  -43.6842,
  -43.571,
  -43.4453,
  -43.3163,
  -43.1919,
  -43.0801,
  -42.9744,
  -42.8786,
  -42.7876,
  -42.7029,
  -42.6225,
  -42.5411,
  -42.4744,
  -42.4058,
  -42.3489,
  -42.2927,
  -42.24,
  -42.1832,
  -42.128,
  -42.0792,
  -42.0326,
  -41.9871,
  -41.9423,
  -41.8998,
  -41.8698,
  -41.8359,
  -41.8012,
  -41.7673,
  -41.7414,
  -41.7215,
  -41.7083,
  -41.687,
  -41.6782,
  -41.6699,
  -41.6575,
  -41.6454,
  -41.6268,
  -41.6074,
  -41.6008,
  -41.5601,
  -41.5192,
  -41.4835,
  -41.4456,
  -41.4128,
  -41.3802,
  -41.3454,
  -41.31,
  -41.2791,
  -41.2463,
  -41.2195,
  -41.2021,
  -41.1607,
  -41.1306,
  -41.1053,
  -41.0825,
  -41.0615,
  -41.0313,
  -41.0108,
  -41.0051,
  -40.9993,
  -41.0027,
  -41.0107,
  -41.0219,
  -41.04,
  -41.063,
  -41.0768,
  -41.0883,
  -41.0999,
  -41.1181,
  -41.1346,
  -41.1472,
  -41.1543,
  -41.1592,
  -41.1589,
  -41.1547,
  -41.1553,
  -41.1567,
  -41.1575,
  -41.1659,
  -41.1783,
  -41.1892,
  -41.2,
  -41.2053,
  -41.2177,
  -41.2328,
  -41.2462,
  -41.2568,
  -41.2806,
  -41.3011,
  -41.3256,
  -41.3515,
  -41.3793,
  -41.4149,
  -41.4604,
  -41.504,
  -41.5529,
  -41.6021,
  -41.6491,
  -41.6977,
  -41.7424,
  -41.7814,
  -41.8146,
  -41.8526,
  -41.8844,
  -41.9084,
  -41.9286,
  -41.9485,
  -41.9679,
  -41.9875,
  -42.0079,
  -42.029,
  -42.0504,
  -42.073,
  -42.0955,
  -42.1168,
  -42.1362,
  -42.1538,
  -42.1699,
  -42.188,
  -42.2074,
  -42.2278,
  -42.2484,
  -42.2714,
  -42.295,
  -42.3194,
  -42.3436,
  -42.3674,
  -42.3885,
  -42.4009,
  -42.4062,
  -42.4042,
  -42.3965,
  -42.3827,
  -42.3682,
  -42.3527,
  -42.3376,
  -42.3222,
  -42.304,
  -42.2923,
  -42.2802,
  -42.2585,
  -42.2493,
  -42.2514,
  -42.2543,
  -42.2463,
  -42.2408,
  -42.2357,
  -42.2295,
  -42.2292,
  -42.2323,
  -42.2358,
  -42.2363,
  -42.2402,
  -42.2374,
  -42.2344,
  -42.237,
  -42.2485,
  -42.2635,
  -42.2867,
  -42.3156,
  -42.3517,
  -42.3979,
  -42.4473,
  -42.5075,
  -42.5744,
  -42.647,
  -42.7245,
  -42.8076,
  -42.8922,
  -42.9805,
  -43.076,
  -43.1777,
  -43.2878,
  -43.4056,
  -43.5288,
  -43.6573,
  -43.7869,
  -43.9143,
  -44.0365,
  -44.1517,
  -44.2587,
  -44.3567,
  -44.4457,
  -44.5257,
  -44.5981,
  -44.6646,
  -44.7266,
  -44.7873,
  -44.8484,
  -44.9111,
  -44.9739,
  -45.0365,
  -45.0965,
  -45.1534,
  -45.2051,
  -45.2504,
  -45.2874,
  -45.3154,
  -45.3341,
  -45.3436,
  -38.1202,
  -38.1884,
  -38.2542,
  -38.3152,
  -38.3684,
  -38.4134,
  -38.4492,
  -38.4787,
  -38.5029,
  -38.5226,
  -38.539,
  -38.5534,
  -38.566,
  -38.5833,
  -38.6076,
  -38.6399,
  -38.6796,
  -38.7256,
  -38.7769,
  -38.8387,
  -38.9078,
  -38.9892,
  -39.0872,
  -39.2036,
  -39.3359,
  -39.4721,
  -39.6113,
  -39.7494,
  -39.884,
  -40.0188,
  -40.1538,
  -40.2945,
  -40.4442,
  -40.6039,
  -40.7608,
  -40.9162,
  -41.0709,
  -41.2221,
  -41.3682,
  -41.5076,
  -41.64,
  -41.7643,
  -41.8793,
  -41.9845,
  -42.0813,
  -42.1715,
  -42.2565,
  -42.3373,
  -42.4142,
  -42.4868,
  -42.5545,
  -42.6167,
  -42.6724,
  -42.7235,
  -42.769,
  -42.81,
  -42.8479,
  -42.8841,
  -42.9205,
  -42.9575,
  -42.9959,
  -43.0359,
  -43.0783,
  -43.1229,
  -43.1694,
  -43.2178,
  -43.2673,
  -43.3183,
  -43.3702,
  -43.4212,
  -43.4719,
  -43.5212,
  -43.5681,
  -43.6119,
  -43.6536,
  -43.6941,
  -43.7342,
  -43.7743,
  -43.8135,
  -43.8522,
  -43.8893,
  -43.9253,
  -43.9584,
  -43.9871,
  -44.0093,
  -44.0229,
  -44.026,
  -44.0186,
  -44.0021,
  -43.979,
  -43.9509,
  -43.9197,
  -43.8906,
  -43.8642,
  -43.8374,
  -43.8101,
  -43.7776,
  -43.7371,
  -43.6854,
  -43.6165,
  -43.5324,
  -43.4309,
  -43.3184,
  -43.1943,
  -43.0649,
  -42.9354,
  -42.82,
  -42.7137,
  -42.6156,
  -42.5237,
  -42.4393,
  -42.3627,
  -42.2824,
  -42.218,
  -42.1562,
  -42.0954,
  -42.0393,
  -41.9865,
  -41.93,
  -41.8785,
  -41.8259,
  -41.7625,
  -41.7065,
  -41.6565,
  -41.6127,
  -41.5737,
  -41.5307,
  -41.4935,
  -41.457,
  -41.4288,
  -41.4068,
  -41.3872,
  -41.3632,
  -41.3527,
  -41.3402,
  -41.3275,
  -41.3151,
  -41.2924,
  -41.2709,
  -41.2564,
  -41.2348,
  -41.186,
  -41.1505,
  -41.1117,
  -41.0737,
  -41.0383,
  -41.0034,
  -40.9675,
  -40.9369,
  -40.9045,
  -40.8779,
  -40.8662,
  -40.8421,
  -40.8069,
  -40.7848,
  -40.7624,
  -40.7372,
  -40.7103,
  -40.6919,
  -40.6837,
  -40.6835,
  -40.6804,
  -40.6916,
  -40.7001,
  -40.7141,
  -40.7406,
  -40.7561,
  -40.7704,
  -40.7833,
  -40.8011,
  -40.822,
  -40.8417,
  -40.8561,
  -40.8678,
  -40.8722,
  -40.8739,
  -40.8788,
  -40.8817,
  -40.8842,
  -40.9013,
  -40.9133,
  -40.921,
  -40.9285,
  -40.9377,
  -40.9482,
  -40.9706,
  -40.9867,
  -40.9966,
  -41.0217,
  -41.0437,
  -41.0685,
  -41.0949,
  -41.1236,
  -41.1563,
  -41.2192,
  -41.2716,
  -41.3297,
  -41.3854,
  -41.4384,
  -41.4939,
  -41.55,
  -41.5958,
  -41.6421,
  -41.6889,
  -41.7271,
  -41.7571,
  -41.7816,
  -41.8059,
  -41.8283,
  -41.8506,
  -41.8726,
  -41.8945,
  -41.9168,
  -41.9393,
  -41.9629,
  -41.9856,
  -42.006,
  -42.0236,
  -42.0403,
  -42.0576,
  -42.0765,
  -42.0976,
  -42.1199,
  -42.1451,
  -42.1717,
  -42.1991,
  -42.2282,
  -42.2569,
  -42.2843,
  -42.3011,
  -42.3104,
  -42.3126,
  -42.3087,
  -42.2994,
  -42.2899,
  -42.2797,
  -42.2703,
  -42.2614,
  -42.2384,
  -42.2264,
  -42.22,
  -42.2015,
  -42.1876,
  -42.1912,
  -42.1948,
  -42.1886,
  -42.1852,
  -42.1885,
  -42.1937,
  -42.1982,
  -42.2022,
  -42.2059,
  -42.2042,
  -42.2037,
  -42.1932,
  -42.1907,
  -42.1995,
  -42.2295,
  -42.2596,
  -42.2909,
  -42.3309,
  -42.3768,
  -42.4306,
  -42.4868,
  -42.5525,
  -42.6296,
  -42.7118,
  -42.8013,
  -42.8949,
  -42.9896,
  -43.0867,
  -43.188,
  -43.2952,
  -43.4088,
  -43.5279,
  -43.6515,
  -43.7766,
  -43.901,
  -44.0203,
  -44.1318,
  -44.233,
  -44.3229,
  -44.4006,
  -44.4669,
  -44.5242,
  -44.5744,
  -44.6211,
  -44.6692,
  -44.7203,
  -44.7772,
  -44.8397,
  -44.9056,
  -44.9719,
  -45.0365,
  -45.0936,
  -45.1447,
  -45.1877,
  -45.2209,
  -45.2441,
  -45.2576,
  -45.2619,
  -38.1985,
  -38.2637,
  -38.3272,
  -38.3853,
  -38.4354,
  -38.4773,
  -38.5106,
  -38.5362,
  -38.5559,
  -38.5708,
  -38.5813,
  -38.5903,
  -38.5964,
  -38.6013,
  -38.6167,
  -38.6407,
  -38.6702,
  -38.7093,
  -38.7559,
  -38.8172,
  -38.8871,
  -38.9713,
  -39.0715,
  -39.1885,
  -39.3228,
  -39.4618,
  -39.6049,
  -39.7469,
  -39.8869,
  -40.0237,
  -40.1621,
  -40.3069,
  -40.4578,
  -40.6134,
  -40.7712,
  -40.9311,
  -41.0873,
  -41.2401,
  -41.3838,
  -41.5212,
  -41.6493,
  -41.769,
  -41.8793,
  -41.9804,
  -42.0735,
  -42.1603,
  -42.2425,
  -42.32,
  -42.3947,
  -42.4647,
  -42.5294,
  -42.5885,
  -42.642,
  -42.6895,
  -42.7314,
  -42.7684,
  -42.8024,
  -42.8341,
  -42.8656,
  -42.8981,
  -42.9315,
  -42.9664,
  -43.0036,
  -43.0414,
  -43.0824,
  -43.125,
  -43.1685,
  -43.2143,
  -43.2612,
  -43.3086,
  -43.3554,
  -43.3989,
  -43.4403,
  -43.4779,
  -43.512,
  -43.5443,
  -43.5757,
  -43.6067,
  -43.6365,
  -43.6656,
  -43.6917,
  -43.7186,
  -43.7423,
  -43.7626,
  -43.7776,
  -43.7849,
  -43.7836,
  -43.7738,
  -43.7559,
  -43.7316,
  -43.7032,
  -43.6737,
  -43.644,
  -43.6168,
  -43.5905,
  -43.5631,
  -43.5314,
  -43.4916,
  -43.4413,
  -43.3745,
  -43.2919,
  -43.1941,
  -43.0837,
  -42.9633,
  -42.838,
  -42.7132,
  -42.5882,
  -42.4711,
  -42.366,
  -42.2699,
  -42.1858,
  -42.1122,
  -42.0388,
  -41.9736,
  -41.9077,
  -41.8444,
  -41.7844,
  -41.732,
  -41.674,
  -41.6244,
  -41.5746,
  -41.5203,
  -41.4597,
  -41.3972,
  -41.3424,
  -41.2946,
  -41.2466,
  -41.2032,
  -41.1678,
  -41.136,
  -41.1127,
  -41.0902,
  -41.0683,
  -41.0529,
  -41.0375,
  -41.021,
  -41.0014,
  -40.981,
  -40.9608,
  -40.9417,
  -40.9314,
  -40.8777,
  -40.8326,
  -40.7935,
  -40.7505,
  -40.7115,
  -40.6748,
  -40.6404,
  -40.6111,
  -40.5814,
  -40.5565,
  -40.5464,
  -40.5324,
  -40.4953,
  -40.4743,
  -40.4498,
  -40.4196,
  -40.3984,
  -40.3819,
  -40.3738,
  -40.3741,
  -40.3753,
  -40.3736,
  -40.3869,
  -40.404,
  -40.4309,
  -40.4558,
  -40.4739,
  -40.4861,
  -40.5014,
  -40.5224,
  -40.5485,
  -40.5713,
  -40.5858,
  -40.6009,
  -40.6062,
  -40.6158,
  -40.6241,
  -40.6289,
  -40.6523,
  -40.6666,
  -40.6777,
  -40.678,
  -40.6895,
  -40.7022,
  -40.7262,
  -40.7432,
  -40.7553,
  -40.774,
  -40.7935,
  -40.8141,
  -40.8311,
  -40.8583,
  -40.8997,
  -40.9732,
  -41.0505,
  -41.1192,
  -41.1813,
  -41.2393,
  -41.3092,
  -41.3801,
  -41.4402,
  -41.4939,
  -41.5464,
  -41.5905,
  -41.6272,
  -41.6572,
  -41.6838,
  -41.7096,
  -41.7339,
  -41.758,
  -41.7808,
  -41.803,
  -41.8263,
  -41.8503,
  -41.8743,
  -41.8958,
  -41.9148,
  -41.9309,
  -41.949,
  -41.966,
  -41.9868,
  -42.0093,
  -42.0374,
  -42.0681,
  -42.101,
  -42.1347,
  -42.168,
  -42.2019,
  -42.2232,
  -42.2361,
  -42.2422,
  -42.2431,
  -42.2394,
  -42.2365,
  -42.2326,
  -42.2299,
  -42.2267,
  -42.2149,
  -42.2128,
  -42.2093,
  -42.2027,
  -42.1967,
  -42.2023,
  -42.1982,
  -42.1828,
  -42.1731,
  -42.1743,
  -42.1726,
  -42.1826,
  -42.1885,
  -42.1908,
  -42.1885,
  -42.1787,
  -42.1729,
  -42.1778,
  -42.1918,
  -42.2218,
  -42.2693,
  -42.3124,
  -42.3593,
  -42.4171,
  -42.4813,
  -42.5477,
  -42.6271,
  -42.7133,
  -42.8052,
  -42.9048,
  -43.0073,
  -43.1087,
  -43.2113,
  -43.3163,
  -43.4247,
  -43.5385,
  -43.6555,
  -43.7747,
  -43.8945,
  -44.0111,
  -44.1209,
  -44.221,
  -44.308,
  -44.3801,
  -44.4391,
  -44.4852,
  -44.5217,
  -44.553,
  -44.5846,
  -44.6223,
  -44.6679,
  -44.7227,
  -44.7878,
  -44.8577,
  -44.9261,
  -44.9915,
  -45.0484,
  -45.0951,
  -45.132,
  -45.1576,
  -45.1731,
  -45.179,
  -45.1769,
  -38.2815,
  -38.3449,
  -38.4047,
  -38.459,
  -38.5052,
  -38.5433,
  -38.5724,
  -38.5937,
  -38.6089,
  -38.6186,
  -38.6233,
  -38.6247,
  -38.6235,
  -38.6235,
  -38.6322,
  -38.6479,
  -38.6699,
  -38.7037,
  -38.7479,
  -38.8061,
  -38.8766,
  -38.9631,
  -39.0672,
  -39.1878,
  -39.3223,
  -39.4639,
  -39.6075,
  -39.752,
  -39.8953,
  -40.0369,
  -40.1801,
  -40.3273,
  -40.4806,
  -40.6396,
  -40.801,
  -40.9598,
  -41.1177,
  -41.2672,
  -41.4078,
  -41.541,
  -41.6646,
  -41.7786,
  -41.8847,
  -41.982,
  -42.0716,
  -42.1552,
  -42.2344,
  -42.3103,
  -42.3821,
  -42.4493,
  -42.5106,
  -42.5658,
  -42.615,
  -42.6578,
  -42.695,
  -42.7272,
  -42.7561,
  -42.7813,
  -42.8067,
  -42.8329,
  -42.8602,
  -42.8892,
  -42.9202,
  -42.9531,
  -42.9884,
  -43.0256,
  -43.0646,
  -43.1054,
  -43.149,
  -43.1924,
  -43.2344,
  -43.2735,
  -43.3089,
  -43.3404,
  -43.3669,
  -43.3917,
  -43.4149,
  -43.4371,
  -43.458,
  -43.4778,
  -43.4967,
  -43.5146,
  -43.53,
  -43.5427,
  -43.5507,
  -43.5524,
  -43.547,
  -43.5346,
  -43.5153,
  -43.4901,
  -43.4613,
  -43.4309,
  -43.4,
  -43.3716,
  -43.3442,
  -43.3162,
  -43.2852,
  -43.247,
  -43.1996,
  -43.1376,
  -43.0592,
  -42.9656,
  -42.8602,
  -42.744,
  -42.6249,
  -42.5019,
  -42.3804,
  -42.261,
  -42.1462,
  -42.0423,
  -41.9614,
  -41.8861,
  -41.8081,
  -41.7373,
  -41.662,
  -41.5942,
  -41.5331,
  -41.4806,
  -41.4273,
  -41.3761,
  -41.3243,
  -41.2724,
  -41.2166,
  -41.1561,
  -41.0926,
  -41.0384,
  -40.9873,
  -40.9365,
  -40.8946,
  -40.8611,
  -40.8363,
  -40.8094,
  -40.7857,
  -40.7735,
  -40.7561,
  -40.7365,
  -40.7177,
  -40.7019,
  -40.6846,
  -40.668,
  -40.648,
  -40.606,
  -40.5523,
  -40.5071,
  -40.4631,
  -40.4185,
  -40.3715,
  -40.3352,
  -40.3055,
  -40.2809,
  -40.261,
  -40.2436,
  -40.2251,
  -40.2039,
  -40.1817,
  -40.1457,
  -40.1145,
  -40.0905,
  -40.0758,
  -40.0657,
  -40.0637,
  -40.0646,
  -40.0674,
  -40.0814,
  -40.1034,
  -40.131,
  -40.1635,
  -40.19,
  -40.2041,
  -40.2164,
  -40.2466,
  -40.2754,
  -40.3027,
  -40.3182,
  -40.3425,
  -40.3578,
  -40.3692,
  -40.3838,
  -40.4039,
  -40.4246,
  -40.4363,
  -40.4496,
  -40.4634,
  -40.4651,
  -40.48,
  -40.5048,
  -40.5263,
  -40.529,
  -40.5298,
  -40.5559,
  -40.5693,
  -40.582,
  -40.6044,
  -40.6644,
  -40.7629,
  -40.851,
  -40.9297,
  -41.0041,
  -41.0793,
  -41.1639,
  -41.2405,
  -41.3073,
  -41.3646,
  -41.4224,
  -41.4725,
  -41.5163,
  -41.5514,
  -41.5821,
  -41.6103,
  -41.6382,
  -41.6629,
  -41.6862,
  -41.7094,
  -41.734,
  -41.7596,
  -41.7852,
  -41.8079,
  -41.8282,
  -41.845,
  -41.8636,
  -41.8819,
  -41.8997,
  -41.9208,
  -41.9504,
  -41.9824,
  -42.0256,
  -42.0642,
  -42.103,
  -42.1397,
  -42.1642,
  -42.1807,
  -42.1911,
  -42.1975,
  -42.2002,
  -42.2038,
  -42.2068,
  -42.2113,
  -42.2156,
  -42.211,
  -42.2146,
  -42.2172,
  -42.2174,
  -42.2134,
  -42.2189,
  -42.2125,
  -42.2012,
  -42.1885,
  -42.1884,
  -42.1874,
  -42.1889,
  -42.1938,
  -42.197,
  -42.1976,
  -42.1995,
  -42.203,
  -42.2146,
  -42.2327,
  -42.2569,
  -42.2978,
  -42.3477,
  -42.4047,
  -42.4721,
  -42.5486,
  -42.6262,
  -42.718,
  -42.8179,
  -42.922,
  -43.0274,
  -43.1359,
  -43.2412,
  -43.3455,
  -43.4497,
  -43.5556,
  -43.6641,
  -43.776,
  -43.8887,
  -44.0004,
  -44.1079,
  -44.2075,
  -44.2957,
  -44.3693,
  -44.4262,
  -44.4685,
  -44.4974,
  -44.5181,
  -44.5361,
  -44.5582,
  -44.5895,
  -44.6332,
  -44.6901,
  -44.7569,
  -44.8282,
  -44.8974,
  -44.9594,
  -45.0116,
  -45.051,
  -45.0784,
  -45.094,
  -45.0992,
  -45.0961,
  -45.0866,
  -38.3691,
  -38.4283,
  -38.4838,
  -38.5332,
  -38.5746,
  -38.6071,
  -38.6304,
  -38.6473,
  -38.6576,
  -38.6622,
  -38.6623,
  -38.6582,
  -38.6519,
  -38.6472,
  -38.6485,
  -38.6576,
  -38.6747,
  -38.7037,
  -38.7461,
  -38.8046,
  -38.8787,
  -38.967,
  -39.0739,
  -39.199,
  -39.334,
  -39.4766,
  -39.623,
  -39.7705,
  -39.9166,
  -40.0622,
  -40.2096,
  -40.3594,
  -40.5155,
  -40.6775,
  -40.8399,
  -41.0004,
  -41.1545,
  -41.3014,
  -41.4394,
  -41.5678,
  -41.6872,
  -41.7977,
  -41.8997,
  -41.9933,
  -42.0798,
  -42.1605,
  -42.237,
  -42.3103,
  -42.3792,
  -42.4428,
  -42.5004,
  -42.5512,
  -42.5944,
  -42.6317,
  -42.663,
  -42.6889,
  -42.7105,
  -42.7295,
  -42.7477,
  -42.7665,
  -42.7862,
  -42.8073,
  -42.8308,
  -42.8567,
  -42.8858,
  -42.9173,
  -42.9515,
  -42.9891,
  -43.027,
  -43.0663,
  -43.1043,
  -43.1399,
  -43.1708,
  -43.1972,
  -43.2196,
  -43.2388,
  -43.2556,
  -43.2709,
  -43.2844,
  -43.2964,
  -43.3074,
  -43.3173,
  -43.3249,
  -43.3304,
  -43.3316,
  -43.3279,
  -43.3171,
  -43.302,
  -43.2806,
  -43.2538,
  -43.2238,
  -43.1923,
  -43.1607,
  -43.1302,
  -43.1009,
  -43.0714,
  -43.0399,
  -43.0033,
  -42.9584,
  -42.8994,
  -42.8264,
  -42.7387,
  -42.6393,
  -42.5292,
  -42.4167,
  -42.2997,
  -42.1829,
  -42.0662,
  -41.9621,
  -41.8644,
  -41.7775,
  -41.6928,
  -41.6033,
  -41.5239,
  -41.4433,
  -41.364,
  -41.3011,
  -41.2473,
  -41.1902,
  -41.1342,
  -41.0814,
  -41.0285,
  -40.9727,
  -40.9217,
  -40.8649,
  -40.806,
  -40.7432,
  -40.694,
  -40.6433,
  -40.6014,
  -40.576,
  -40.5504,
  -40.5247,
  -40.5145,
  -40.4918,
  -40.4756,
  -40.4628,
  -40.4601,
  -40.4507,
  -40.4145,
  -40.3719,
  -40.3352,
  -40.2761,
  -40.2217,
  -40.1668,
  -40.1259,
  -40.0875,
  -40.0506,
  -40.0243,
  -40.004,
  -39.9781,
  -39.9559,
  -39.9426,
  -39.918,
  -39.8953,
  -39.86,
  -39.8281,
  -39.7927,
  -39.7719,
  -39.7575,
  -39.7534,
  -39.7529,
  -39.7625,
  -39.7731,
  -39.806,
  -39.8487,
  -39.8865,
  -39.9197,
  -39.9359,
  -39.9461,
  -39.9641,
  -40.0036,
  -40.0458,
  -40.0728,
  -40.0998,
  -40.1266,
  -40.1572,
  -40.1841,
  -40.2041,
  -40.2157,
  -40.2285,
  -40.2378,
  -40.2583,
  -40.2695,
  -40.2919,
  -40.3212,
  -40.3327,
  -40.3341,
  -40.3384,
  -40.3476,
  -40.3672,
  -40.3824,
  -40.4251,
  -40.4991,
  -40.5942,
  -40.6684,
  -40.7605,
  -40.8632,
  -40.9629,
  -41.0503,
  -41.1243,
  -41.1923,
  -41.2539,
  -41.3183,
  -41.3741,
  -41.4223,
  -41.4631,
  -41.498,
  -41.5303,
  -41.5589,
  -41.5851,
  -41.6098,
  -41.6352,
  -41.6607,
  -41.6873,
  -41.7144,
  -41.74,
  -41.762,
  -41.7803,
  -41.7999,
  -41.8195,
  -41.8431,
  -41.8681,
  -41.8985,
  -41.9289,
  -41.9714,
  -42.0149,
  -42.0554,
  -42.0936,
  -42.1206,
  -42.1411,
  -42.1564,
  -42.1686,
  -42.1779,
  -42.1888,
  -42.2003,
  -42.2124,
  -42.2244,
  -42.2263,
  -42.2358,
  -42.2434,
  -42.2477,
  -42.2483,
  -42.2539,
  -42.2473,
  -42.2365,
  -42.2274,
  -42.2215,
  -42.2179,
  -42.2181,
  -42.2197,
  -42.2229,
  -42.2262,
  -42.2338,
  -42.2414,
  -42.2557,
  -42.2776,
  -42.3088,
  -42.3473,
  -42.3998,
  -42.4657,
  -42.5437,
  -42.6315,
  -42.7227,
  -42.8274,
  -42.9373,
  -43.0492,
  -43.1599,
  -43.2706,
  -43.3758,
  -43.4777,
  -43.5775,
  -43.6775,
  -43.7797,
  -43.8833,
  -43.9873,
  -44.0894,
  -44.1866,
  -44.2751,
  -44.3515,
  -44.4128,
  -44.4574,
  -44.4869,
  -44.5047,
  -44.5157,
  -44.527,
  -44.5451,
  -44.575,
  -44.6181,
  -44.6754,
  -44.7412,
  -44.8103,
  -44.8752,
  -44.9309,
  -44.9741,
  -45.0034,
  -45.0193,
  -45.0235,
  -45.0182,
  -45.006,
  -44.9887,
  -38.4571,
  -38.5104,
  -38.5603,
  -38.6036,
  -38.6384,
  -38.6651,
  -38.6838,
  -38.6955,
  -38.7013,
  -38.7011,
  -38.6964,
  -38.6882,
  -38.6778,
  -38.6701,
  -38.6641,
  -38.6667,
  -38.6796,
  -38.7084,
  -38.7528,
  -38.8101,
  -38.8865,
  -38.9803,
  -39.0911,
  -39.217,
  -39.3531,
  -39.4977,
  -39.647,
  -39.7977,
  -39.9486,
  -40.0988,
  -40.249,
  -40.4027,
  -40.562,
  -40.7259,
  -40.8893,
  -41.0489,
  -41.2021,
  -41.3464,
  -41.4809,
  -41.6059,
  -41.7211,
  -41.8275,
  -41.9257,
  -42.0162,
  -42.1,
  -42.1784,
  -42.2517,
  -42.3225,
  -42.3884,
  -42.4484,
  -42.5016,
  -42.5472,
  -42.5856,
  -42.6162,
  -42.6402,
  -42.6578,
  -42.6707,
  -42.6811,
  -42.6906,
  -42.7,
  -42.7103,
  -42.7223,
  -42.7371,
  -42.7543,
  -42.7765,
  -42.8026,
  -42.8329,
  -42.8663,
  -42.9019,
  -42.9374,
  -42.9714,
  -43.003,
  -43.0304,
  -43.0534,
  -43.072,
  -43.0869,
  -43.0991,
  -43.109,
  -43.1165,
  -43.1222,
  -43.1256,
  -43.1286,
  -43.1293,
  -43.1278,
  -43.1231,
  -43.1142,
  -43.1004,
  -43.0813,
  -43.0574,
  -43.0284,
  -42.9961,
  -42.9621,
  -42.9273,
  -42.8927,
  -42.859,
  -42.8261,
  -42.7926,
  -42.7561,
  -42.7134,
  -42.6585,
  -42.5906,
  -42.5099,
  -42.4176,
  -42.3122,
  -42.2072,
  -42.1006,
  -41.9919,
  -41.8844,
  -41.7849,
  -41.6854,
  -41.5927,
  -41.5027,
  -41.4151,
  -41.3347,
  -41.2529,
  -41.1696,
  -41.1029,
  -41.0403,
  -40.9714,
  -40.9116,
  -40.8537,
  -40.8004,
  -40.7455,
  -40.6947,
  -40.6407,
  -40.5812,
  -40.5131,
  -40.4612,
  -40.4136,
  -40.3637,
  -40.3344,
  -40.3026,
  -40.278,
  -40.2609,
  -40.2445,
  -40.2335,
  -40.2298,
  -40.2322,
  -40.2181,
  -40.1657,
  -40.1121,
  -40.0772,
  -40.0098,
  -39.9446,
  -39.891,
  -39.8405,
  -39.8048,
  -39.7765,
  -39.7566,
  -39.739,
  -39.7226,
  -39.6932,
  -39.6771,
  -39.6335,
  -39.6015,
  -39.5766,
  -39.5463,
  -39.5224,
  -39.5045,
  -39.478,
  -39.4677,
  -39.4646,
  -39.4752,
  -39.4957,
  -39.5237,
  -39.5575,
  -39.5966,
  -39.6474,
  -39.6811,
  -39.6855,
  -39.7064,
  -39.7493,
  -39.7942,
  -39.8237,
  -39.8578,
  -39.9001,
  -39.9458,
  -39.99,
  -40.0237,
  -40.0513,
  -40.071,
  -40.0871,
  -40.096,
  -40.1145,
  -40.1394,
  -40.1726,
  -40.187,
  -40.1839,
  -40.1823,
  -40.1823,
  -40.2007,
  -40.2401,
  -40.307,
  -40.3765,
  -40.447,
  -40.5491,
  -40.6632,
  -40.7749,
  -40.8718,
  -40.9465,
  -41.0195,
  -41.0999,
  -41.1697,
  -41.2356,
  -41.2936,
  -41.345,
  -41.3909,
  -41.4307,
  -41.4663,
  -41.4972,
  -41.525,
  -41.5516,
  -41.5776,
  -41.6029,
  -41.6318,
  -41.6605,
  -41.6878,
  -41.7123,
  -41.7334,
  -41.7554,
  -41.7783,
  -41.8031,
  -41.8302,
  -41.8612,
  -41.8975,
  -41.94,
  -41.9829,
  -42.024,
  -42.0615,
  -42.0917,
  -42.1169,
  -42.1381,
  -42.1571,
  -42.1744,
  -42.1929,
  -42.2128,
  -42.2335,
  -42.2535,
  -42.265,
  -42.2798,
  -42.2913,
  -42.2985,
  -42.3,
  -42.3022,
  -42.2941,
  -42.283,
  -42.2727,
  -42.2657,
  -42.2617,
  -42.2603,
  -42.2603,
  -42.2618,
  -42.2645,
  -42.2731,
  -42.2832,
  -42.3001,
  -42.3251,
  -42.36,
  -42.4042,
  -42.4648,
  -42.5401,
  -42.6274,
  -42.7282,
  -42.8327,
  -42.9484,
  -43.0667,
  -43.1834,
  -43.2956,
  -43.4041,
  -43.5048,
  -43.6001,
  -43.6919,
  -43.7828,
  -43.8753,
  -43.9687,
  -44.0625,
  -44.1541,
  -44.2401,
  -44.3182,
  -44.3845,
  -44.4357,
  -44.4714,
  -44.4934,
  -44.5054,
  -44.5133,
  -44.5236,
  -44.5433,
  -44.5751,
  -44.6187,
  -44.6742,
  -44.7367,
  -44.7987,
  -44.8543,
  -44.8991,
  -44.9302,
  -44.9469,
  -44.9504,
  -44.9431,
  -44.928,
  -44.9075,
  -44.8835,
  -38.5417,
  -38.5905,
  -38.634,
  -38.6701,
  -38.6978,
  -38.7174,
  -38.7304,
  -38.7364,
  -38.7367,
  -38.7319,
  -38.7219,
  -38.7099,
  -38.6965,
  -38.6853,
  -38.6763,
  -38.6768,
  -38.6882,
  -38.7163,
  -38.76,
  -38.8202,
  -38.9001,
  -38.996,
  -39.1099,
  -39.2371,
  -39.3747,
  -39.5196,
  -39.6711,
  -39.8254,
  -39.9803,
  -40.1351,
  -40.2911,
  -40.4499,
  -40.6128,
  -40.7772,
  -40.941,
  -41.1005,
  -41.2529,
  -41.3966,
  -41.5299,
  -41.653,
  -41.7659,
  -41.8683,
  -41.9637,
  -42.0516,
  -42.1332,
  -42.21,
  -42.2822,
  -42.3509,
  -42.4137,
  -42.4699,
  -42.518,
  -42.5579,
  -42.5898,
  -42.6129,
  -42.6282,
  -42.6361,
  -42.6391,
  -42.6381,
  -42.6366,
  -42.6349,
  -42.634,
  -42.6352,
  -42.6396,
  -42.6486,
  -42.6633,
  -42.683,
  -42.7085,
  -42.7376,
  -42.7697,
  -42.8016,
  -42.8332,
  -42.8617,
  -42.8871,
  -42.9085,
  -42.9244,
  -42.9374,
  -42.9472,
  -42.9538,
  -42.9571,
  -42.9583,
  -42.958,
  -42.955,
  -42.9501,
  -42.9427,
  -42.9322,
  -42.9184,
  -42.9001,
  -42.8781,
  -42.8507,
  -42.8185,
  -42.7827,
  -42.7447,
  -42.704,
  -42.664,
  -42.6253,
  -42.588,
  -42.5515,
  -42.5132,
  -42.472,
  -42.4209,
  -42.3584,
  -42.2836,
  -42.1976,
  -42.0989,
  -42.0012,
  -41.9013,
  -41.8008,
  -41.7003,
  -41.6014,
  -41.5013,
  -41.4023,
  -41.309,
  -41.222,
  -41.1409,
  -41.0541,
  -40.9712,
  -40.8959,
  -40.8177,
  -40.7394,
  -40.6816,
  -40.6319,
  -40.5778,
  -40.5312,
  -40.4827,
  -40.4322,
  -40.3716,
  -40.3139,
  -40.25,
  -40.1977,
  -40.1444,
  -40.1035,
  -40.0698,
  -40.0403,
  -40.0192,
  -40.0081,
  -40.0148,
  -40.0299,
  -40.036,
  -40.0156,
  -39.9695,
  -39.9075,
  -39.8614,
  -39.7699,
  -39.6918,
  -39.6377,
  -39.5838,
  -39.5466,
  -39.5156,
  -39.4919,
  -39.4919,
  -39.4772,
  -39.4438,
  -39.4321,
  -39.3929,
  -39.3474,
  -39.309,
  -39.2753,
  -39.2647,
  -39.2387,
  -39.2283,
  -39.2119,
  -39.2075,
  -39.2221,
  -39.2386,
  -39.265,
  -39.301,
  -39.3455,
  -39.3993,
  -39.4323,
  -39.4446,
  -39.4782,
  -39.525,
  -39.5699,
  -39.601,
  -39.6439,
  -39.6974,
  -39.7506,
  -39.8064,
  -39.8529,
  -39.8929,
  -39.9265,
  -39.9529,
  -39.9765,
  -40.0035,
  -40.0253,
  -40.0415,
  -40.0531,
  -40.0588,
  -40.0695,
  -40.0784,
  -40.1004,
  -40.1527,
  -40.2351,
  -40.3038,
  -40.3641,
  -40.464,
  -40.5972,
  -40.7106,
  -40.794,
  -40.8647,
  -40.942,
  -41.0269,
  -41.0995,
  -41.1649,
  -41.2247,
  -41.28,
  -41.3295,
  -41.3737,
  -41.4125,
  -41.4449,
  -41.4745,
  -41.5019,
  -41.5287,
  -41.5574,
  -41.5879,
  -41.6187,
  -41.6483,
  -41.6753,
  -41.698,
  -41.7233,
  -41.7494,
  -41.7775,
  -41.8065,
  -41.8405,
  -41.8777,
  -41.9184,
  -41.9616,
  -42.0017,
  -42.0417,
  -42.0758,
  -42.1065,
  -42.1341,
  -42.1601,
  -42.1852,
  -42.2117,
  -42.2397,
  -42.269,
  -42.2962,
  -42.3153,
  -42.3354,
  -42.3511,
  -42.3608,
  -42.3635,
  -42.3662,
  -42.3599,
  -42.35,
  -42.341,
  -42.3339,
  -42.3302,
  -42.3274,
  -42.3258,
  -42.326,
  -42.3278,
  -42.3363,
  -42.3477,
  -42.3666,
  -42.3954,
  -42.4352,
  -42.4854,
  -42.5535,
  -42.6373,
  -42.7345,
  -42.8428,
  -42.9572,
  -43.0786,
  -43.2,
  -43.3167,
  -43.4256,
  -43.5275,
  -43.6196,
  -43.7049,
  -43.7857,
  -43.8641,
  -43.9444,
  -44.0262,
  -44.1087,
  -44.189,
  -44.265,
  -44.3331,
  -44.3907,
  -44.4352,
  -44.4665,
  -44.4862,
  -44.4986,
  -44.509,
  -44.5235,
  -44.5479,
  -44.5832,
  -44.6274,
  -44.6803,
  -44.7359,
  -44.7881,
  -44.8316,
  -44.8627,
  -44.8794,
  -44.8818,
  -44.873,
  -44.8555,
  -44.8319,
  -44.8049,
  -44.7763,
  -38.6215,
  -38.664,
  -38.7004,
  -38.7293,
  -38.7492,
  -38.7608,
  -38.7666,
  -38.7666,
  -38.7617,
  -38.7524,
  -38.7398,
  -38.7252,
  -38.7104,
  -38.696,
  -38.6864,
  -38.6871,
  -38.6966,
  -38.7255,
  -38.7686,
  -38.8309,
  -38.9119,
  -39.0094,
  -39.124,
  -39.2521,
  -39.3897,
  -39.5356,
  -39.6879,
  -39.8447,
  -40.0043,
  -40.1649,
  -40.3271,
  -40.4914,
  -40.6579,
  -40.825,
  -40.99,
  -41.15,
  -41.3037,
  -41.4483,
  -41.5825,
  -41.7065,
  -41.8191,
  -41.9218,
  -42.0156,
  -42.1019,
  -42.1822,
  -42.2576,
  -42.3287,
  -42.3951,
  -42.4548,
  -42.5066,
  -42.5495,
  -42.5821,
  -42.6064,
  -42.621,
  -42.6265,
  -42.6245,
  -42.6163,
  -42.6045,
  -42.5903,
  -42.5758,
  -42.5622,
  -42.5508,
  -42.5436,
  -42.5426,
  -42.5484,
  -42.5615,
  -42.581,
  -42.6057,
  -42.6333,
  -42.6626,
  -42.6917,
  -42.7189,
  -42.7438,
  -42.765,
  -42.7822,
  -42.7949,
  -42.8042,
  -42.8096,
  -42.8108,
  -42.8093,
  -42.8053,
  -42.7981,
  -42.7886,
  -42.7769,
  -42.762,
  -42.7427,
  -42.7203,
  -42.6936,
  -42.6622,
  -42.6263,
  -42.5861,
  -42.5426,
  -42.4966,
  -42.45,
  -42.4042,
  -42.3608,
  -42.3195,
  -42.2784,
  -42.2364,
  -42.187,
  -42.1286,
  -42.0592,
  -41.9797,
  -41.8874,
  -41.7953,
  -41.7018,
  -41.6072,
  -41.5122,
  -41.4181,
  -41.3171,
  -41.218,
  -41.1237,
  -41.0359,
  -40.953,
  -40.8557,
  -40.7732,
  -40.6909,
  -40.6119,
  -40.5295,
  -40.4672,
  -40.4141,
  -40.3615,
  -40.3089,
  -40.263,
  -40.2268,
  -40.1796,
  -40.128,
  -40.0705,
  -40.0122,
  -39.9447,
  -39.8942,
  -39.8527,
  -39.8249,
  -39.8038,
  -39.7899,
  -39.8029,
  -39.8296,
  -39.8328,
  -39.8105,
  -39.7784,
  -39.7276,
  -39.6721,
  -39.5772,
  -39.478,
  -39.4165,
  -39.3584,
  -39.3204,
  -39.2847,
  -39.2611,
  -39.2557,
  -39.2503,
  -39.2205,
  -39.2029,
  -39.1853,
  -39.1384,
  -39.0876,
  -39.058,
  -39.0429,
  -39.0129,
  -38.9939,
  -38.9794,
  -38.9859,
  -38.9998,
  -39.018,
  -39.0455,
  -39.0833,
  -39.1319,
  -39.1915,
  -39.2258,
  -39.2353,
  -39.2721,
  -39.3228,
  -39.3753,
  -39.4197,
  -39.4774,
  -39.5403,
  -39.6045,
  -39.6614,
  -39.7147,
  -39.7566,
  -39.7891,
  -39.8214,
  -39.8531,
  -39.8956,
  -39.9323,
  -39.9599,
  -39.9796,
  -39.9898,
  -40.0169,
  -40.0494,
  -40.0782,
  -40.1272,
  -40.2199,
  -40.2995,
  -40.3548,
  -40.4584,
  -40.5633,
  -40.6615,
  -40.7408,
  -40.8132,
  -40.8847,
  -40.9705,
  -41.0406,
  -41.1067,
  -41.1684,
  -41.2265,
  -41.2811,
  -41.328,
  -41.369,
  -41.4028,
  -41.4329,
  -41.4611,
  -41.4902,
  -41.5215,
  -41.5543,
  -41.5872,
  -41.6187,
  -41.6478,
  -41.6727,
  -41.6998,
  -41.7273,
  -41.7572,
  -41.7895,
  -41.8244,
  -41.8629,
  -41.904,
  -41.9463,
  -41.9884,
  -42.0315,
  -42.0713,
  -42.109,
  -42.144,
  -42.1783,
  -42.2129,
  -42.2495,
  -42.2868,
  -42.3239,
  -42.358,
  -42.3836,
  -42.4094,
  -42.4296,
  -42.4421,
  -42.4472,
  -42.4511,
  -42.4468,
  -42.4393,
  -42.4316,
  -42.4251,
  -42.4209,
  -42.4165,
  -42.4137,
  -42.4121,
  -42.4131,
  -42.421,
  -42.4329,
  -42.4541,
  -42.4863,
  -42.5315,
  -42.5874,
  -42.6624,
  -42.7525,
  -42.8563,
  -42.9705,
  -43.0883,
  -43.2108,
  -43.3298,
  -43.4412,
  -43.5417,
  -43.6332,
  -43.7133,
  -43.7858,
  -43.8534,
  -43.9194,
  -43.9867,
  -44.0554,
  -44.1258,
  -44.1962,
  -44.263,
  -44.3235,
  -44.375,
  -44.4158,
  -44.446,
  -44.4683,
  -44.4865,
  -44.5041,
  -44.5265,
  -44.5573,
  -44.5964,
  -44.6416,
  -44.6894,
  -44.7356,
  -44.7747,
  -44.8031,
  -44.8182,
  -44.8197,
  -44.8088,
  -44.7885,
  -44.7618,
  -44.7321,
  -44.7011,
  -44.67,
  -38.6917,
  -38.7276,
  -38.7568,
  -38.778,
  -38.791,
  -38.7964,
  -38.7957,
  -38.7896,
  -38.7789,
  -38.7656,
  -38.7496,
  -38.733,
  -38.7162,
  -38.7018,
  -38.692,
  -38.6907,
  -38.7028,
  -38.7317,
  -38.7766,
  -38.8386,
  -38.9197,
  -39.0183,
  -39.132,
  -39.2589,
  -39.3949,
  -39.5392,
  -39.6903,
  -39.8484,
  -40.0116,
  -40.1784,
  -40.3462,
  -40.5169,
  -40.6888,
  -40.861,
  -41.0301,
  -41.1954,
  -41.353,
  -41.5008,
  -41.6388,
  -41.7661,
  -41.8806,
  -41.9844,
  -42.0787,
  -42.1649,
  -42.2449,
  -42.3199,
  -42.3887,
  -42.4526,
  -42.5093,
  -42.5566,
  -42.594,
  -42.6209,
  -42.637,
  -42.6425,
  -42.6377,
  -42.6246,
  -42.6043,
  -42.5794,
  -42.5515,
  -42.5229,
  -42.495,
  -42.4701,
  -42.4494,
  -42.437,
  -42.4335,
  -42.439,
  -42.4524,
  -42.4724,
  -42.4979,
  -42.5246,
  -42.552,
  -42.5794,
  -42.6053,
  -42.6275,
  -42.646,
  -42.66,
  -42.6699,
  -42.6754,
  -42.6764,
  -42.6732,
  -42.6675,
  -42.6575,
  -42.6453,
  -42.6307,
  -42.6128,
  -42.5912,
  -42.5651,
  -42.5341,
  -42.498,
  -42.4569,
  -42.4107,
  -42.3605,
  -42.3071,
  -42.2532,
  -42.1993,
  -42.1488,
  -42.1013,
  -42.0559,
  -42.0123,
  -41.9632,
  -41.9066,
  -41.841,
  -41.7672,
  -41.6809,
  -41.5949,
  -41.5078,
  -41.4193,
  -41.3303,
  -41.2406,
  -41.1448,
  -41.0471,
  -40.9529,
  -40.8624,
  -40.7815,
  -40.6837,
  -40.5967,
  -40.5097,
  -40.4239,
  -40.342,
  -40.2724,
  -40.2156,
  -40.1579,
  -40.1054,
  -40.0728,
  -40.0393,
  -39.986,
  -39.9307,
  -39.8839,
  -39.8294,
  -39.78,
  -39.7204,
  -39.668,
  -39.6384,
  -39.6098,
  -39.5822,
  -39.5913,
  -39.6206,
  -39.6297,
  -39.6047,
  -39.5764,
  -39.5358,
  -39.4855,
  -39.4217,
  -39.3287,
  -39.2497,
  -39.1887,
  -39.1332,
  -39.0925,
  -39.0712,
  -39.0654,
  -39.0485,
  -39.0105,
  -39.0088,
  -38.9885,
  -38.9279,
  -38.8914,
  -38.8757,
  -38.8636,
  -38.8419,
  -38.8207,
  -38.7959,
  -38.7957,
  -38.81,
  -38.8428,
  -38.8756,
  -38.9149,
  -38.9651,
  -39.0206,
  -39.0458,
  -39.0601,
  -39.0936,
  -39.1454,
  -39.1941,
  -39.2432,
  -39.3036,
  -39.3747,
  -39.4579,
  -39.5261,
  -39.5821,
  -39.6285,
  -39.6638,
  -39.6939,
  -39.7294,
  -39.7852,
  -39.8366,
  -39.8837,
  -39.9184,
  -39.9551,
  -39.9921,
  -40.035,
  -40.0751,
  -40.1223,
  -40.2064,
  -40.3041,
  -40.3827,
  -40.4632,
  -40.5517,
  -40.6357,
  -40.7127,
  -40.7812,
  -40.8577,
  -40.9302,
  -40.9971,
  -41.0623,
  -41.1256,
  -41.187,
  -41.2439,
  -41.2921,
  -41.3334,
  -41.3677,
  -41.3984,
  -41.4277,
  -41.4575,
  -41.4922,
  -41.5277,
  -41.5628,
  -41.5963,
  -41.6275,
  -41.6537,
  -41.6818,
  -41.7104,
  -41.7411,
  -41.7751,
  -41.813,
  -41.8536,
  -41.8967,
  -41.9415,
  -41.9878,
  -42.0366,
  -42.0831,
  -42.1285,
  -42.1726,
  -42.2167,
  -42.2618,
  -42.3086,
  -42.3553,
  -42.4009,
  -42.4427,
  -42.4754,
  -42.5063,
  -42.5302,
  -42.5455,
  -42.5545,
  -42.56,
  -42.5584,
  -42.5519,
  -42.546,
  -42.5402,
  -42.5361,
  -42.5313,
  -42.527,
  -42.5239,
  -42.5238,
  -42.5306,
  -42.5428,
  -42.5651,
  -42.6007,
  -42.6502,
  -42.7128,
  -42.7927,
  -42.8873,
  -42.994,
  -43.1088,
  -43.2248,
  -43.3422,
  -43.4531,
  -43.5542,
  -43.6424,
  -43.7192,
  -43.7846,
  -43.842,
  -43.8945,
  -43.9457,
  -43.9994,
  -44.0558,
  -44.115,
  -44.176,
  -44.2355,
  -44.2911,
  -44.3404,
  -44.3817,
  -44.4147,
  -44.4434,
  -44.4704,
  -44.4978,
  -44.5294,
  -44.5657,
  -44.6081,
  -44.6524,
  -44.6944,
  -44.7303,
  -44.7565,
  -44.7694,
  -44.7693,
  -44.7553,
  -44.7314,
  -44.7,
  -44.6662,
  -44.6322,
  -44.5995,
  -44.5685,
  -38.7518,
  -38.7814,
  -38.8041,
  -38.8183,
  -38.8245,
  -38.8235,
  -38.8165,
  -38.8046,
  -38.7892,
  -38.7718,
  -38.7525,
  -38.7339,
  -38.7159,
  -38.6996,
  -38.6899,
  -38.6914,
  -38.7055,
  -38.7361,
  -38.783,
  -38.8441,
  -38.9237,
  -39.0199,
  -39.1295,
  -39.2518,
  -39.3829,
  -39.5222,
  -39.6717,
  -39.8306,
  -39.9965,
  -40.1686,
  -40.3447,
  -40.5235,
  -40.7036,
  -40.8833,
  -41.0599,
  -41.2312,
  -41.3949,
  -41.5502,
  -41.6947,
  -41.8267,
  -41.945,
  -42.0524,
  -42.1492,
  -42.2374,
  -42.3182,
  -42.3931,
  -42.4621,
  -42.5238,
  -42.5767,
  -42.6197,
  -42.6509,
  -42.6703,
  -42.6781,
  -42.6739,
  -42.6585,
  -42.6337,
  -42.5995,
  -42.5609,
  -42.5189,
  -42.4751,
  -42.4324,
  -42.3929,
  -42.3596,
  -42.3355,
  -42.3223,
  -42.32,
  -42.3271,
  -42.3418,
  -42.3644,
  -42.3898,
  -42.4172,
  -42.445,
  -42.473,
  -42.4967,
  -42.5172,
  -42.5334,
  -42.5451,
  -42.5521,
  -42.5542,
  -42.5519,
  -42.5456,
  -42.5356,
  -42.5222,
  -42.5061,
  -42.4863,
  -42.4625,
  -42.4331,
  -42.3979,
  -42.3567,
  -42.3093,
  -42.2562,
  -42.1975,
  -42.1363,
  -42.0733,
  -42.0114,
  -41.9532,
  -41.8999,
  -41.8504,
  -41.8036,
  -41.7532,
  -41.6975,
  -41.6347,
  -41.5643,
  -41.4833,
  -41.4033,
  -41.3217,
  -41.2392,
  -41.1562,
  -41.0737,
  -40.985,
  -40.8927,
  -40.8012,
  -40.7108,
  -40.6255,
  -40.5282,
  -40.4396,
  -40.3498,
  -40.2645,
  -40.1725,
  -40.0992,
  -40.0317,
  -39.9796,
  -39.9384,
  -39.9031,
  -39.857,
  -39.7971,
  -39.735,
  -39.7032,
  -39.6634,
  -39.606,
  -39.5659,
  -39.5178,
  -39.4761,
  -39.4442,
  -39.4164,
  -39.4076,
  -39.4289,
  -39.4412,
  -39.4114,
  -39.3747,
  -39.3442,
  -39.3095,
  -39.2626,
  -39.1993,
  -39.1316,
  -39.064,
  -38.9984,
  -38.9263,
  -38.8876,
  -38.8974,
  -38.872,
  -38.8345,
  -38.8182,
  -38.8137,
  -38.7666,
  -38.7315,
  -38.7218,
  -38.7019,
  -38.6786,
  -38.6668,
  -38.6494,
  -38.6496,
  -38.6686,
  -38.701,
  -38.7489,
  -38.7975,
  -38.8405,
  -38.8659,
  -38.8852,
  -38.8947,
  -38.9307,
  -38.9809,
  -39.0273,
  -39.078,
  -39.1354,
  -39.2224,
  -39.3114,
  -39.3854,
  -39.4468,
  -39.4984,
  -39.5452,
  -39.5874,
  -39.634,
  -39.6872,
  -39.7476,
  -39.803,
  -39.854,
  -39.9028,
  -39.9493,
  -39.9988,
  -40.057,
  -40.1261,
  -40.2084,
  -40.2968,
  -40.3806,
  -40.4616,
  -40.541,
  -40.6193,
  -40.6967,
  -40.7707,
  -40.8419,
  -40.9086,
  -40.9734,
  -41.0384,
  -41.1,
  -41.1601,
  -41.2181,
  -41.2641,
  -41.3051,
  -41.3387,
  -41.3694,
  -41.3997,
  -41.4341,
  -41.4718,
  -41.5103,
  -41.5484,
  -41.5844,
  -41.6172,
  -41.6444,
  -41.6731,
  -41.7023,
  -41.7338,
  -41.7694,
  -41.8096,
  -41.8533,
  -41.9001,
  -41.9497,
  -42.002,
  -42.0575,
  -42.1121,
  -42.1671,
  -42.2218,
  -42.277,
  -42.3323,
  -42.3894,
  -42.446,
  -42.5005,
  -42.5502,
  -42.5903,
  -42.6261,
  -42.6539,
  -42.6731,
  -42.6848,
  -42.693,
  -42.6944,
  -42.6919,
  -42.6881,
  -42.6839,
  -42.6802,
  -42.675,
  -42.6697,
  -42.665,
  -42.663,
  -42.668,
  -42.6798,
  -42.7033,
  -42.7408,
  -42.7933,
  -42.8599,
  -42.9424,
  -43.0372,
  -43.142,
  -43.2521,
  -43.3611,
  -43.4676,
  -43.5654,
  -43.6512,
  -43.7231,
  -43.783,
  -43.8315,
  -43.8714,
  -43.9082,
  -43.945,
  -43.9853,
  -44.0304,
  -44.0804,
  -44.1343,
  -44.1893,
  -44.2428,
  -44.293,
  -44.3379,
  -44.378,
  -44.4153,
  -44.4517,
  -44.4898,
  -44.5306,
  -44.5744,
  -44.6189,
  -44.6609,
  -44.6963,
  -44.722,
  -44.7348,
  -44.7336,
  -44.7182,
  -44.6903,
  -44.655,
  -44.615,
  -44.5758,
  -44.5396,
  -44.5076,
  -44.479,
  -38.7995,
  -38.8236,
  -38.8407,
  -38.849,
  -38.8496,
  -38.8425,
  -38.8301,
  -38.8132,
  -38.7939,
  -38.773,
  -38.7525,
  -38.7331,
  -38.7143,
  -38.698,
  -38.6898,
  -38.6919,
  -38.7071,
  -38.7393,
  -38.7847,
  -38.8456,
  -38.9208,
  -39.0122,
  -39.1154,
  -39.2292,
  -39.3537,
  -39.4888,
  -39.6335,
  -39.791,
  -39.9592,
  -40.1366,
  -40.3204,
  -40.5088,
  -40.6987,
  -40.8882,
  -41.0746,
  -41.2544,
  -41.4275,
  -41.5915,
  -41.7442,
  -41.8842,
  -42.0105,
  -42.124,
  -42.2258,
  -42.3174,
  -42.4006,
  -42.4761,
  -42.5439,
  -42.6036,
  -42.6527,
  -42.6902,
  -42.7147,
  -42.7255,
  -42.7247,
  -42.7109,
  -42.6845,
  -42.6477,
  -42.6013,
  -42.5486,
  -42.4921,
  -42.4331,
  -42.3751,
  -42.3207,
  -42.2737,
  -42.2379,
  -42.2147,
  -42.2035,
  -42.2049,
  -42.2137,
  -42.2328,
  -42.2568,
  -42.2852,
  -42.3167,
  -42.3474,
  -42.3755,
  -42.3989,
  -42.4179,
  -42.4323,
  -42.4415,
  -42.4452,
  -42.4445,
  -42.4395,
  -42.4302,
  -42.4172,
  -42.401,
  -42.3804,
  -42.3542,
  -42.3219,
  -42.2825,
  -42.2357,
  -42.1817,
  -42.1211,
  -42.0549,
  -41.9846,
  -41.9133,
  -41.8432,
  -41.7777,
  -41.7179,
  -41.6634,
  -41.6125,
  -41.5593,
  -41.5032,
  -41.4415,
  -41.3745,
  -41.2973,
  -41.2228,
  -41.1465,
  -41.0699,
  -40.9919,
  -40.9147,
  -40.8344,
  -40.7483,
  -40.661,
  -40.5706,
  -40.4844,
  -40.3956,
  -40.3083,
  -40.2162,
  -40.1284,
  -40.0384,
  -39.9541,
  -39.8815,
  -39.821,
  -39.7887,
  -39.7408,
  -39.6902,
  -39.6327,
  -39.5739,
  -39.5472,
  -39.5019,
  -39.4564,
  -39.422,
  -39.3729,
  -39.3442,
  -39.3062,
  -39.268,
  -39.2598,
  -39.2788,
  -39.2664,
  -39.2546,
  -39.2099,
  -39.1687,
  -39.1453,
  -39.1118,
  -39.0597,
  -38.987,
  -38.917,
  -38.8578,
  -38.8029,
  -38.7501,
  -38.7564,
  -38.7173,
  -38.6959,
  -38.6764,
  -38.6778,
  -38.6491,
  -38.6113,
  -38.5941,
  -38.5682,
  -38.5478,
  -38.5407,
  -38.5245,
  -38.5337,
  -38.548,
  -38.5781,
  -38.6165,
  -38.6756,
  -38.7118,
  -38.725,
  -38.7355,
  -38.7489,
  -38.7833,
  -38.8304,
  -38.8792,
  -38.9332,
  -38.9973,
  -39.0782,
  -39.1607,
  -39.2458,
  -39.3095,
  -39.3602,
  -39.4175,
  -39.4884,
  -39.5529,
  -39.6091,
  -39.6635,
  -39.7283,
  -39.784,
  -39.8419,
  -39.8957,
  -39.9499,
  -40.0145,
  -40.0922,
  -40.1797,
  -40.2728,
  -40.3616,
  -40.4518,
  -40.5352,
  -40.6126,
  -40.6907,
  -40.7682,
  -40.8393,
  -40.9069,
  -40.973,
  -41.0327,
  -41.0936,
  -41.1521,
  -41.2044,
  -41.2485,
  -41.2877,
  -41.3219,
  -41.3536,
  -41.3863,
  -41.4249,
  -41.4668,
  -41.5085,
  -41.5495,
  -41.5877,
  -41.6221,
  -41.6494,
  -41.6783,
  -41.7081,
  -41.7411,
  -41.7773,
  -41.8202,
  -41.8675,
  -41.9195,
  -41.9753,
  -42.0345,
  -42.098,
  -42.1622,
  -42.2282,
  -42.2942,
  -42.3614,
  -42.4289,
  -42.4968,
  -42.5642,
  -42.6283,
  -42.686,
  -42.7346,
  -42.7765,
  -42.8087,
  -42.8317,
  -42.8473,
  -42.8578,
  -42.8623,
  -42.8625,
  -42.8608,
  -42.8578,
  -42.8533,
  -42.8472,
  -42.8406,
  -42.8336,
  -42.8288,
  -42.8304,
  -42.841,
  -42.8641,
  -42.9009,
  -42.9548,
  -43.0225,
  -43.1041,
  -43.1961,
  -43.2939,
  -43.3946,
  -43.4914,
  -43.5822,
  -43.6624,
  -43.7298,
  -43.783,
  -43.824,
  -43.8547,
  -43.8788,
  -43.9004,
  -43.9238,
  -43.9524,
  -43.9883,
  -44.0309,
  -44.0809,
  -44.134,
  -44.1891,
  -44.2427,
  -44.2934,
  -44.3418,
  -44.3893,
  -44.4364,
  -44.4839,
  -44.5328,
  -44.5814,
  -44.6266,
  -44.6652,
  -44.6949,
  -44.7109,
  -44.7119,
  -44.6973,
  -44.6687,
  -44.6297,
  -44.5844,
  -44.5379,
  -44.4946,
  -44.458,
  -44.4281,
  -44.4034,
  -38.8342,
  -38.8537,
  -38.866,
  -38.8702,
  -38.8672,
  -38.8569,
  -38.8403,
  -38.8202,
  -38.7981,
  -38.7753,
  -38.7536,
  -38.7334,
  -38.7148,
  -38.6989,
  -38.6895,
  -38.6926,
  -38.7094,
  -38.7403,
  -38.7842,
  -38.8422,
  -38.9128,
  -38.9961,
  -39.0906,
  -39.1966,
  -39.313,
  -39.4411,
  -39.5816,
  -39.7362,
  -39.9048,
  -40.0862,
  -40.2764,
  -40.4739,
  -40.6747,
  -40.8757,
  -41.0737,
  -41.2661,
  -41.4505,
  -41.6253,
  -41.7886,
  -41.9382,
  -42.0739,
  -42.1951,
  -42.3034,
  -42.3996,
  -42.4855,
  -42.5611,
  -42.6285,
  -42.6857,
  -42.7307,
  -42.7628,
  -42.781,
  -42.7856,
  -42.7761,
  -42.7526,
  -42.7153,
  -42.6663,
  -42.6072,
  -42.5408,
  -42.4695,
  -42.3964,
  -42.3238,
  -42.2551,
  -42.194,
  -42.1462,
  -42.113,
  -42.0935,
  -42.0888,
  -42.0952,
  -42.1119,
  -42.1352,
  -42.1628,
  -42.1973,
  -42.2323,
  -42.2644,
  -42.2924,
  -42.3146,
  -42.3314,
  -42.3426,
  -42.3492,
  -42.3498,
  -42.3468,
  -42.3392,
  -42.3279,
  -42.3122,
  -42.2917,
  -42.2645,
  -42.2294,
  -42.1864,
  -42.1345,
  -42.0741,
  -42.0054,
  -41.9306,
  -41.8516,
  -41.7715,
  -41.6937,
  -41.6213,
  -41.5552,
  -41.4939,
  -41.4381,
  -41.3823,
  -41.325,
  -41.2638,
  -41.1991,
  -41.1272,
  -41.0568,
  -40.9856,
  -40.9139,
  -40.8417,
  -40.7694,
  -40.6946,
  -40.6108,
  -40.5252,
  -40.4373,
  -40.3484,
  -40.2582,
  -40.1784,
  -40.0975,
  -40.0124,
  -39.9281,
  -39.8342,
  -39.7576,
  -39.6945,
  -39.6456,
  -39.5924,
  -39.5314,
  -39.4857,
  -39.4274,
  -39.3955,
  -39.3625,
  -39.3188,
  -39.2906,
  -39.2454,
  -39.2146,
  -39.1791,
  -39.1624,
  -39.1509,
  -39.142,
  -39.1096,
  -39.1011,
  -39.0792,
  -39.0441,
  -39.004,
  -38.9728,
  -38.9146,
  -38.8386,
  -38.7713,
  -38.7244,
  -38.6826,
  -38.6449,
  -38.6496,
  -38.6222,
  -38.6041,
  -38.5912,
  -38.5783,
  -38.5719,
  -38.5416,
  -38.5097,
  -38.4801,
  -38.4653,
  -38.4571,
  -38.4489,
  -38.4543,
  -38.4693,
  -38.4907,
  -38.5276,
  -38.5697,
  -38.5939,
  -38.5981,
  -38.6043,
  -38.6376,
  -38.6662,
  -38.7077,
  -38.7521,
  -38.8059,
  -38.8696,
  -38.9449,
  -39.0339,
  -39.1124,
  -39.1764,
  -39.2346,
  -39.3106,
  -39.392,
  -39.4685,
  -39.5356,
  -39.5955,
  -39.6624,
  -39.7305,
  -39.7956,
  -39.8537,
  -39.918,
  -39.9881,
  -40.0793,
  -40.1712,
  -40.2634,
  -40.3597,
  -40.453,
  -40.5397,
  -40.62,
  -40.6987,
  -40.7745,
  -40.8469,
  -40.915,
  -40.9808,
  -41.0409,
  -41.0989,
  -41.1515,
  -41.1985,
  -41.2402,
  -41.279,
  -41.3137,
  -41.3488,
  -41.3851,
  -41.4262,
  -41.4717,
  -41.5151,
  -41.5584,
  -41.5988,
  -41.6351,
  -41.6648,
  -41.6961,
  -41.7284,
  -41.7631,
  -41.8036,
  -41.8502,
  -41.9029,
  -41.9614,
  -42.0244,
  -42.0925,
  -42.1648,
  -42.2395,
  -42.3163,
  -42.3938,
  -42.4722,
  -42.5509,
  -42.6295,
  -42.7065,
  -42.7791,
  -42.8442,
  -42.8997,
  -42.9462,
  -42.9826,
  -43.0095,
  -43.0282,
  -43.0416,
  -43.0484,
  -43.0516,
  -43.0523,
  -43.0513,
  -43.0479,
  -43.0424,
  -43.0347,
  -43.0259,
  -43.019,
  -43.0184,
  -43.027,
  -43.0485,
  -43.0855,
  -43.1376,
  -43.203,
  -43.2794,
  -43.3636,
  -43.4504,
  -43.536,
  -43.6156,
  -43.687,
  -43.7465,
  -43.7926,
  -43.8255,
  -43.8471,
  -43.8599,
  -43.8682,
  -43.8762,
  -43.8876,
  -43.9074,
  -43.9366,
  -43.9761,
  -44.0241,
  -44.078,
  -44.1369,
  -44.1961,
  -44.2545,
  -44.3119,
  -44.3689,
  -44.4253,
  -44.4798,
  -44.5343,
  -44.5859,
  -44.6312,
  -44.6663,
  -44.6897,
  -44.6976,
  -44.6887,
  -44.6638,
  -44.6253,
  -44.577,
  -44.5244,
  -44.4727,
  -44.4269,
  -44.3906,
  -44.3636,
  -44.3433,
  -38.8594,
  -38.875,
  -38.884,
  -38.8855,
  -38.8799,
  -38.8678,
  -38.8493,
  -38.8275,
  -38.804,
  -38.7798,
  -38.7577,
  -38.7374,
  -38.7193,
  -38.7053,
  -38.6954,
  -38.699,
  -38.7148,
  -38.7439,
  -38.7856,
  -38.838,
  -38.901,
  -38.9761,
  -39.0617,
  -39.1583,
  -39.2657,
  -39.3865,
  -39.521,
  -39.6716,
  -39.8395,
  -40.0231,
  -40.2198,
  -40.4256,
  -40.6368,
  -40.8498,
  -41.0605,
  -41.2658,
  -41.4628,
  -41.6496,
  -41.8247,
  -41.9856,
  -42.13,
  -42.2608,
  -42.3765,
  -42.4784,
  -42.5678,
  -42.6458,
  -42.7123,
  -42.767,
  -42.8084,
  -42.8355,
  -42.8478,
  -42.8455,
  -42.8278,
  -42.7948,
  -42.7469,
  -42.6869,
  -42.6151,
  -42.5362,
  -42.4518,
  -42.3651,
  -42.2789,
  -42.1968,
  -42.1243,
  -42.065,
  -42.0223,
  -41.9955,
  -41.9834,
  -41.9864,
  -42.0004,
  -42.0245,
  -42.0554,
  -42.0919,
  -42.13,
  -42.1654,
  -42.1972,
  -42.2229,
  -42.2426,
  -42.2567,
  -42.2651,
  -42.2696,
  -42.269,
  -42.2637,
  -42.2541,
  -42.2394,
  -42.2186,
  -42.1901,
  -42.1532,
  -42.1067,
  -42.0498,
  -41.9828,
  -41.9068,
  -41.8223,
  -41.7348,
  -41.6467,
  -41.5617,
  -41.4828,
  -41.411,
  -41.3454,
  -41.2852,
  -41.2258,
  -41.1671,
  -41.1067,
  -41.0437,
  -40.9751,
  -40.9078,
  -40.8401,
  -40.7722,
  -40.7045,
  -40.6363,
  -40.5656,
  -40.4882,
  -40.4076,
  -40.3267,
  -40.2466,
  -40.162,
  -40.0871,
  -40.0047,
  -39.919,
  -39.8215,
  -39.7256,
  -39.6461,
  -39.5802,
  -39.5343,
  -39.4786,
  -39.423,
  -39.3693,
  -39.3161,
  -39.2776,
  -39.2474,
  -39.201,
  -39.1631,
  -39.1277,
  -39.0977,
  -39.0695,
  -39.0476,
  -39.0371,
  -39.039,
  -39.0101,
  -38.9745,
  -38.962,
  -38.9396,
  -38.9081,
  -38.8657,
  -38.8085,
  -38.747,
  -38.6834,
  -38.6371,
  -38.6072,
  -38.586,
  -38.5918,
  -38.5811,
  -38.569,
  -38.5801,
  -38.5587,
  -38.5396,
  -38.5084,
  -38.4763,
  -38.4488,
  -38.4352,
  -38.4131,
  -38.4025,
  -38.404,
  -38.4155,
  -38.4327,
  -38.4527,
  -38.4861,
  -38.5038,
  -38.5127,
  -38.5059,
  -38.5301,
  -38.5643,
  -38.5994,
  -38.6387,
  -38.6867,
  -38.742,
  -38.8101,
  -38.8879,
  -38.9744,
  -39.0523,
  -39.1249,
  -39.2185,
  -39.3079,
  -39.3878,
  -39.4548,
  -39.5187,
  -39.5992,
  -39.6758,
  -39.7525,
  -39.8242,
  -39.9021,
  -39.9794,
  -40.069,
  -40.1646,
  -40.2631,
  -40.366,
  -40.4621,
  -40.553,
  -40.635,
  -40.7154,
  -40.7898,
  -40.8614,
  -40.9283,
  -40.9925,
  -41.05,
  -41.1061,
  -41.1564,
  -41.2014,
  -41.2429,
  -41.283,
  -41.3206,
  -41.3598,
  -41.402,
  -41.4472,
  -41.4955,
  -41.5404,
  -41.5842,
  -41.6264,
  -41.6668,
  -41.7006,
  -41.7356,
  -41.7715,
  -41.8106,
  -41.8545,
  -41.9061,
  -41.9659,
  -42.0316,
  -42.1033,
  -42.1802,
  -42.2619,
  -42.3462,
  -42.4334,
  -42.5216,
  -42.609,
  -42.6979,
  -42.7857,
  -42.8712,
  -42.9504,
  -43.0218,
  -43.0836,
  -43.1348,
  -43.1748,
  -43.2056,
  -43.2279,
  -43.2438,
  -43.2543,
  -43.26,
  -43.2628,
  -43.2634,
  -43.261,
  -43.2555,
  -43.2471,
  -43.237,
  -43.2283,
  -43.2254,
  -43.2315,
  -43.2505,
  -43.2843,
  -43.3322,
  -43.3915,
  -43.4594,
  -43.5315,
  -43.6033,
  -43.6707,
  -43.7298,
  -43.779,
  -43.816,
  -43.84,
  -43.852,
  -43.8546,
  -43.85,
  -43.8446,
  -43.8413,
  -43.8446,
  -43.8579,
  -43.8834,
  -43.9222,
  -43.9713,
  -44.0286,
  -44.092,
  -44.1579,
  -44.2243,
  -44.2901,
  -44.3551,
  -44.4187,
  -44.48,
  -44.5379,
  -44.5902,
  -44.6345,
  -44.6665,
  -44.6847,
  -44.6864,
  -44.6706,
  -44.6386,
  -44.593,
  -44.5385,
  -44.4806,
  -44.4251,
  -44.3776,
  -44.3414,
  -44.3165,
  -44.3,
  -38.8761,
  -38.8889,
  -38.8959,
  -38.8964,
  -38.8903,
  -38.8764,
  -38.8582,
  -38.8368,
  -38.8139,
  -38.7914,
  -38.7701,
  -38.75,
  -38.733,
  -38.7203,
  -38.7135,
  -38.7163,
  -38.7296,
  -38.7551,
  -38.7918,
  -38.8383,
  -38.894,
  -38.9609,
  -39.0378,
  -39.1242,
  -39.2225,
  -39.3367,
  -39.4654,
  -39.6107,
  -39.7752,
  -39.9586,
  -40.1578,
  -40.3696,
  -40.5897,
  -40.8136,
  -41.0358,
  -41.2541,
  -41.4645,
  -41.6645,
  -41.8518,
  -42.0243,
  -42.1805,
  -42.3204,
  -42.4442,
  -42.5521,
  -42.6452,
  -42.7248,
  -42.7908,
  -42.8431,
  -42.8806,
  -42.9036,
  -42.9105,
  -42.9019,
  -42.8767,
  -42.8351,
  -42.7779,
  -42.7078,
  -42.6265,
  -42.5372,
  -42.4416,
  -42.3434,
  -42.245,
  -42.1511,
  -42.0673,
  -41.9976,
  -41.9461,
  -41.9122,
  -41.8954,
  -41.8929,
  -41.9058,
  -41.9286,
  -41.9609,
  -41.9996,
  -42.0405,
  -42.0807,
  -42.1169,
  -42.1463,
  -42.1692,
  -42.1862,
  -42.1973,
  -42.2037,
  -42.2045,
  -42.2011,
  -42.1929,
  -42.1791,
  -42.1571,
  -42.128,
  -42.0896,
  -42.0398,
  -41.9785,
  -41.9056,
  -41.8225,
  -41.732,
  -41.6365,
  -41.5415,
  -41.4502,
  -41.3652,
  -41.2877,
  -41.217,
  -41.1526,
  -41.0906,
  -41.0302,
  -40.9704,
  -40.9088,
  -40.8419,
  -40.7767,
  -40.711,
  -40.6454,
  -40.5802,
  -40.5151,
  -40.4493,
  -40.3782,
  -40.3044,
  -40.229,
  -40.1554,
  -40.0805,
  -40.0074,
  -39.931,
  -39.8471,
  -39.7464,
  -39.6553,
  -39.57,
  -39.4974,
  -39.4445,
  -39.3988,
  -39.3537,
  -39.3011,
  -39.2492,
  -39.2025,
  -39.1671,
  -39.1273,
  -39.0794,
  -39.0345,
  -38.9983,
  -38.9731,
  -38.9528,
  -38.9499,
  -38.9437,
  -38.9339,
  -38.9025,
  -38.8848,
  -38.8726,
  -38.8662,
  -38.8323,
  -38.7982,
  -38.7512,
  -38.6994,
  -38.6434,
  -38.6075,
  -38.5938,
  -38.5965,
  -38.6212,
  -38.6166,
  -38.616,
  -38.5956,
  -38.5636,
  -38.5367,
  -38.4941,
  -38.4696,
  -38.4568,
  -38.4235,
  -38.3864,
  -38.3748,
  -38.3727,
  -38.3776,
  -38.3839,
  -38.4017,
  -38.4356,
  -38.4437,
  -38.4491,
  -38.4627,
  -38.4885,
  -38.5157,
  -38.5478,
  -38.5918,
  -38.6387,
  -38.6805,
  -38.757,
  -38.8573,
  -38.9424,
  -39.0194,
  -39.1293,
  -39.2302,
  -39.3112,
  -39.3898,
  -39.4537,
  -39.5364,
  -39.6219,
  -39.7103,
  -39.7981,
  -39.8935,
  -39.9891,
  -40.0814,
  -40.176,
  -40.2774,
  -40.381,
  -40.4811,
  -40.5739,
  -40.6582,
  -40.7395,
  -40.8143,
  -40.8852,
  -40.9521,
  -41.0149,
  -41.0713,
  -41.1254,
  -41.1746,
  -41.2193,
  -41.2614,
  -41.3037,
  -41.3461,
  -41.3915,
  -41.4385,
  -41.4871,
  -41.5376,
  -41.5809,
  -41.625,
  -41.6703,
  -41.7179,
  -41.7591,
  -41.8005,
  -41.8417,
  -41.885,
  -41.9355,
  -41.9942,
  -42.0615,
  -42.1355,
  -42.2157,
  -42.301,
  -42.3908,
  -42.4837,
  -42.5792,
  -42.6759,
  -42.7725,
  -42.8694,
  -42.9643,
  -43.0557,
  -43.1408,
  -43.2169,
  -43.2831,
  -43.3385,
  -43.3825,
  -43.4161,
  -43.4415,
  -43.4597,
  -43.4723,
  -43.4799,
  -43.4841,
  -43.4854,
  -43.4831,
  -43.4777,
  -43.4687,
  -43.4574,
  -43.447,
  -43.4413,
  -43.4447,
  -43.4592,
  -43.4881,
  -43.529,
  -43.5793,
  -43.6354,
  -43.6928,
  -43.7464,
  -43.7932,
  -43.8301,
  -43.8562,
  -43.87,
  -43.872,
  -43.8643,
  -43.8496,
  -43.832,
  -43.8158,
  -43.8048,
  -43.8031,
  -43.8141,
  -43.8396,
  -43.8792,
  -43.9308,
  -43.9924,
  -44.0606,
  -44.1327,
  -44.2056,
  -44.2779,
  -44.3492,
  -44.4175,
  -44.4819,
  -44.5412,
  -44.5932,
  -44.6354,
  -44.6648,
  -44.6794,
  -44.6772,
  -44.6574,
  -44.6217,
  -44.5724,
  -44.5142,
  -44.453,
  -44.3952,
  -44.3464,
  -44.3101,
  -44.2863,
  -44.2698,
  -38.8861,
  -38.8973,
  -38.9036,
  -38.9043,
  -38.8989,
  -38.8873,
  -38.8714,
  -38.8521,
  -38.8316,
  -38.8112,
  -38.7916,
  -38.773,
  -38.7571,
  -38.7454,
  -38.7391,
  -38.7418,
  -38.7535,
  -38.7753,
  -38.8077,
  -38.8489,
  -38.899,
  -38.9589,
  -39.0286,
  -39.1075,
  -39.1979,
  -39.3021,
  -39.4238,
  -39.562,
  -39.721,
  -39.9002,
  -40.0991,
  -40.3135,
  -40.5394,
  -40.7721,
  -41.0064,
  -41.2374,
  -41.4609,
  -41.6733,
  -41.8731,
  -42.0569,
  -42.2234,
  -42.3723,
  -42.5036,
  -42.6173,
  -42.7141,
  -42.7939,
  -42.8593,
  -42.9104,
  -42.9461,
  -42.9655,
  -42.969,
  -42.9556,
  -42.9241,
  -42.8752,
  -42.8099,
  -42.7315,
  -42.6418,
  -42.5439,
  -42.4393,
  -42.332,
  -42.2241,
  -42.1193,
  -42.026,
  -41.9477,
  -41.8887,
  -41.8478,
  -41.827,
  -41.8224,
  -41.8323,
  -41.8542,
  -41.8865,
  -41.9262,
  -41.9694,
  -42.0126,
  -42.0521,
  -42.0855,
  -42.1118,
  -42.1313,
  -42.1436,
  -42.1513,
  -42.1533,
  -42.1505,
  -42.1426,
  -42.1289,
  -42.1077,
  -42.0781,
  -42.0382,
  -41.9859,
  -41.921,
  -41.8433,
  -41.7546,
  -41.6579,
  -41.5564,
  -41.4558,
  -41.3587,
  -41.2683,
  -41.1847,
  -41.1092,
  -41.0405,
  -40.9762,
  -40.9145,
  -40.8547,
  -40.794,
  -40.7298,
  -40.6657,
  -40.6008,
  -40.5361,
  -40.4714,
  -40.4075,
  -40.3447,
  -40.2773,
  -40.2154,
  -40.1459,
  -40.0818,
  -40.0112,
  -39.9381,
  -39.8665,
  -39.7868,
  -39.7089,
  -39.6279,
  -39.5469,
  -39.4777,
  -39.4263,
  -39.3863,
  -39.3502,
  -39.2921,
  -39.2486,
  -39.2029,
  -39.1506,
  -39.1062,
  -39.0566,
  -39.0063,
  -38.9671,
  -38.9369,
  -38.9086,
  -38.9013,
  -38.8862,
  -38.8692,
  -38.8521,
  -38.8596,
  -38.8662,
  -38.8507,
  -38.8436,
  -38.8327,
  -38.7973,
  -38.7707,
  -38.7258,
  -38.679,
  -38.662,
  -38.6634,
  -38.6931,
  -38.6892,
  -38.666,
  -38.6435,
  -38.6053,
  -38.5706,
  -38.5331,
  -38.5172,
  -38.4922,
  -38.454,
  -38.4129,
  -38.3806,
  -38.3656,
  -38.3549,
  -38.3477,
  -38.3467,
  -38.362,
  -38.392,
  -38.4015,
  -38.4159,
  -38.4347,
  -38.4555,
  -38.4859,
  -38.5214,
  -38.5559,
  -38.5971,
  -38.6604,
  -38.7533,
  -38.8458,
  -38.9545,
  -39.0652,
  -39.1688,
  -39.2527,
  -39.3339,
  -39.4084,
  -39.4962,
  -39.5923,
  -39.6907,
  -39.7873,
  -39.8919,
  -39.9978,
  -40.1008,
  -40.2042,
  -40.3071,
  -40.4104,
  -40.5117,
  -40.6064,
  -40.693,
  -40.7775,
  -40.8542,
  -40.9257,
  -40.9923,
  -41.0541,
  -41.1093,
  -41.1618,
  -41.2095,
  -41.2529,
  -41.296,
  -41.3422,
  -41.3894,
  -41.4368,
  -41.4872,
  -41.5396,
  -41.5945,
  -41.6418,
  -41.6892,
  -41.7402,
  -41.7947,
  -41.8446,
  -41.8935,
  -41.9415,
  -41.9922,
  -42.0545,
  -42.121,
  -42.1963,
  -42.2781,
  -42.3659,
  -42.4583,
  -42.5546,
  -42.6535,
  -42.7547,
  -42.8567,
  -42.9586,
  -43.0605,
  -43.1598,
  -43.2548,
  -43.3431,
  -43.4224,
  -43.4917,
  -43.5496,
  -43.5965,
  -43.6329,
  -43.6597,
  -43.6799,
  -43.694,
  -43.7025,
  -43.7069,
  -43.7077,
  -43.7052,
  -43.6993,
  -43.6895,
  -43.677,
  -43.6649,
  -43.6568,
  -43.6568,
  -43.6677,
  -43.6899,
  -43.7216,
  -43.7604,
  -43.8022,
  -43.8425,
  -43.8765,
  -43.9016,
  -43.9161,
  -43.9191,
  -43.9111,
  -43.8924,
  -43.8668,
  -43.8375,
  -43.809,
  -43.7856,
  -43.7708,
  -43.768,
  -43.7796,
  -43.8068,
  -43.8491,
  -43.9037,
  -43.9684,
  -44.0409,
  -44.1172,
  -44.195,
  -44.2713,
  -44.3457,
  -44.4156,
  -44.4813,
  -44.5403,
  -44.5909,
  -44.6312,
  -44.6586,
  -44.6713,
  -44.6676,
  -44.646,
  -44.6092,
  -44.559,
  -44.5007,
  -44.4383,
  -44.3796,
  -44.3298,
  -44.2926,
  -44.2678,
  -44.252,
  -38.8954,
  -38.9063,
  -38.9131,
  -38.9147,
  -38.9109,
  -38.9024,
  -38.8898,
  -38.8744,
  -38.8575,
  -38.8394,
  -38.822,
  -38.8057,
  -38.792,
  -38.7826,
  -38.778,
  -38.7802,
  -38.7914,
  -38.8099,
  -38.8372,
  -38.8733,
  -38.9179,
  -38.9711,
  -39.0337,
  -39.1066,
  -39.1897,
  -39.2866,
  -39.3998,
  -39.5318,
  -39.6839,
  -39.8585,
  -40.054,
  -40.2675,
  -40.496,
  -40.7343,
  -40.9777,
  -41.2193,
  -41.4543,
  -41.679,
  -41.8897,
  -42.0827,
  -42.2584,
  -42.4153,
  -42.5531,
  -42.6714,
  -42.7717,
  -42.8544,
  -42.9206,
  -42.9707,
  -43.0053,
  -43.0227,
  -43.0231,
  -43.0057,
  -42.9693,
  -42.9153,
  -42.8436,
  -42.7577,
  -42.6615,
  -42.5566,
  -42.4445,
  -42.33,
  -42.2148,
  -42.1041,
  -42.0035,
  -41.9181,
  -41.851,
  -41.8014,
  -41.7774,
  -41.7725,
  -41.7789,
  -41.8035,
  -41.8337,
  -41.872,
  -41.9151,
  -41.9604,
  -42.0029,
  -42.0398,
  -42.0695,
  -42.0914,
  -42.1059,
  -42.1144,
  -42.1166,
  -42.1132,
  -42.105,
  -42.091,
  -42.0694,
  -42.0389,
  -41.9976,
  -41.9435,
  -41.8757,
  -41.7946,
  -41.7009,
  -41.5997,
  -41.4937,
  -41.3886,
  -41.2871,
  -41.1921,
  -41.1048,
  -41.025,
  -40.9523,
  -40.885,
  -40.8224,
  -40.7617,
  -40.7012,
  -40.6384,
  -40.5747,
  -40.5101,
  -40.4442,
  -40.3793,
  -40.3147,
  -40.252,
  -40.1896,
  -40.1279,
  -40.0711,
  -40.0093,
  -39.9457,
  -39.8806,
  -39.8129,
  -39.7455,
  -39.6762,
  -39.6102,
  -39.5483,
  -39.4962,
  -39.4485,
  -39.3983,
  -39.3633,
  -39.3029,
  -39.2777,
  -39.247,
  -39.1997,
  -39.1504,
  -39.0956,
  -39.0365,
  -38.9995,
  -38.9777,
  -38.9182,
  -38.8882,
  -38.8753,
  -38.8768,
  -38.8679,
  -38.8677,
  -38.8825,
  -38.8833,
  -38.8616,
  -38.863,
  -38.8571,
  -38.8302,
  -38.8055,
  -38.7822,
  -38.7714,
  -38.7685,
  -38.7692,
  -38.7477,
  -38.7153,
  -38.689,
  -38.6367,
  -38.6155,
  -38.5819,
  -38.56,
  -38.5524,
  -38.5207,
  -38.4806,
  -38.4354,
  -38.3969,
  -38.3694,
  -38.3423,
  -38.3265,
  -38.321,
  -38.3331,
  -38.3503,
  -38.3656,
  -38.3818,
  -38.3996,
  -38.4229,
  -38.4512,
  -38.4732,
  -38.5074,
  -38.5665,
  -38.6513,
  -38.7684,
  -38.8881,
  -39.0089,
  -39.1172,
  -39.2066,
  -39.2987,
  -39.3853,
  -39.4861,
  -39.5915,
  -39.6967,
  -39.8017,
  -39.9111,
  -40.028,
  -40.1421,
  -40.2523,
  -40.3558,
  -40.4582,
  -40.5592,
  -40.6546,
  -40.7451,
  -40.8336,
  -40.9142,
  -40.987,
  -41.0528,
  -41.1139,
  -41.1684,
  -41.2183,
  -41.2631,
  -41.3058,
  -41.3485,
  -41.3945,
  -41.4418,
  -41.4962,
  -41.5545,
  -41.6166,
  -41.6785,
  -41.7354,
  -41.7908,
  -41.8466,
  -41.9073,
  -41.9658,
  -42.0247,
  -42.082,
  -42.143,
  -42.2108,
  -42.2858,
  -42.3683,
  -42.4574,
  -42.5519,
  -42.6497,
  -42.75,
  -42.8521,
  -42.9558,
  -43.0584,
  -43.1619,
  -43.2648,
  -43.3651,
  -43.4609,
  -43.5499,
  -43.6297,
  -43.6999,
  -43.7591,
  -43.8075,
  -43.8458,
  -43.8756,
  -43.8977,
  -43.9128,
  -43.9214,
  -43.9257,
  -43.9266,
  -43.9233,
  -43.9158,
  -43.9046,
  -43.8907,
  -43.8774,
  -43.8672,
  -43.8633,
  -43.8681,
  -43.882,
  -43.903,
  -43.9278,
  -43.9536,
  -43.9755,
  -43.9895,
  -43.9929,
  -43.985,
  -43.9662,
  -43.9375,
  -43.9009,
  -43.8601,
  -43.8186,
  -43.7825,
  -43.7553,
  -43.74,
  -43.7386,
  -43.7531,
  -43.783,
  -43.8265,
  -43.8833,
  -43.9505,
  -44.0251,
  -44.1039,
  -44.1836,
  -44.2623,
  -44.3378,
  -44.4091,
  -44.4744,
  -44.5323,
  -44.5815,
  -44.6202,
  -44.6466,
  -44.6587,
  -44.6549,
  -44.6346,
  -44.5986,
  -44.5507,
  -44.4936,
  -44.4332,
  -44.3747,
  -44.3245,
  -44.2858,
  -44.2584,
  -44.2399,
  -38.9075,
  -38.9193,
  -38.9273,
  -38.9306,
  -38.9283,
  -38.9236,
  -38.9153,
  -38.9043,
  -38.8919,
  -38.8783,
  -38.8641,
  -38.8509,
  -38.8398,
  -38.8322,
  -38.8291,
  -38.8311,
  -38.8401,
  -38.8561,
  -38.8796,
  -38.9102,
  -38.9496,
  -38.9982,
  -39.0555,
  -39.1224,
  -39.2019,
  -39.2935,
  -39.4005,
  -39.5252,
  -39.6705,
  -39.8381,
  -40.0277,
  -40.2381,
  -40.4657,
  -40.7076,
  -40.9548,
  -41.2047,
  -41.4492,
  -41.6833,
  -41.9037,
  -42.106,
  -42.2892,
  -42.4524,
  -42.5954,
  -42.7177,
  -42.8213,
  -42.9063,
  -42.9738,
  -43.0244,
  -43.0585,
  -43.0751,
  -43.0725,
  -43.0523,
  -43.0129,
  -42.9556,
  -42.8801,
  -42.7914,
  -42.6903,
  -42.5807,
  -42.4638,
  -42.345,
  -42.2253,
  -42.1101,
  -42.005,
  -41.9135,
  -41.8388,
  -41.7841,
  -41.7532,
  -41.744,
  -41.7517,
  -41.77,
  -41.8019,
  -41.8382,
  -41.8813,
  -41.9272,
  -41.9716,
  -42.0108,
  -42.0434,
  -42.0672,
  -42.083,
  -42.0918,
  -42.0934,
  -42.0893,
  -42.08,
  -42.0647,
  -42.041,
  -42.0094,
  -41.9671,
  -41.9118,
  -41.8426,
  -41.7596,
  -41.6643,
  -41.5599,
  -41.4518,
  -41.3434,
  -41.2384,
  -41.1397,
  -41.0481,
  -40.9634,
  -40.8864,
  -40.8162,
  -40.7513,
  -40.6888,
  -40.6263,
  -40.5635,
  -40.4996,
  -40.4342,
  -40.367,
  -40.3007,
  -40.2358,
  -40.1732,
  -40.1136,
  -40.0602,
  -40.0047,
  -39.9454,
  -39.8875,
  -39.8292,
  -39.7728,
  -39.7181,
  -39.6658,
  -39.6093,
  -39.5612,
  -39.5175,
  -39.4759,
  -39.4342,
  -39.3906,
  -39.3419,
  -39.3116,
  -39.2856,
  -39.2572,
  -39.2088,
  -39.153,
  -39.0905,
  -39.0623,
  -39.0261,
  -38.9676,
  -38.9325,
  -38.9259,
  -38.9248,
  -38.948,
  -38.938,
  -38.9379,
  -38.9332,
  -38.9198,
  -38.9076,
  -38.907,
  -38.9118,
  -38.8948,
  -38.8668,
  -38.8562,
  -38.8529,
  -38.8433,
  -38.8129,
  -38.7822,
  -38.7479,
  -38.7055,
  -38.6822,
  -38.6579,
  -38.6314,
  -38.6168,
  -38.5875,
  -38.547,
  -38.5066,
  -38.4644,
  -38.4229,
  -38.3726,
  -38.3467,
  -38.3213,
  -38.3177,
  -38.3141,
  -38.328,
  -38.339,
  -38.3448,
  -38.3737,
  -38.4129,
  -38.4371,
  -38.4725,
  -38.5328,
  -38.6121,
  -38.7163,
  -38.826,
  -38.9624,
  -39.0802,
  -39.1825,
  -39.2842,
  -39.3887,
  -39.4993,
  -39.6162,
  -39.7315,
  -39.8446,
  -39.9617,
  -40.0794,
  -40.1971,
  -40.3081,
  -40.4125,
  -40.5153,
  -40.6181,
  -40.7188,
  -40.8164,
  -40.9107,
  -40.9965,
  -41.0738,
  -41.1415,
  -41.2021,
  -41.2561,
  -41.3052,
  -41.3491,
  -41.3898,
  -41.4311,
  -41.485,
  -41.544,
  -41.6015,
  -41.6684,
  -41.7325,
  -41.7974,
  -41.8591,
  -41.9233,
  -41.9881,
  -42.0541,
  -42.1196,
  -42.1863,
  -42.2525,
  -42.325,
  -42.4015,
  -42.484,
  -42.5737,
  -42.6692,
  -42.7683,
  -42.8695,
  -42.971,
  -43.073,
  -43.1756,
  -43.278,
  -43.3798,
  -43.4809,
  -43.5793,
  -43.6731,
  -43.7607,
  -43.8403,
  -43.9096,
  -43.9687,
  -44.0175,
  -44.0571,
  -44.0877,
  -44.1098,
  -44.1248,
  -44.133,
  -44.1365,
  -44.1349,
  -44.1292,
  -44.1197,
  -44.1063,
  -44.0904,
  -44.0739,
  -44.0605,
  -44.0509,
  -44.0482,
  -44.0525,
  -44.0615,
  -44.072,
  -44.0812,
  -44.0842,
  -44.0781,
  -44.0608,
  -44.0326,
  -43.9942,
  -43.9474,
  -43.8959,
  -43.8438,
  -43.7953,
  -43.7549,
  -43.7263,
  -43.7126,
  -43.7136,
  -43.7293,
  -43.7609,
  -43.8065,
  -43.8646,
  -43.9315,
  -44.0065,
  -44.0853,
  -44.1654,
  -44.2441,
  -44.3198,
  -44.3906,
  -44.4549,
  -44.5116,
  -44.5596,
  -44.5975,
  -44.6237,
  -44.6357,
  -44.6335,
  -44.6159,
  -44.5833,
  -44.5389,
  -44.4858,
  -44.4282,
  -44.3721,
  -44.3217,
  -44.2803,
  -44.2497,
  -44.227,
  -38.9266,
  -38.94,
  -38.9497,
  -38.956,
  -38.9581,
  -38.9571,
  -38.9531,
  -38.9466,
  -38.9387,
  -38.9289,
  -38.9177,
  -38.9072,
  -38.899,
  -38.8929,
  -38.8896,
  -38.8914,
  -38.8991,
  -38.913,
  -38.9338,
  -38.9624,
  -38.9986,
  -39.0434,
  -39.0971,
  -39.1605,
  -39.2352,
  -39.3223,
  -39.4237,
  -39.5428,
  -39.6819,
  -39.8413,
  -40.0243,
  -40.2297,
  -40.4548,
  -40.6964,
  -40.9472,
  -41.2009,
  -41.4512,
  -41.692,
  -41.9195,
  -42.1279,
  -42.3167,
  -42.4848,
  -42.6314,
  -42.7574,
  -42.8626,
  -42.95,
  -43.0196,
  -43.0713,
  -43.1061,
  -43.1223,
  -43.1196,
  -43.0979,
  -43.0575,
  -42.9996,
  -42.9225,
  -42.8322,
  -42.729,
  -42.6167,
  -42.4974,
  -42.3763,
  -42.2547,
  -42.1361,
  -42.0277,
  -41.9326,
  -41.8532,
  -41.7953,
  -41.7612,
  -41.7464,
  -41.75,
  -41.7638,
  -41.7915,
  -41.8245,
  -41.8656,
  -41.9115,
  -41.9561,
  -41.9971,
  -42.0307,
  -42.0563,
  -42.0722,
  -42.0811,
  -42.0821,
  -42.0767,
  -42.0659,
  -42.0488,
  -42.0246,
  -41.9919,
  -41.9487,
  -41.8932,
  -41.8238,
  -41.7406,
  -41.6446,
  -41.54,
  -41.4301,
  -41.3198,
  -41.2122,
  -41.1098,
  -41.0126,
  -40.9234,
  -40.8418,
  -40.7676,
  -40.699,
  -40.6339,
  -40.5705,
  -40.5071,
  -40.4423,
  -40.3758,
  -40.3078,
  -40.2399,
  -40.1742,
  -40.1114,
  -40.0531,
  -39.9976,
  -39.9406,
  -39.8822,
  -39.8264,
  -39.7762,
  -39.7326,
  -39.6902,
  -39.6525,
  -39.6095,
  -39.5716,
  -39.5376,
  -39.5033,
  -39.4701,
  -39.4268,
  -39.388,
  -39.3643,
  -39.336,
  -39.3106,
  -39.2655,
  -39.2248,
  -39.1913,
  -39.1585,
  -39.1159,
  -39.0642,
  -39.0374,
  -39.0393,
  -39.029,
  -39.0384,
  -39.0375,
  -39.0316,
  -39.0218,
  -39.0112,
  -39.0017,
  -38.9883,
  -38.9941,
  -38.9899,
  -38.9694,
  -38.9542,
  -38.9346,
  -38.9238,
  -38.8764,
  -38.8281,
  -38.8084,
  -38.7928,
  -38.7652,
  -38.7339,
  -38.7097,
  -38.6805,
  -38.6491,
  -38.608,
  -38.5679,
  -38.5241,
  -38.4832,
  -38.4376,
  -38.3961,
  -38.377,
  -38.3554,
  -38.3168,
  -38.3116,
  -38.3251,
  -38.3322,
  -38.358,
  -38.3974,
  -38.435,
  -38.4779,
  -38.5477,
  -38.6429,
  -38.7221,
  -38.8179,
  -38.9439,
  -39.0662,
  -39.1792,
  -39.2935,
  -39.4093,
  -39.5365,
  -39.6699,
  -39.7914,
  -39.9087,
  -40.0263,
  -40.1384,
  -40.2556,
  -40.3731,
  -40.4812,
  -40.5887,
  -40.6969,
  -40.8053,
  -40.9104,
  -41.0115,
  -41.1026,
  -41.1842,
  -41.2544,
  -41.3166,
  -41.3705,
  -41.4202,
  -41.4665,
  -41.5125,
  -41.5608,
  -41.6157,
  -41.6795,
  -41.7411,
  -41.8062,
  -41.8717,
  -41.9412,
  -42.0101,
  -42.0808,
  -42.1533,
  -42.2261,
  -42.299,
  -42.3745,
  -42.4533,
  -42.5357,
  -42.6215,
  -42.7116,
  -42.8075,
  -42.9069,
  -43.0082,
  -43.1095,
  -43.2103,
  -43.3101,
  -43.4092,
  -43.5075,
  -43.6049,
  -43.7016,
  -43.7963,
  -43.8869,
  -43.971,
  -44.0476,
  -44.1151,
  -44.1729,
  -44.2208,
  -44.2593,
  -44.2893,
  -44.3112,
  -44.3253,
  -44.3322,
  -44.3335,
  -44.3292,
  -44.3203,
  -44.3074,
  -44.2906,
  -44.2715,
  -44.2517,
  -44.2334,
  -44.2186,
  -44.2081,
  -44.2016,
  -44.1969,
  -44.1925,
  -44.1844,
  -44.1688,
  -44.1434,
  -44.1066,
  -44.0597,
  -44.0044,
  -43.9431,
  -43.8797,
  -43.8192,
  -43.7657,
  -43.723,
  -43.6941,
  -43.6809,
  -43.6827,
  -43.7,
  -43.732,
  -43.7771,
  -43.8334,
  -43.8993,
  -43.9724,
  -44.0506,
  -44.1301,
  -44.2076,
  -44.2829,
  -44.3532,
  -44.417,
  -44.473,
  -44.5204,
  -44.5578,
  -44.5838,
  -44.5973,
  -44.5973,
  -44.5833,
  -44.556,
  -44.5167,
  -44.4687,
  -44.4155,
  -44.3619,
  -44.3126,
  -44.2703,
  -44.236,
  -44.2084,
  -38.9595,
  -38.9749,
  -38.9871,
  -38.9961,
  -39.0016,
  -39.0041,
  -39.0042,
  -39.002,
  -38.9976,
  -38.9898,
  -38.9817,
  -38.9737,
  -38.9674,
  -38.963,
  -38.961,
  -38.9627,
  -38.9693,
  -38.9817,
  -39.001,
  -39.0277,
  -39.0622,
  -39.105,
  -39.1566,
  -39.2166,
  -39.2884,
  -39.3722,
  -39.4701,
  -39.5843,
  -39.718,
  -39.8724,
  -40.0496,
  -40.2491,
  -40.4695,
  -40.7069,
  -40.9564,
  -41.211,
  -41.4632,
  -41.707,
  -41.9376,
  -42.149,
  -42.3416,
  -42.5126,
  -42.6619,
  -42.7907,
  -42.8997,
  -42.9894,
  -43.0606,
  -43.1139,
  -43.1492,
  -43.1657,
  -43.1639,
  -43.1431,
  -43.103,
  -43.0457,
  -42.97,
  -42.8788,
  -42.7763,
  -42.6642,
  -42.5444,
  -42.4236,
  -42.3022,
  -42.1846,
  -42.0752,
  -41.9783,
  -41.8995,
  -41.8377,
  -41.7947,
  -41.7725,
  -41.7713,
  -41.7815,
  -41.8006,
  -41.8306,
  -41.8676,
  -41.9101,
  -41.954,
  -41.9947,
  -42.0291,
  -42.056,
  -42.0734,
  -42.0827,
  -42.0827,
  -42.0759,
  -42.0633,
  -42.0444,
  -42.0187,
  -41.9851,
  -41.9418,
  -41.8868,
  -41.8185,
  -41.7355,
  -41.6411,
  -41.5374,
  -41.4282,
  -41.3168,
  -41.2067,
  -41.1005,
  -40.9995,
  -40.9052,
  -40.8186,
  -40.7394,
  -40.6662,
  -40.5976,
  -40.5315,
  -40.4664,
  -40.4009,
  -40.3337,
  -40.2647,
  -40.1961,
  -40.1289,
  -40.0662,
  -40.0049,
  -39.9458,
  -39.883,
  -39.8233,
  -39.7735,
  -39.7303,
  -39.6963,
  -39.6659,
  -39.6379,
  -39.6061,
  -39.5816,
  -39.5556,
  -39.5279,
  -39.5011,
  -39.4707,
  -39.4427,
  -39.4237,
  -39.4042,
  -39.3739,
  -39.3496,
  -39.3095,
  -39.2738,
  -39.2546,
  -39.2285,
  -39.1961,
  -39.1705,
  -39.1652,
  -39.1576,
  -39.1522,
  -39.1425,
  -39.1394,
  -39.1318,
  -39.124,
  -39.1144,
  -39.1097,
  -39.1052,
  -39.0952,
  -39.0835,
  -39.0659,
  -39.0425,
  -39.0149,
  -38.9683,
  -38.927,
  -38.8967,
  -38.8826,
  -38.8508,
  -38.8126,
  -38.7871,
  -38.7542,
  -38.708,
  -38.6618,
  -38.6204,
  -38.5787,
  -38.5376,
  -38.5003,
  -38.4841,
  -38.4595,
  -38.4077,
  -38.3656,
  -38.3671,
  -38.3791,
  -38.3733,
  -38.371,
  -38.413,
  -38.4629,
  -38.5188,
  -38.609,
  -38.7064,
  -38.7815,
  -38.8595,
  -38.9618,
  -39.0804,
  -39.2001,
  -39.3253,
  -39.4546,
  -39.5832,
  -39.7156,
  -39.8446,
  -39.9665,
  -40.0898,
  -40.2116,
  -40.3332,
  -40.4524,
  -40.566,
  -40.68,
  -40.7957,
  -40.9114,
  -41.0239,
  -41.1325,
  -41.229,
  -41.3136,
  -41.3866,
  -41.4502,
  -41.5051,
  -41.5563,
  -41.6066,
  -41.6583,
  -41.7133,
  -41.7709,
  -41.8319,
  -41.8974,
  -41.9644,
  -42.0329,
  -42.1064,
  -42.1809,
  -42.2574,
  -42.3359,
  -42.4166,
  -42.4986,
  -42.5843,
  -42.6734,
  -42.7661,
  -42.8613,
  -42.9576,
  -43.0568,
  -43.1586,
  -43.2594,
  -43.3591,
  -43.4567,
  -43.5524,
  -43.6454,
  -43.738,
  -43.8297,
  -43.9208,
  -44.0101,
  -44.0957,
  -44.1757,
  -44.2485,
  -44.313,
  -44.3682,
  -44.4143,
  -44.4517,
  -44.4804,
  -44.5007,
  -44.5128,
  -44.5177,
  -44.5158,
  -44.508,
  -44.4955,
  -44.4779,
  -44.4569,
  -44.4333,
  -44.4085,
  -44.3842,
  -44.3617,
  -44.3419,
  -44.3238,
  -44.3057,
  -44.2857,
  -44.2601,
  -44.2266,
  -44.1826,
  -44.1283,
  -44.0651,
  -43.9954,
  -43.9226,
  -43.8496,
  -43.7833,
  -43.7265,
  -43.6824,
  -43.6531,
  -43.6394,
  -43.6405,
  -43.6561,
  -43.6859,
  -43.728,
  -43.7807,
  -43.844,
  -43.9152,
  -43.9919,
  -44.0711,
  -44.1497,
  -44.2254,
  -44.2961,
  -44.36,
  -44.4161,
  -44.4634,
  -44.5007,
  -44.5273,
  -44.5424,
  -44.5453,
  -44.5356,
  -44.5137,
  -44.4805,
  -44.4384,
  -44.3903,
  -44.34,
  -44.2913,
  -44.2473,
  -44.2094,
  -44.1769,
  -39.0086,
  -39.0261,
  -39.0405,
  -39.0521,
  -39.0595,
  -39.0651,
  -39.0687,
  -39.0698,
  -39.0678,
  -39.0634,
  -39.0578,
  -39.0522,
  -39.0475,
  -39.0437,
  -39.0421,
  -39.0437,
  -39.0493,
  -39.0607,
  -39.0781,
  -39.1038,
  -39.1375,
  -39.1799,
  -39.2307,
  -39.2905,
  -39.3612,
  -39.4431,
  -39.538,
  -39.6493,
  -39.7794,
  -39.9292,
  -40.1009,
  -40.2949,
  -40.5093,
  -40.7414,
  -40.985,
  -41.2356,
  -41.4854,
  -41.7282,
  -41.9588,
  -42.1721,
  -42.3661,
  -42.5388,
  -42.6902,
  -42.8211,
  -42.9318,
  -43.0238,
  -43.0968,
  -43.1513,
  -43.1877,
  -43.2044,
  -43.2043,
  -43.1854,
  -43.1479,
  -43.0938,
  -43.0213,
  -42.9339,
  -42.834,
  -42.724,
  -42.6067,
  -42.4874,
  -42.3687,
  -42.2528,
  -42.1447,
  -42.0481,
  -41.9676,
  -41.9038,
  -41.856,
  -41.8271,
  -41.8174,
  -41.8182,
  -41.8317,
  -41.8563,
  -41.8887,
  -41.926,
  -41.9662,
  -42.0044,
  -42.0384,
  -42.0651,
  -42.0829,
  -42.092,
  -42.0916,
  -42.0832,
  -42.0689,
  -42.0473,
  -42.0205,
  -41.9865,
  -41.944,
  -41.8905,
  -41.8247,
  -41.7455,
  -41.654,
  -41.5528,
  -41.4456,
  -41.334,
  -41.2221,
  -41.1123,
  -41.0065,
  -40.9068,
  -40.8141,
  -40.729,
  -40.6502,
  -40.5768,
  -40.5063,
  -40.4395,
  -40.3731,
  -40.3055,
  -40.2367,
  -40.1676,
  -40.1005,
  -40.0349,
  -39.9745,
  -39.9174,
  -39.8602,
  -39.8067,
  -39.7634,
  -39.7273,
  -39.6962,
  -39.6691,
  -39.6444,
  -39.6193,
  -39.5962,
  -39.5782,
  -39.559,
  -39.5379,
  -39.515,
  -39.4916,
  -39.4837,
  -39.4724,
  -39.455,
  -39.4353,
  -39.4065,
  -39.3841,
  -39.3628,
  -39.3362,
  -39.3118,
  -39.2883,
  -39.2745,
  -39.269,
  -39.2545,
  -39.2443,
  -39.2477,
  -39.2443,
  -39.2389,
  -39.2326,
  -39.2259,
  -39.2226,
  -39.2105,
  -39.1976,
  -39.1774,
  -39.1526,
  -39.1191,
  -39.0792,
  -39.0399,
  -39.0054,
  -38.9788,
  -38.9451,
  -38.9054,
  -38.8709,
  -38.8298,
  -38.7783,
  -38.7243,
  -38.6839,
  -38.6409,
  -38.6183,
  -38.6017,
  -38.5742,
  -38.5391,
  -38.498,
  -38.4753,
  -38.4515,
  -38.4268,
  -38.4302,
  -38.4321,
  -38.477,
  -38.5305,
  -38.5955,
  -38.6863,
  -38.7782,
  -38.8639,
  -38.9322,
  -39.0211,
  -39.1209,
  -39.2442,
  -39.3672,
  -39.4997,
  -39.6403,
  -39.7688,
  -39.8983,
  -40.0281,
  -40.1615,
  -40.2945,
  -40.4254,
  -40.5519,
  -40.6693,
  -40.7903,
  -40.9122,
  -41.034,
  -41.1526,
  -41.2661,
  -41.3675,
  -41.4565,
  -41.5325,
  -41.598,
  -41.6558,
  -41.7086,
  -41.7623,
  -41.8187,
  -41.8776,
  -41.9395,
  -42.0053,
  -42.0729,
  -42.142,
  -42.2139,
  -42.2908,
  -42.369,
  -42.4501,
  -42.5343,
  -42.6222,
  -42.7132,
  -42.807,
  -42.9049,
  -43.0053,
  -43.1064,
  -43.2074,
  -43.3091,
  -43.4103,
  -43.5099,
  -43.6064,
  -43.6997,
  -43.79,
  -43.8781,
  -43.9643,
  -44.0494,
  -44.1342,
  -44.2176,
  -44.2977,
  -44.3724,
  -44.4406,
  -44.5013,
  -44.5533,
  -44.5967,
  -44.6309,
  -44.6567,
  -44.6747,
  -44.6839,
  -44.6856,
  -44.6798,
  -44.6679,
  -44.6504,
  -44.6282,
  -44.602,
  -44.5727,
  -44.5413,
  -44.5086,
  -44.4774,
  -44.447,
  -44.4165,
  -44.3844,
  -44.3488,
  -44.3065,
  -44.2558,
  -44.195,
  -44.1248,
  -44.048,
  -43.9668,
  -43.8851,
  -43.8067,
  -43.7365,
  -43.6775,
  -43.6318,
  -43.6012,
  -43.5852,
  -43.5831,
  -43.5943,
  -43.6192,
  -43.656,
  -43.7039,
  -43.7634,
  -43.8329,
  -43.9089,
  -43.988,
  -44.0679,
  -44.1452,
  -44.2173,
  -44.2824,
  -44.3394,
  -44.3872,
  -44.4248,
  -44.4521,
  -44.4687,
  -44.4743,
  -44.469,
  -44.4519,
  -44.4252,
  -44.3888,
  -44.3457,
  -44.2984,
  -44.2496,
  -44.2039,
  -44.1622,
  -44.125,
  -39.0746,
  -39.0938,
  -39.1101,
  -39.1237,
  -39.1344,
  -39.1423,
  -39.1481,
  -39.1508,
  -39.1503,
  -39.1473,
  -39.1433,
  -39.1395,
  -39.1361,
  -39.1326,
  -39.1311,
  -39.1324,
  -39.1373,
  -39.1482,
  -39.1662,
  -39.192,
  -39.2256,
  -39.2679,
  -39.3193,
  -39.3792,
  -39.4498,
  -39.5312,
  -39.625,
  -39.7351,
  -39.8611,
  -40.0082,
  -40.1762,
  -40.3646,
  -40.5723,
  -40.7968,
  -41.0336,
  -41.2766,
  -41.5197,
  -41.7572,
  -41.9843,
  -42.1959,
  -42.3892,
  -42.562,
  -42.7142,
  -42.847,
  -42.9583,
  -43.051,
  -43.1256,
  -43.1814,
  -43.2194,
  -43.2388,
  -43.2407,
  -43.225,
  -43.1916,
  -43.1416,
  -43.0744,
  -42.9924,
  -42.8982,
  -42.7933,
  -42.6814,
  -42.5673,
  -42.4517,
  -42.34,
  -42.2351,
  -42.1402,
  -42.0589,
  -41.9931,
  -41.941,
  -41.9058,
  -41.8868,
  -41.8794,
  -41.8842,
  -41.9004,
  -41.9246,
  -41.9548,
  -41.9887,
  -42.0228,
  -42.0544,
  -42.0788,
  -42.0962,
  -42.105,
  -42.1039,
  -42.0946,
  -42.0788,
  -42.057,
  -42.0293,
  -41.9956,
  -41.9545,
  -41.9035,
  -41.8406,
  -41.7654,
  -41.6782,
  -41.5809,
  -41.4762,
  -41.3668,
  -41.2543,
  -41.1406,
  -41.0303,
  -40.9248,
  -40.8255,
  -40.7334,
  -40.6481,
  -40.5691,
  -40.4958,
  -40.4266,
  -40.3592,
  -40.2918,
  -40.2237,
  -40.1559,
  -40.0907,
  -40.0287,
  -39.971,
  -39.9155,
  -39.8631,
  -39.8126,
  -39.7716,
  -39.7387,
  -39.7098,
  -39.6869,
  -39.6655,
  -39.6475,
  -39.6311,
  -39.6185,
  -39.6052,
  -39.5945,
  -39.5781,
  -39.5629,
  -39.5528,
  -39.5445,
  -39.5357,
  -39.524,
  -39.5073,
  -39.4864,
  -39.4765,
  -39.4544,
  -39.4381,
  -39.417,
  -39.4009,
  -39.3773,
  -39.3582,
  -39.3572,
  -39.364,
  -39.3659,
  -39.3673,
  -39.3655,
  -39.3584,
  -39.3459,
  -39.3311,
  -39.317,
  -39.2959,
  -39.2652,
  -39.2317,
  -39.1937,
  -39.158,
  -39.1182,
  -39.0815,
  -39.0434,
  -38.9978,
  -38.9557,
  -38.903,
  -38.8456,
  -38.8025,
  -38.7643,
  -38.7302,
  -38.7182,
  -38.7005,
  -38.6756,
  -38.6466,
  -38.6153,
  -38.5815,
  -38.5536,
  -38.5421,
  -38.5339,
  -38.5555,
  -38.6052,
  -38.6483,
  -38.6839,
  -38.7668,
  -38.8475,
  -38.9547,
  -39.0348,
  -39.1106,
  -39.1887,
  -39.3102,
  -39.435,
  -39.551,
  -39.6802,
  -39.81,
  -39.9472,
  -40.0907,
  -40.2505,
  -40.4034,
  -40.5467,
  -40.6791,
  -40.799,
  -40.9237,
  -41.0488,
  -41.1732,
  -41.2944,
  -41.4086,
  -41.5116,
  -41.6025,
  -41.681,
  -41.7487,
  -41.8103,
  -41.8673,
  -41.9242,
  -41.9861,
  -42.0507,
  -42.1183,
  -42.1878,
  -42.2597,
  -42.333,
  -42.4083,
  -42.4873,
  -42.5685,
  -42.653,
  -42.7418,
  -42.8348,
  -42.9322,
  -43.0333,
  -43.1375,
  -43.2428,
  -43.3478,
  -43.4515,
  -43.5537,
  -43.6535,
  -43.7503,
  -43.843,
  -43.9315,
  -44.0165,
  -44.0985,
  -44.1783,
  -44.2571,
  -44.3355,
  -44.4126,
  -44.4869,
  -44.556,
  -44.6193,
  -44.6754,
  -44.7227,
  -44.761,
  -44.7912,
  -44.8131,
  -44.827,
  -44.8315,
  -44.8292,
  -44.8198,
  -44.8033,
  -44.7801,
  -44.7526,
  -44.7207,
  -44.6842,
  -44.6457,
  -44.6054,
  -44.5649,
  -44.5235,
  -44.4807,
  -44.435,
  -44.3842,
  -44.3261,
  -44.2596,
  -44.1836,
  -44.1,
  -44.0118,
  -43.9217,
  -43.8332,
  -43.7504,
  -43.6777,
  -43.6168,
  -43.5689,
  -43.5358,
  -43.5162,
  -43.5096,
  -43.5149,
  -43.5321,
  -43.5625,
  -43.6069,
  -43.6613,
  -43.7282,
  -43.8037,
  -43.8833,
  -43.965,
  -44.0445,
  -44.1184,
  -44.1852,
  -44.2434,
  -44.2919,
  -44.3303,
  -44.3588,
  -44.3771,
  -44.3855,
  -44.3832,
  -44.3715,
  -44.3492,
  -44.3178,
  -44.2783,
  -44.2329,
  -44.1846,
  -44.1368,
  -44.0914,
  -44.0497,
  -39.158,
  -39.1786,
  -39.1963,
  -39.2106,
  -39.2226,
  -39.2322,
  -39.2388,
  -39.2427,
  -39.2421,
  -39.2404,
  -39.2379,
  -39.2353,
  -39.2325,
  -39.2311,
  -39.2303,
  -39.2311,
  -39.2357,
  -39.2464,
  -39.2642,
  -39.2904,
  -39.325,
  -39.3679,
  -39.4199,
  -39.4797,
  -39.5508,
  -39.6324,
  -39.7272,
  -39.8356,
  -39.9621,
  -40.1073,
  -40.2713,
  -40.4546,
  -40.6557,
  -40.8713,
  -41.0977,
  -41.3303,
  -41.5639,
  -41.7933,
  -42.0132,
  -42.2207,
  -42.411,
  -42.5827,
  -42.7348,
  -42.8679,
  -42.9807,
  -43.074,
  -43.1493,
  -43.2064,
  -43.2458,
  -43.2673,
  -43.2717,
  -43.2597,
  -43.2312,
  -43.1868,
  -43.1261,
  -43.0502,
  -42.9633,
  -42.8658,
  -42.761,
  -42.6536,
  -42.5451,
  -42.439,
  -42.3384,
  -42.2457,
  -42.1648,
  -42.0971,
  -42.0414,
  -41.9996,
  -41.9717,
  -41.9555,
  -41.9508,
  -41.9559,
  -41.9708,
  -41.9924,
  -42.0182,
  -42.0468,
  -42.0744,
  -42.0978,
  -42.1141,
  -42.1221,
  -42.1203,
  -42.11,
  -42.093,
  -42.0699,
  -42.042,
  -42.0087,
  -41.9689,
  -41.9204,
  -41.8614,
  -41.7901,
  -41.7082,
  -41.6167,
  -41.5172,
  -41.4109,
  -41.2981,
  -41.1836,
  -41.0693,
  -40.9581,
  -40.8521,
  -40.7533,
  -40.6609,
  -40.5758,
  -40.498,
  -40.4262,
  -40.358,
  -40.2912,
  -40.2244,
  -40.1577,
  -40.093,
  -40.0336,
  -39.9772,
  -39.9245,
  -39.8755,
  -39.8267,
  -39.79,
  -39.7613,
  -39.7395,
  -39.7213,
  -39.7037,
  -39.6901,
  -39.6779,
  -39.6692,
  -39.6606,
  -39.6565,
  -39.6492,
  -39.6405,
  -39.6312,
  -39.6255,
  -39.6143,
  -39.6081,
  -39.6047,
  -39.5955,
  -39.5956,
  -39.588,
  -39.5713,
  -39.5486,
  -39.5317,
  -39.5104,
  -39.4891,
  -39.4802,
  -39.483,
  -39.4934,
  -39.4959,
  -39.4958,
  -39.4911,
  -39.4773,
  -39.4633,
  -39.4423,
  -39.4168,
  -39.3857,
  -39.3517,
  -39.3182,
  -39.2824,
  -39.2435,
  -39.2009,
  -39.1566,
  -39.1065,
  -39.0605,
  -39.0043,
  -38.9516,
  -38.9129,
  -38.8758,
  -38.8487,
  -38.8297,
  -38.807,
  -38.7796,
  -38.7481,
  -38.7183,
  -38.6897,
  -38.6687,
  -38.6631,
  -38.6712,
  -38.6872,
  -38.7337,
  -38.7502,
  -38.797,
  -38.8863,
  -38.97,
  -39.0587,
  -39.143,
  -39.2157,
  -39.2992,
  -39.3946,
  -39.5128,
  -39.6503,
  -39.781,
  -39.9173,
  -40.0478,
  -40.2066,
  -40.3741,
  -40.5347,
  -40.681,
  -40.8153,
  -40.9378,
  -41.0644,
  -41.1909,
  -41.3153,
  -41.4358,
  -41.5493,
  -41.6509,
  -41.7424,
  -41.8223,
  -41.8923,
  -41.9572,
  -42.0188,
  -42.0814,
  -42.1485,
  -42.2193,
  -42.2927,
  -42.3694,
  -42.4476,
  -42.5258,
  -42.6057,
  -42.6884,
  -42.773,
  -42.8608,
  -42.9529,
  -43.0493,
  -43.1501,
  -43.2543,
  -43.3617,
  -43.4693,
  -43.5754,
  -43.6792,
  -43.7806,
  -43.8781,
  -43.9719,
  -44.0606,
  -44.1445,
  -44.2233,
  -44.2998,
  -44.3737,
  -44.4464,
  -44.5188,
  -44.5894,
  -44.6575,
  -44.7212,
  -44.7789,
  -44.8293,
  -44.8718,
  -44.9063,
  -44.9319,
  -44.9481,
  -44.9564,
  -44.956,
  -44.9484,
  -44.9339,
  -44.9123,
  -44.884,
  -44.8501,
  -44.8114,
  -44.7679,
  -44.7212,
  -44.6722,
  -44.6216,
  -44.5695,
  -44.5151,
  -44.4563,
  -44.3916,
  -44.3194,
  -44.239,
  -44.1504,
  -44.0559,
  -43.9583,
  -43.8606,
  -43.7659,
  -43.6793,
  -43.6047,
  -43.5419,
  -43.4922,
  -43.4567,
  -43.433,
  -43.4204,
  -43.4192,
  -43.4294,
  -43.4538,
  -43.4914,
  -43.5438,
  -43.6083,
  -43.6837,
  -43.7647,
  -43.8481,
  -43.9294,
  -44.0053,
  -44.0735,
  -44.1328,
  -44.1823,
  -44.2216,
  -44.251,
  -44.2708,
  -44.2808,
  -44.2814,
  -44.2727,
  -44.2539,
  -44.2251,
  -44.1872,
  -44.1419,
  -44.0921,
  -44.0413,
  -43.9914,
  -43.9455,
  -39.2555,
  -39.2773,
  -39.295,
  -39.3091,
  -39.3213,
  -39.3315,
  -39.3387,
  -39.3429,
  -39.3445,
  -39.3441,
  -39.3429,
  -39.3417,
  -39.3398,
  -39.3386,
  -39.3384,
  -39.3396,
  -39.3444,
  -39.3552,
  -39.3721,
  -39.3986,
  -39.4335,
  -39.4773,
  -39.5299,
  -39.5916,
  -39.6636,
  -39.7459,
  -39.8413,
  -39.9505,
  -40.0762,
  -40.2196,
  -40.3806,
  -40.5587,
  -40.752,
  -40.9573,
  -41.1727,
  -41.3932,
  -41.6154,
  -41.835,
  -42.0478,
  -42.2489,
  -42.4352,
  -42.6042,
  -42.7551,
  -42.8869,
  -42.9993,
  -43.0932,
  -43.1686,
  -43.2262,
  -43.267,
  -43.2896,
  -43.2967,
  -43.2884,
  -43.2646,
  -43.2268,
  -43.1733,
  -43.1066,
  -43.028,
  -42.9395,
  -42.8431,
  -42.7432,
  -42.6427,
  -42.5434,
  -42.4481,
  -42.3591,
  -42.2797,
  -42.21,
  -42.1511,
  -42.1032,
  -42.0676,
  -42.0422,
  -42.0271,
  -42.0226,
  -42.0265,
  -42.0379,
  -42.0557,
  -42.0777,
  -42.0999,
  -42.1194,
  -42.1335,
  -42.1403,
  -42.1382,
  -42.1269,
  -42.1089,
  -42.0839,
  -42.0554,
  -42.0222,
  -41.9839,
  -41.9379,
  -41.8832,
  -41.8184,
  -41.7432,
  -41.6591,
  -41.5648,
  -41.4625,
  -41.3538,
  -41.2387,
  -41.1213,
  -41.0051,
  -40.8928,
  -40.786,
  -40.6866,
  -40.5944,
  -40.5113,
  -40.4367,
  -40.3672,
  -40.3015,
  -40.2364,
  -40.1711,
  -40.1071,
  -40.0475,
  -39.9953,
  -39.9429,
  -39.8903,
  -39.8364,
  -39.8097,
  -39.7892,
  -39.7746,
  -39.7592,
  -39.747,
  -39.7371,
  -39.7289,
  -39.7222,
  -39.7173,
  -39.718,
  -39.7191,
  -39.7172,
  -39.713,
  -39.709,
  -39.6943,
  -39.6946,
  -39.7016,
  -39.7078,
  -39.719,
  -39.7163,
  -39.7053,
  -39.6906,
  -39.6751,
  -39.651,
  -39.6252,
  -39.6095,
  -39.6126,
  -39.6172,
  -39.6222,
  -39.6228,
  -39.6179,
  -39.6063,
  -39.589,
  -39.5638,
  -39.5319,
  -39.4998,
  -39.4679,
  -39.4376,
  -39.4035,
  -39.3668,
  -39.3237,
  -39.2746,
  -39.2256,
  -39.1768,
  -39.1205,
  -39.0744,
  -39.0311,
  -38.9924,
  -38.966,
  -38.9452,
  -38.9161,
  -38.8874,
  -38.8604,
  -38.8368,
  -38.8174,
  -38.8046,
  -38.806,
  -38.8045,
  -38.8334,
  -38.8694,
  -38.9051,
  -38.9454,
  -39.021,
  -39.0977,
  -39.1764,
  -39.2612,
  -39.3397,
  -39.4134,
  -39.5079,
  -39.6051,
  -39.7423,
  -39.892,
  -40.0443,
  -40.2015,
  -40.3683,
  -40.5283,
  -40.6823,
  -40.826,
  -40.9604,
  -41.084,
  -41.2104,
  -41.3349,
  -41.456,
  -41.572,
  -41.6813,
  -41.7811,
  -41.8708,
  -41.9505,
  -42.0225,
  -42.091,
  -42.1574,
  -42.2262,
  -42.2991,
  -42.3766,
  -42.4575,
  -42.5415,
  -42.6265,
  -42.7117,
  -42.7977,
  -42.8846,
  -42.9727,
  -43.0637,
  -43.1579,
  -43.2558,
  -43.3569,
  -43.462,
  -43.5692,
  -43.6756,
  -43.7808,
  -43.8829,
  -43.9814,
  -44.0764,
  -44.1663,
  -44.2509,
  -44.3313,
  -44.4066,
  -44.4781,
  -44.5469,
  -44.6141,
  -44.6807,
  -44.7453,
  -44.8074,
  -44.865,
  -44.9164,
  -44.9613,
  -44.9985,
  -45.0267,
  -45.0457,
  -45.0562,
  -45.0584,
  -45.0526,
  -45.0396,
  -45.0193,
  -44.9921,
  -44.9583,
  -44.9177,
  -44.8719,
  -44.8208,
  -44.7645,
  -44.7071,
  -44.6469,
  -44.5849,
  -44.5193,
  -44.4489,
  -44.3723,
  -44.2882,
  -44.1963,
  -44.0972,
  -43.9935,
  -43.8883,
  -43.7847,
  -43.6867,
  -43.5966,
  -43.5193,
  -43.4547,
  -43.4037,
  -43.3645,
  -43.3366,
  -43.319,
  -43.3122,
  -43.3169,
  -43.3354,
  -43.3687,
  -43.4179,
  -43.4814,
  -43.556,
  -43.6376,
  -43.7217,
  -43.8042,
  -43.8812,
  -43.9505,
  -44.0104,
  -44.06,
  -44.0997,
  -44.1295,
  -44.1496,
  -44.1602,
  -44.1617,
  -44.154,
  -44.1362,
  -44.108,
  -44.0685,
  -44.0216,
  -43.9694,
  -43.9142,
  -43.8602,
  -43.8105,
  -39.362,
  -39.3833,
  -39.4018,
  -39.4169,
  -39.4298,
  -39.4399,
  -39.4476,
  -39.4525,
  -39.4551,
  -39.4563,
  -39.4571,
  -39.4572,
  -39.4571,
  -39.4557,
  -39.456,
  -39.4578,
  -39.4635,
  -39.4745,
  -39.4925,
  -39.5189,
  -39.5538,
  -39.5976,
  -39.6505,
  -39.7129,
  -39.7857,
  -39.8694,
  -39.9654,
  -40.075,
  -40.1989,
  -40.3402,
  -40.4977,
  -40.6697,
  -40.8554,
  -41.0518,
  -41.2556,
  -41.4643,
  -41.6746,
  -41.8836,
  -42.0874,
  -42.2813,
  -42.4621,
  -42.6273,
  -42.7753,
  -42.9042,
  -43.0154,
  -43.1084,
  -43.1835,
  -43.2414,
  -43.2831,
  -43.3086,
  -43.3185,
  -43.3135,
  -43.295,
  -43.2628,
  -43.2171,
  -43.1587,
  -43.0889,
  -43.0092,
  -42.9221,
  -42.8309,
  -42.7375,
  -42.6452,
  -42.556,
  -42.4715,
  -42.3945,
  -42.3255,
  -42.2645,
  -42.2123,
  -42.1699,
  -42.136,
  -42.1109,
  -42.0951,
  -42.0893,
  -42.0901,
  -42.0987,
  -42.1123,
  -42.1278,
  -42.1416,
  -42.1526,
  -42.1578,
  -42.1548,
  -42.1436,
  -42.1248,
  -42.1003,
  -42.0711,
  -42.0376,
  -41.9999,
  -41.9562,
  -41.9057,
  -41.8467,
  -41.7791,
  -41.7023,
  -41.616,
  -41.5195,
  -41.4145,
  -41.3004,
  -41.1822,
  -41.0628,
  -40.9445,
  -40.8311,
  -40.7244,
  -40.6267,
  -40.5382,
  -40.4602,
  -40.3897,
  -40.3246,
  -40.2621,
  -40.1994,
  -40.1385,
  -40.0823,
  -40.0315,
  -39.9773,
  -39.9296,
  -39.8881,
  -39.8628,
  -39.8439,
  -39.8266,
  -39.8129,
  -39.806,
  -39.7987,
  -39.794,
  -39.7884,
  -39.7863,
  -39.7882,
  -39.7908,
  -39.8015,
  -39.8039,
  -39.7946,
  -39.7901,
  -39.798,
  -39.8135,
  -39.8323,
  -39.845,
  -39.8494,
  -39.8437,
  -39.8309,
  -39.8159,
  -39.7954,
  -39.7709,
  -39.7557,
  -39.7541,
  -39.7535,
  -39.7507,
  -39.7477,
  -39.74,
  -39.728,
  -39.7085,
  -39.6819,
  -39.6481,
  -39.6148,
  -39.5821,
  -39.5504,
  -39.5154,
  -39.4792,
  -39.4363,
  -39.3899,
  -39.3409,
  -39.2937,
  -39.239,
  -39.1929,
  -39.1506,
  -39.114,
  -39.0816,
  -39.0584,
  -39.0292,
  -39.0004,
  -38.9767,
  -38.9589,
  -38.9494,
  -38.9445,
  -38.9475,
  -38.9559,
  -38.9797,
  -39.01,
  -39.0507,
  -39.1046,
  -39.1657,
  -39.2355,
  -39.3101,
  -39.3897,
  -39.4694,
  -39.5512,
  -39.6501,
  -39.7445,
  -39.8737,
  -40.0188,
  -40.1896,
  -40.3529,
  -40.5239,
  -40.6844,
  -40.8347,
  -40.9762,
  -41.1104,
  -41.2332,
  -41.357,
  -41.4768,
  -41.5916,
  -41.7006,
  -41.8021,
  -41.8964,
  -41.982,
  -42.0598,
  -42.1322,
  -42.2045,
  -42.276,
  -42.3513,
  -42.4312,
  -42.5157,
  -42.6034,
  -42.6963,
  -42.7893,
  -42.8813,
  -42.9742,
  -43.0661,
  -43.1584,
  -43.2529,
  -43.3486,
  -43.4466,
  -43.5482,
  -43.6516,
  -43.7557,
  -43.8588,
  -43.9605,
  -44.0584,
  -44.1539,
  -44.2456,
  -44.332,
  -44.413,
  -44.4892,
  -44.5609,
  -44.6288,
  -44.6928,
  -44.7548,
  -44.8157,
  -44.8744,
  -44.9304,
  -44.9815,
  -45.0269,
  -45.0655,
  -45.0951,
  -45.117,
  -45.1292,
  -45.1335,
  -45.1295,
  -45.117,
  -45.0991,
  -45.073,
  -45.0396,
  -44.9999,
  -44.9525,
  -44.8999,
  -44.8408,
  -44.7769,
  -44.7115,
  -44.6431,
  -44.5717,
  -44.4964,
  -44.4161,
  -44.3299,
  -44.2365,
  -44.1358,
  -44.0285,
  -43.9178,
  -43.8063,
  -43.6975,
  -43.5952,
  -43.5026,
  -43.4227,
  -43.3563,
  -43.3031,
  -43.2618,
  -43.2307,
  -43.2093,
  -43.1983,
  -43.199,
  -43.2138,
  -43.2444,
  -43.2915,
  -43.3535,
  -43.4266,
  -43.5075,
  -43.5912,
  -43.6735,
  -43.7501,
  -43.8189,
  -43.878,
  -43.9266,
  -43.9654,
  -43.9945,
  -44.0136,
  -44.0232,
  -44.0236,
  -44.0147,
  -43.9956,
  -43.9652,
  -43.9242,
  -43.8738,
  -43.817,
  -43.7576,
  -43.6998,
  -43.6468,
  -39.4751,
  -39.4962,
  -39.5143,
  -39.53,
  -39.5431,
  -39.5539,
  -39.5624,
  -39.5686,
  -39.5724,
  -39.5755,
  -39.5784,
  -39.5803,
  -39.5821,
  -39.5837,
  -39.5851,
  -39.5881,
  -39.5943,
  -39.6059,
  -39.6241,
  -39.6501,
  -39.6845,
  -39.7276,
  -39.7802,
  -39.842,
  -39.9152,
  -39.9995,
  -40.096,
  -40.2053,
  -40.3289,
  -40.4674,
  -40.6202,
  -40.7862,
  -40.9639,
  -41.1507,
  -41.3439,
  -41.5412,
  -41.7404,
  -41.9385,
  -42.1314,
  -42.3175,
  -42.4918,
  -42.652,
  -42.7962,
  -42.9231,
  -43.0322,
  -43.1236,
  -43.1979,
  -43.2557,
  -43.2979,
  -43.325,
  -43.3373,
  -43.3356,
  -43.3212,
  -43.2947,
  -43.2545,
  -43.2039,
  -43.1427,
  -43.0721,
  -42.9936,
  -42.911,
  -42.8265,
  -42.7413,
  -42.6584,
  -42.5788,
  -42.5049,
  -42.437,
  -42.3754,
  -42.3208,
  -42.2729,
  -42.232,
  -42.1982,
  -42.173,
  -42.1559,
  -42.1467,
  -42.1451,
  -42.1495,
  -42.1577,
  -42.1664,
  -42.1733,
  -42.1761,
  -42.1723,
  -42.1608,
  -42.1425,
  -42.118,
  -42.0879,
  -42.0539,
  -42.0161,
  -41.9747,
  -41.9285,
  -41.8744,
  -41.8137,
  -41.7451,
  -41.6672,
  -41.5786,
  -41.4788,
  -41.3698,
  -41.2526,
  -41.1314,
  -41.0096,
  -40.8905,
  -40.7774,
  -40.6734,
  -40.5794,
  -40.4977,
  -40.426,
  -40.3617,
  -40.3017,
  -40.2429,
  -40.1888,
  -40.1385,
  -40.0898,
  -40.0401,
  -40.0002,
  -39.9654,
  -39.9408,
  -39.9274,
  -39.914,
  -39.9025,
  -39.8954,
  -39.8917,
  -39.8885,
  -39.8842,
  -39.8763,
  -39.8768,
  -39.8893,
  -39.9005,
  -39.9034,
  -39.9002,
  -39.9087,
  -39.9238,
  -39.9426,
  -39.9644,
  -39.9814,
  -39.9905,
  -39.9863,
  -39.9755,
  -39.9601,
  -39.9409,
  -39.9229,
  -39.9083,
  -39.8962,
  -39.8872,
  -39.8801,
  -39.8721,
  -39.8619,
  -39.8474,
  -39.8272,
  -39.8,
  -39.7669,
  -39.7311,
  -39.6957,
  -39.6607,
  -39.6233,
  -39.5841,
  -39.5398,
  -39.4951,
  -39.4496,
  -39.405,
  -39.353,
  -39.3079,
  -39.2652,
  -39.2284,
  -39.1964,
  -39.173,
  -39.1419,
  -39.114,
  -39.0909,
  -39.0771,
  -39.0729,
  -39.0716,
  -39.0785,
  -39.0936,
  -39.1171,
  -39.1487,
  -39.1957,
  -39.2503,
  -39.3122,
  -39.3809,
  -39.4549,
  -39.5344,
  -39.6199,
  -39.7109,
  -39.8139,
  -39.9264,
  -40.055,
  -40.1955,
  -40.3524,
  -40.5147,
  -40.6803,
  -40.836,
  -40.9845,
  -41.125,
  -41.2574,
  -41.3777,
  -41.4965,
  -41.6092,
  -41.7152,
  -41.8144,
  -41.9052,
  -41.9908,
  -42.0704,
  -42.1454,
  -42.2187,
  -42.2938,
  -42.3708,
  -42.4532,
  -42.5409,
  -42.6344,
  -42.7316,
  -42.8317,
  -42.9318,
  -43.0323,
  -43.133,
  -43.2298,
  -43.3271,
  -43.4238,
  -43.5214,
  -43.6188,
  -43.7174,
  -43.817,
  -43.9165,
  -44.0137,
  -44.1095,
  -44.203,
  -44.2939,
  -44.3811,
  -44.4639,
  -44.5414,
  -44.6131,
  -44.6816,
  -44.7455,
  -44.8061,
  -44.8636,
  -44.9184,
  -44.9708,
  -45.0203,
  -45.0651,
  -45.1039,
  -45.1359,
  -45.1604,
  -45.1755,
  -45.1814,
  -45.1787,
  -45.1686,
  -45.1504,
  -45.1255,
  -45.0949,
  -45.0559,
  -45.0093,
  -44.955,
  -44.8945,
  -44.8286,
  -44.7586,
  -44.6848,
  -44.6083,
  -44.5289,
  -44.4458,
  -44.3577,
  -44.2641,
  -44.1641,
  -44.0572,
  -43.9447,
  -43.8289,
  -43.7119,
  -43.5972,
  -43.4904,
  -43.3947,
  -43.3124,
  -43.2441,
  -43.1896,
  -43.1467,
  -43.1145,
  -43.0915,
  -43.0796,
  -43.0783,
  -43.092,
  -43.1218,
  -43.1684,
  -43.2287,
  -43.3009,
  -43.3805,
  -43.4627,
  -43.5431,
  -43.6174,
  -43.6835,
  -43.7399,
  -43.786,
  -43.8219,
  -43.8484,
  -43.8652,
  -43.8722,
  -43.8699,
  -43.8578,
  -43.8353,
  -43.8005,
  -43.7546,
  -43.6995,
  -43.6376,
  -43.5737,
  -43.5122,
  -43.4574,
  -39.5908,
  -39.6114,
  -39.6295,
  -39.6447,
  -39.6585,
  -39.6705,
  -39.6808,
  -39.6893,
  -39.6964,
  -39.7023,
  -39.7077,
  -39.7124,
  -39.7165,
  -39.7201,
  -39.7236,
  -39.7281,
  -39.7354,
  -39.7474,
  -39.7647,
  -39.7902,
  -39.8235,
  -39.8658,
  -39.9178,
  -39.98,
  -40.0531,
  -40.1372,
  -40.2331,
  -40.3416,
  -40.463,
  -40.5975,
  -40.7456,
  -40.9058,
  -41.0756,
  -41.2518,
  -41.4351,
  -41.6219,
  -41.8105,
  -41.9982,
  -42.1825,
  -42.3601,
  -42.5273,
  -42.6816,
  -42.8208,
  -42.9439,
  -43.0499,
  -43.1391,
  -43.212,
  -43.2694,
  -43.3116,
  -43.3389,
  -43.3532,
  -43.3543,
  -43.3436,
  -43.3214,
  -43.2886,
  -43.2446,
  -43.1911,
  -43.1285,
  -43.0583,
  -42.9833,
  -42.9062,
  -42.8286,
  -42.7516,
  -42.6776,
  -42.6082,
  -42.5417,
  -42.4808,
  -42.4249,
  -42.3738,
  -42.3275,
  -42.288,
  -42.2549,
  -42.2287,
  -42.2095,
  -42.1978,
  -42.1922,
  -42.1914,
  -42.193,
  -42.1949,
  -42.195,
  -42.1901,
  -42.1789,
  -42.16,
  -42.1359,
  -42.1062,
  -42.0721,
  -42.0347,
  -41.9944,
  -41.9516,
  -41.9038,
  -41.8501,
  -41.7897,
  -41.7206,
  -41.6405,
  -41.5485,
  -41.445,
  -41.3314,
  -41.211,
  -41.0873,
  -40.9647,
  -40.8472,
  -40.7365,
  -40.638,
  -40.5527,
  -40.4787,
  -40.4143,
  -40.3568,
  -40.304,
  -40.2549,
  -40.2096,
  -40.1679,
  -40.1267,
  -40.0915,
  -40.0623,
  -40.0417,
  -40.0285,
  -40.0184,
  -40.0113,
  -40.0077,
  -40.0061,
  -40.0036,
  -40.0014,
  -39.9965,
  -39.9998,
  -40.0083,
  -40.0192,
  -40.032,
  -40.0462,
  -40.0608,
  -40.0788,
  -40.0994,
  -40.1201,
  -40.1354,
  -40.1427,
  -40.1398,
  -40.1297,
  -40.114,
  -40.0953,
  -40.0783,
  -40.0596,
  -40.042,
  -40.0257,
  -40.0134,
  -40.0008,
  -39.9865,
  -39.9697,
  -39.948,
  -39.921,
  -39.8873,
  -39.8523,
  -39.8149,
  -39.7754,
  -39.7337,
  -39.6923,
  -39.6479,
  -39.6028,
  -39.5584,
  -39.517,
  -39.4699,
  -39.4264,
  -39.3861,
  -39.3488,
  -39.3161,
  -39.2897,
  -39.2585,
  -39.2311,
  -39.2079,
  -39.1941,
  -39.1911,
  -39.1927,
  -39.2032,
  -39.223,
  -39.2527,
  -39.2903,
  -39.3429,
  -39.4033,
  -39.4689,
  -39.5389,
  -39.6148,
  -39.6964,
  -39.784,
  -39.8781,
  -39.9819,
  -40.0983,
  -40.2254,
  -40.3652,
  -40.5133,
  -40.6664,
  -40.8226,
  -40.9731,
  -41.1187,
  -41.2567,
  -41.3861,
  -41.5043,
  -41.6167,
  -41.7214,
  -41.8175,
  -41.9059,
  -41.9873,
  -42.0638,
  -42.1369,
  -42.209,
  -42.2832,
  -42.3619,
  -42.4458,
  -42.5365,
  -42.6339,
  -42.7371,
  -42.8434,
  -42.9515,
  -43.0587,
  -43.1664,
  -43.273,
  -43.3766,
  -43.4767,
  -43.5757,
  -43.6726,
  -43.7673,
  -43.8616,
  -43.9547,
  -44.0472,
  -44.1377,
  -44.2261,
  -44.3129,
  -44.3975,
  -44.4797,
  -44.5585,
  -44.6327,
  -44.7021,
  -44.7672,
  -44.8278,
  -44.8847,
  -44.9378,
  -44.9871,
  -45.0335,
  -45.0758,
  -45.1145,
  -45.1472,
  -45.1724,
  -45.1901,
  -45.1986,
  -45.1987,
  -45.1899,
  -45.1733,
  -45.1498,
  -45.1191,
  -45.082,
  -45.0363,
  -44.984,
  -44.9233,
  -44.8558,
  -44.7818,
  -44.7042,
  -44.6226,
  -44.5391,
  -44.453,
  -44.3635,
  -44.2699,
  -44.1711,
  -44.0673,
  -43.9571,
  -43.842,
  -43.7234,
  -43.6024,
  -43.4843,
  -43.3738,
  -43.2748,
  -43.1901,
  -43.1197,
  -43.0645,
  -43.0218,
  -42.9892,
  -42.9673,
  -42.9566,
  -42.9582,
  -42.9731,
  -43.0042,
  -43.051,
  -43.1114,
  -43.181,
  -43.258,
  -43.3371,
  -43.4141,
  -43.4839,
  -43.5451,
  -43.5966,
  -43.6377,
  -43.6688,
  -43.6909,
  -43.7032,
  -43.7061,
  -43.6995,
  -43.6829,
  -43.6556,
  -43.6145,
  -43.5633,
  -43.5025,
  -43.4358,
  -43.3677,
  -43.3037,
  -43.249,
  -39.7055,
  -39.7259,
  -39.7446,
  -39.7613,
  -39.7763,
  -39.7904,
  -39.8028,
  -39.814,
  -39.8242,
  -39.8336,
  -39.8421,
  -39.8501,
  -39.8571,
  -39.8622,
  -39.8683,
  -39.8744,
  -39.8834,
  -39.8964,
  -39.9152,
  -39.94,
  -39.9723,
  -40.0135,
  -40.0641,
  -40.1255,
  -40.1974,
  -40.2807,
  -40.3752,
  -40.4815,
  -40.599,
  -40.73,
  -40.8727,
  -41.0261,
  -41.1881,
  -41.3564,
  -41.5302,
  -41.7075,
  -41.8859,
  -42.0638,
  -42.2387,
  -42.4076,
  -42.5672,
  -42.7147,
  -42.8485,
  -42.9658,
  -43.0683,
  -43.1548,
  -43.226,
  -43.2825,
  -43.3247,
  -43.3536,
  -43.3693,
  -43.3726,
  -43.365,
  -43.347,
  -43.3189,
  -43.2808,
  -43.2338,
  -43.1782,
  -43.1153,
  -43.0465,
  -42.9763,
  -42.9053,
  -42.8347,
  -42.7669,
  -42.702,
  -42.6407,
  -42.5821,
  -42.5264,
  -42.4744,
  -42.4253,
  -42.3803,
  -42.3401,
  -42.3057,
  -42.2772,
  -42.2552,
  -42.2392,
  -42.228,
  -42.2216,
  -42.2178,
  -42.2146,
  -42.2087,
  -42.198,
  -42.1813,
  -42.1583,
  -42.1298,
  -42.0963,
  -42.0594,
  -42.0205,
  -41.9794,
  -41.9363,
  -41.8903,
  -41.8372,
  -41.7768,
  -41.7062,
  -41.622,
  -41.5258,
  -41.4184,
  -41.3014,
  -41.1786,
  -41.0554,
  -40.9354,
  -40.8226,
  -40.7201,
  -40.6311,
  -40.5546,
  -40.4892,
  -40.4325,
  -40.382,
  -40.3375,
  -40.2965,
  -40.2597,
  -40.2259,
  -40.1962,
  -40.1695,
  -40.1522,
  -40.1402,
  -40.1331,
  -40.1298,
  -40.1292,
  -40.1308,
  -40.1334,
  -40.1361,
  -40.1382,
  -40.1447,
  -40.1523,
  -40.1671,
  -40.1826,
  -40.2005,
  -40.2192,
  -40.2407,
  -40.2639,
  -40.2844,
  -40.2994,
  -40.306,
  -40.3035,
  -40.294,
  -40.2779,
  -40.2575,
  -40.2375,
  -40.215,
  -40.1923,
  -40.1713,
  -40.1531,
  -40.1344,
  -40.1159,
  -40.0955,
  -40.0717,
  -40.0438,
  -40.0094,
  -39.9732,
  -39.9339,
  -39.8921,
  -39.8481,
  -39.8041,
  -39.7574,
  -39.7117,
  -39.667,
  -39.6249,
  -39.5795,
  -39.5386,
  -39.5006,
  -39.4652,
  -39.4338,
  -39.4072,
  -39.3792,
  -39.3533,
  -39.3327,
  -39.3192,
  -39.3173,
  -39.3212,
  -39.3351,
  -39.3598,
  -39.3957,
  -39.4401,
  -39.4972,
  -39.562,
  -39.6321,
  -39.706,
  -39.7837,
  -39.8665,
  -39.9536,
  -40.0487,
  -40.1523,
  -40.2663,
  -40.3904,
  -40.5248,
  -40.6674,
  -40.8153,
  -40.9661,
  -41.1134,
  -41.2545,
  -41.3876,
  -41.5111,
  -41.6229,
  -41.7261,
  -41.8192,
  -41.9033,
  -41.979,
  -42.0486,
  -42.115,
  -42.1816,
  -42.2516,
  -42.3275,
  -42.4124,
  -42.5049,
  -42.6053,
  -42.7126,
  -42.8242,
  -42.9391,
  -43.054,
  -43.1694,
  -43.2829,
  -43.394,
  -43.5007,
  -43.6034,
  -43.702,
  -43.7975,
  -43.8894,
  -43.978,
  -44.0637,
  -44.1468,
  -44.2281,
  -44.3083,
  -44.3873,
  -44.4651,
  -44.5414,
  -44.6155,
  -44.6862,
  -44.7525,
  -44.8142,
  -44.8712,
  -44.9241,
  -44.9728,
  -45.0168,
  -45.0573,
  -45.093,
  -45.1245,
  -45.1514,
  -45.1708,
  -45.181,
  -45.1835,
  -45.1777,
  -45.1634,
  -45.1411,
  -45.1117,
  -45.0752,
  -45.0313,
  -44.9797,
  -44.9206,
  -44.8537,
  -44.779,
  -44.6994,
  -44.6156,
  -44.5283,
  -44.4388,
  -44.3471,
  -44.2529,
  -44.1558,
  -44.0543,
  -43.9484,
  -43.8378,
  -43.7207,
  -43.601,
  -43.4775,
  -43.3569,
  -43.2428,
  -43.1406,
  -43.0523,
  -42.9802,
  -42.9234,
  -42.8816,
  -42.8522,
  -42.8336,
  -42.8272,
  -42.834,
  -42.8542,
  -42.889,
  -42.9358,
  -42.9956,
  -43.0648,
  -43.1387,
  -43.2133,
  -43.2847,
  -43.3487,
  -43.4032,
  -43.4475,
  -43.4816,
  -43.5064,
  -43.522,
  -43.5287,
  -43.5265,
  -43.5148,
  -43.4931,
  -43.4602,
  -43.4147,
  -43.3581,
  -43.2923,
  -43.2218,
  -43.1513,
  -43.0871,
  -43.0333,
  -39.8211,
  -39.8416,
  -39.8609,
  -39.8784,
  -39.8947,
  -39.9107,
  -39.9256,
  -39.9401,
  -39.9526,
  -39.9655,
  -39.9779,
  -39.9894,
  -39.9995,
  -40.0092,
  -40.0176,
  -40.0267,
  -40.0382,
  -40.0525,
  -40.0724,
  -40.0969,
  -40.1287,
  -40.1688,
  -40.217,
  -40.2766,
  -40.3471,
  -40.4286,
  -40.5212,
  -40.6248,
  -40.7398,
  -40.8661,
  -41.0032,
  -41.1494,
  -41.3036,
  -41.4637,
  -41.6283,
  -41.7962,
  -41.9651,
  -42.1336,
  -42.2983,
  -42.4585,
  -42.61,
  -42.75,
  -42.8778,
  -42.9909,
  -43.0895,
  -43.1731,
  -43.2425,
  -43.2978,
  -43.3395,
  -43.3687,
  -43.3854,
  -43.3904,
  -43.3851,
  -43.3704,
  -43.3454,
  -43.3119,
  -43.2705,
  -43.2212,
  -43.165,
  -43.1041,
  -43.0404,
  -42.9759,
  -42.9119,
  -42.8497,
  -42.7905,
  -42.7335,
  -42.6784,
  -42.625,
  -42.5732,
  -42.5229,
  -42.4734,
  -42.4277,
  -42.3858,
  -42.3484,
  -42.3162,
  -42.2903,
  -42.2703,
  -42.2559,
  -42.2464,
  -42.2395,
  -42.2325,
  -42.2228,
  -42.2077,
  -42.1871,
  -42.1607,
  -42.1291,
  -42.0935,
  -42.0561,
  -42.0163,
  -41.9769,
  -41.9354,
  -41.89,
  -41.8379,
  -41.7765,
  -41.7029,
  -41.6168,
  -41.5171,
  -41.4067,
  -41.2884,
  -41.1674,
  -41.0477,
  -40.9338,
  -40.8291,
  -40.7368,
  -40.6571,
  -40.5897,
  -40.5326,
  -40.4823,
  -40.4394,
  -40.402,
  -40.3694,
  -40.3402,
  -40.3155,
  -40.2941,
  -40.2797,
  -40.2708,
  -40.2668,
  -40.267,
  -40.2698,
  -40.275,
  -40.281,
  -40.2872,
  -40.2936,
  -40.3043,
  -40.3156,
  -40.3295,
  -40.3464,
  -40.3655,
  -40.3866,
  -40.4105,
  -40.4341,
  -40.4549,
  -40.4703,
  -40.4776,
  -40.4772,
  -40.4683,
  -40.452,
  -40.4303,
  -40.4078,
  -40.3811,
  -40.3542,
  -40.3284,
  -40.3041,
  -40.2805,
  -40.2569,
  -40.232,
  -40.2044,
  -40.1732,
  -40.1347,
  -40.0964,
  -40.0555,
  -40.0123,
  -39.9667,
  -39.9213,
  -39.8736,
  -39.8262,
  -39.7815,
  -39.7397,
  -39.6959,
  -39.6576,
  -39.6225,
  -39.5892,
  -39.5593,
  -39.533,
  -39.5064,
  -39.4821,
  -39.4621,
  -39.4489,
  -39.4477,
  -39.453,
  -39.4695,
  -39.497,
  -39.538,
  -39.5883,
  -39.6507,
  -39.7206,
  -39.7954,
  -39.8735,
  -39.9539,
  -40.0377,
  -40.1253,
  -40.2183,
  -40.3184,
  -40.4275,
  -40.5458,
  -40.6741,
  -40.8104,
  -40.9525,
  -41.0973,
  -41.2389,
  -41.3746,
  -41.5016,
  -41.6175,
  -41.7203,
  -41.813,
  -41.8944,
  -41.9652,
  -42.0271,
  -42.0853,
  -42.143,
  -42.2048,
  -42.2747,
  -42.3552,
  -42.4478,
  -42.551,
  -42.6629,
  -42.7807,
  -42.9026,
  -43.0258,
  -43.1481,
  -43.2681,
  -43.3852,
  -43.4985,
  -43.6068,
  -43.7094,
  -43.8059,
  -43.8969,
  -43.983,
  -44.064,
  -44.1406,
  -44.2132,
  -44.2836,
  -44.3537,
  -44.4239,
  -44.4944,
  -44.5645,
  -44.6329,
  -44.698,
  -44.7611,
  -44.8199,
  -44.8733,
  -44.9219,
  -44.9659,
  -45.005,
  -45.0394,
  -45.0691,
  -45.0942,
  -45.1143,
  -45.1279,
  -45.1333,
  -45.13,
  -45.1184,
  -45.099,
  -45.0712,
  -45.0363,
  -44.9936,
  -44.9433,
  -44.8851,
  -44.8195,
  -44.7458,
  -44.6647,
  -44.5781,
  -44.488,
  -44.3953,
  -44.3008,
  -44.2047,
  -44.1073,
  -44.008,
  -43.906,
  -43.8006,
  -43.6893,
  -43.5734,
  -43.4534,
  -43.3291,
  -43.2075,
  -43.0905,
  -42.9859,
  -42.8968,
  -42.8233,
  -42.766,
  -42.7255,
  -42.6998,
  -42.6885,
  -42.6904,
  -42.7046,
  -42.7321,
  -42.7723,
  -42.8236,
  -42.8846,
  -42.9524,
  -43.0232,
  -43.0928,
  -43.1573,
  -43.2138,
  -43.2604,
  -43.2962,
  -43.3216,
  -43.3382,
  -43.3459,
  -43.3458,
  -43.3376,
  -43.3204,
  -43.2933,
  -43.2549,
  -43.2052,
  -43.1447,
  -43.0764,
  -43.0044,
  -42.9345,
  -42.8718,
  -42.8211,
  -39.9367,
  -39.9574,
  -39.9768,
  -39.9941,
  -40.0121,
  -40.0298,
  -40.0474,
  -40.0648,
  -40.0816,
  -40.098,
  -40.114,
  -40.1288,
  -40.1427,
  -40.1554,
  -40.1679,
  -40.1805,
  -40.1947,
  -40.2113,
  -40.2319,
  -40.2566,
  -40.2887,
  -40.3278,
  -40.3761,
  -40.4342,
  -40.5032,
  -40.5827,
  -40.6726,
  -40.7731,
  -40.8839,
  -41.005,
  -41.1358,
  -41.2749,
  -41.42,
  -41.5718,
  -41.7279,
  -41.8866,
  -42.0465,
  -42.2055,
  -42.3621,
  -42.5133,
  -42.6564,
  -42.7894,
  -42.9104,
  -43.0183,
  -43.1126,
  -43.1934,
  -43.2604,
  -43.3142,
  -43.3541,
  -43.3829,
  -43.4004,
  -43.4066,
  -43.4032,
  -43.3907,
  -43.3699,
  -43.3409,
  -43.3046,
  -43.2611,
  -43.2113,
  -43.1571,
  -43.0998,
  -43.042,
  -42.9846,
  -42.9285,
  -42.8747,
  -42.8215,
  -42.7706,
  -42.7202,
  -42.6697,
  -42.6192,
  -42.5692,
  -42.5191,
  -42.4703,
  -42.4248,
  -42.3837,
  -42.3483,
  -42.3196,
  -42.2976,
  -42.2822,
  -42.2722,
  -42.2643,
  -42.2551,
  -42.2418,
  -42.2242,
  -42.2011,
  -42.172,
  -42.1387,
  -42.103,
  -42.0662,
  -42.0297,
  -41.9922,
  -41.9532,
  -41.9099,
  -41.8577,
  -41.794,
  -41.7176,
  -41.6281,
  -41.5262,
  -41.4158,
  -41.3001,
  -41.1826,
  -41.0701,
  -40.9647,
  -40.8701,
  -40.7878,
  -40.7177,
  -40.6587,
  -40.609,
  -40.5673,
  -40.5316,
  -40.5011,
  -40.4752,
  -40.4539,
  -40.4366,
  -40.4257,
  -40.4202,
  -40.4193,
  -40.4225,
  -40.4283,
  -40.4365,
  -40.4446,
  -40.4539,
  -40.4634,
  -40.4762,
  -40.4885,
  -40.503,
  -40.5203,
  -40.5408,
  -40.5626,
  -40.5871,
  -40.6113,
  -40.6327,
  -40.6489,
  -40.6574,
  -40.6581,
  -40.6501,
  -40.6342,
  -40.6117,
  -40.5873,
  -40.5576,
  -40.5268,
  -40.4951,
  -40.4652,
  -40.4362,
  -40.4072,
  -40.3774,
  -40.3453,
  -40.3093,
  -40.2683,
  -40.2275,
  -40.1865,
  -40.142,
  -40.0949,
  -40.0486,
  -40.0005,
  -39.9534,
  -39.9085,
  -39.8667,
  -39.8229,
  -39.787,
  -39.7541,
  -39.7238,
  -39.6954,
  -39.6695,
  -39.6436,
  -39.6198,
  -39.5997,
  -39.586,
  -39.5845,
  -39.5903,
  -39.6083,
  -39.6396,
  -39.6842,
  -39.7391,
  -39.8062,
  -39.8809,
  -39.9599,
  -40.0415,
  -40.1236,
  -40.207,
  -40.2922,
  -40.3808,
  -40.4749,
  -40.5765,
  -40.6868,
  -40.807,
  -40.9356,
  -41.0704,
  -41.2076,
  -41.3433,
  -41.472,
  -41.5916,
  -41.699,
  -41.7928,
  -41.874,
  -41.9428,
  -42.0009,
  -42.0519,
  -42.1,
  -42.1518,
  -42.2119,
  -42.2849,
  -42.3728,
  -42.4758,
  -42.5913,
  -42.7154,
  -42.8444,
  -42.9751,
  -43.1053,
  -43.2323,
  -43.3554,
  -43.4738,
  -43.587,
  -43.6938,
  -43.793,
  -43.8855,
  -43.9696,
  -44.0457,
  -44.1162,
  -44.1821,
  -44.2433,
  -44.3019,
  -44.3609,
  -44.4214,
  -44.4837,
  -44.5471,
  -44.61,
  -44.6712,
  -44.7302,
  -44.7853,
  -44.835,
  -44.8794,
  -44.9183,
  -44.952,
  -44.9807,
  -45.0044,
  -45.0232,
  -45.0367,
  -45.0444,
  -45.0441,
  -45.0351,
  -45.0181,
  -44.9929,
  -44.9601,
  -44.92,
  -44.8704,
  -44.8133,
  -44.7486,
  -44.6762,
  -44.5954,
  -44.506,
  -44.4133,
  -44.3168,
  -44.2188,
  -44.1207,
  -44.021,
  -43.9216,
  -43.8217,
  -43.7203,
  -43.6159,
  -43.5066,
  -43.3929,
  -43.2744,
  -43.1525,
  -43.0313,
  -42.9161,
  -42.8112,
  -42.7214,
  -42.6493,
  -42.5944,
  -42.5571,
  -42.5372,
  -42.5338,
  -42.5457,
  -42.5708,
  -42.608,
  -42.656,
  -42.7127,
  -42.7757,
  -42.8429,
  -42.9102,
  -42.974,
  -43.0313,
  -43.0794,
  -43.1168,
  -43.143,
  -43.159,
  -43.1662,
  -43.1657,
  -43.1579,
  -43.1429,
  -43.1199,
  -43.0869,
  -43.0446,
  -42.9922,
  -42.9304,
  -42.8625,
  -42.7926,
  -42.7257,
  -42.6669,
  -42.6207,
  -40.0506,
  -40.0714,
  -40.0911,
  -40.11,
  -40.1292,
  -40.1483,
  -40.1684,
  -40.188,
  -40.2078,
  -40.2273,
  -40.246,
  -40.2644,
  -40.2815,
  -40.2985,
  -40.315,
  -40.3316,
  -40.3495,
  -40.3695,
  -40.3921,
  -40.4187,
  -40.4512,
  -40.4907,
  -40.5383,
  -40.5954,
  -40.6625,
  -40.7397,
  -40.8271,
  -40.923,
  -41.0294,
  -41.145,
  -41.2694,
  -41.4012,
  -41.5396,
  -41.6831,
  -41.8303,
  -41.9802,
  -42.1309,
  -42.2808,
  -42.428,
  -42.5703,
  -42.7053,
  -42.8306,
  -42.9448,
  -43.0464,
  -43.1365,
  -43.2138,
  -43.2783,
  -43.3304,
  -43.37,
  -43.3982,
  -43.4158,
  -43.4229,
  -43.4207,
  -43.4102,
  -43.3927,
  -43.3676,
  -43.336,
  -43.2983,
  -43.255,
  -43.2064,
  -43.1562,
  -43.105,
  -43.054,
  -43.0041,
  -42.9554,
  -42.9079,
  -42.8612,
  -42.8141,
  -42.7662,
  -42.7164,
  -42.6647,
  -42.612,
  -42.5585,
  -42.5063,
  -42.4575,
  -42.414,
  -42.3771,
  -42.349,
  -42.3287,
  -42.3156,
  -42.3063,
  -42.2978,
  -42.2878,
  -42.2741,
  -42.2549,
  -42.2294,
  -42.1992,
  -42.1652,
  -42.1307,
  -42.0963,
  -42.0629,
  -42.0291,
  -41.9923,
  -41.9484,
  -41.894,
  -41.8281,
  -41.7496,
  -41.6591,
  -41.5582,
  -41.4508,
  -41.3402,
  -41.2308,
  -41.1273,
  -41.032,
  -40.9473,
  -40.8751,
  -40.8137,
  -40.7629,
  -40.7203,
  -40.6852,
  -40.6559,
  -40.6319,
  -40.613,
  -40.5974,
  -40.5891,
  -40.5862,
  -40.5881,
  -40.5937,
  -40.6017,
  -40.6123,
  -40.6237,
  -40.6352,
  -40.6467,
  -40.66,
  -40.6728,
  -40.6872,
  -40.704,
  -40.7236,
  -40.7447,
  -40.7686,
  -40.7926,
  -40.8142,
  -40.8311,
  -40.8398,
  -40.8419,
  -40.8353,
  -40.8203,
  -40.798,
  -40.7724,
  -40.7406,
  -40.7064,
  -40.6717,
  -40.6371,
  -40.6026,
  -40.5685,
  -40.534,
  -40.4976,
  -40.4581,
  -40.4145,
  -40.372,
  -40.3295,
  -40.2837,
  -40.2361,
  -40.1894,
  -40.1418,
  -40.0944,
  -40.0504,
  -40.0093,
  -39.968,
  -39.9339,
  -39.9027,
  -39.8739,
  -39.8465,
  -39.8215,
  -39.7958,
  -39.7717,
  -39.751,
  -39.7363,
  -39.7332,
  -39.7383,
  -39.7565,
  -39.7889,
  -39.8354,
  -39.8932,
  -39.9631,
  -40.0405,
  -40.1219,
  -40.2047,
  -40.2865,
  -40.3663,
  -40.4466,
  -40.5282,
  -40.6135,
  -40.7054,
  -40.8058,
  -40.9161,
  -41.0356,
  -41.162,
  -41.2922,
  -41.421,
  -41.5439,
  -41.6572,
  -41.7559,
  -41.8409,
  -41.9105,
  -41.9673,
  -42.0136,
  -42.0549,
  -42.0958,
  -42.1452,
  -42.2068,
  -42.2865,
  -42.3847,
  -42.4999,
  -42.6283,
  -42.7648,
  -42.9038,
  -43.0421,
  -43.1771,
  -43.3066,
  -43.4303,
  -43.5467,
  -43.6567,
  -43.7586,
  -43.8521,
  -43.9362,
  -44.0107,
  -44.0777,
  -44.1362,
  -44.1892,
  -44.238,
  -44.2848,
  -44.3325,
  -44.3827,
  -44.4364,
  -44.4927,
  -44.5498,
  -44.6061,
  -44.6604,
  -44.711,
  -44.7567,
  -44.7966,
  -44.8305,
  -44.8583,
  -44.8805,
  -44.8979,
  -44.911,
  -44.9169,
  -44.9168,
  -44.9106,
  -44.8964,
  -44.8743,
  -44.8434,
  -44.8057,
  -44.7599,
  -44.7036,
  -44.6389,
  -44.5681,
  -44.4869,
  -44.3985,
  -44.3028,
  -44.2032,
  -44.1016,
  -43.9986,
  -43.8965,
  -43.7953,
  -43.6953,
  -43.5966,
  -43.4963,
  -43.394,
  -43.2876,
  -43.1774,
  -43.0622,
  -42.9435,
  -42.8269,
  -42.7154,
  -42.6143,
  -42.5277,
  -42.4587,
  -42.4087,
  -42.3781,
  -42.3666,
  -42.3735,
  -42.3967,
  -42.4343,
  -42.4832,
  -42.5402,
  -42.6033,
  -42.6691,
  -42.7359,
  -42.7999,
  -42.8578,
  -42.9071,
  -42.9462,
  -42.9741,
  -42.9906,
  -42.997,
  -42.9947,
  -42.985,
  -42.9692,
  -42.9468,
  -42.9182,
  -42.8823,
  -42.8374,
  -42.7848,
  -42.7247,
  -42.6604,
  -42.5955,
  -42.5346,
  -42.4822,
  -42.4412,
  -40.1639,
  -40.1847,
  -40.2046,
  -40.2241,
  -40.2438,
  -40.2642,
  -40.2855,
  -40.3061,
  -40.3279,
  -40.3498,
  -40.3713,
  -40.393,
  -40.4143,
  -40.4353,
  -40.4565,
  -40.478,
  -40.5002,
  -40.524,
  -40.5497,
  -40.5786,
  -40.6125,
  -40.6529,
  -40.6996,
  -40.7561,
  -40.822,
  -40.8969,
  -40.9812,
  -41.0745,
  -41.1764,
  -41.2866,
  -41.4046,
  -41.5295,
  -41.6601,
  -41.7954,
  -41.9339,
  -42.0746,
  -42.2161,
  -42.3558,
  -42.4939,
  -42.6276,
  -42.7545,
  -42.8724,
  -42.9801,
  -43.0769,
  -43.1622,
  -43.2357,
  -43.2973,
  -43.3473,
  -43.3857,
  -43.413,
  -43.43,
  -43.4373,
  -43.4362,
  -43.4268,
  -43.412,
  -43.3912,
  -43.3645,
  -43.3328,
  -43.2962,
  -43.2557,
  -43.2124,
  -43.1678,
  -43.1234,
  -43.0788,
  -43.0349,
  -42.992,
  -42.949,
  -42.9053,
  -42.8596,
  -42.8109,
  -42.7588,
  -42.7042,
  -42.6474,
  -42.591,
  -42.5369,
  -42.4878,
  -42.4465,
  -42.4141,
  -42.3902,
  -42.374,
  -42.3632,
  -42.355,
  -42.347,
  -42.3367,
  -42.3216,
  -42.3006,
  -42.2732,
  -42.2428,
  -42.2087,
  -42.1768,
  -42.146,
  -42.1164,
  -42.0851,
  -42.0487,
  -42.0039,
  -41.9487,
  -41.8819,
  -41.8032,
  -41.7138,
  -41.616,
  -41.5133,
  -41.4103,
  -41.3104,
  -41.2166,
  -41.1315,
  -41.0568,
  -40.993,
  -40.9402,
  -40.8966,
  -40.8608,
  -40.8315,
  -40.8087,
  -40.7909,
  -40.7778,
  -40.7707,
  -40.7691,
  -40.7725,
  -40.7797,
  -40.7895,
  -40.8012,
  -40.8139,
  -40.8267,
  -40.8389,
  -40.8516,
  -40.8637,
  -40.8769,
  -40.891,
  -40.9086,
  -40.9281,
  -40.9501,
  -40.9727,
  -40.9939,
  -41.0112,
  -41.0222,
  -41.0257,
  -41.0207,
  -41.0069,
  -40.9851,
  -40.9581,
  -40.9248,
  -40.8883,
  -40.8503,
  -40.8119,
  -40.7734,
  -40.7352,
  -40.6969,
  -40.658,
  -40.6174,
  -40.5724,
  -40.5289,
  -40.4853,
  -40.4395,
  -40.3924,
  -40.3459,
  -40.2994,
  -40.2547,
  -40.2125,
  -40.1734,
  -40.1358,
  -40.1033,
  -40.0735,
  -40.0456,
  -40.0184,
  -39.9925,
  -39.9659,
  -39.9404,
  -39.918,
  -39.901,
  -39.894,
  -39.8969,
  -39.9134,
  -39.9436,
  -39.9896,
  -40.0481,
  -40.1182,
  -40.1956,
  -40.2765,
  -40.3577,
  -40.4364,
  -40.5121,
  -40.5851,
  -40.6573,
  -40.7319,
  -40.8123,
  -40.9011,
  -41,
  -41.1091,
  -41.2268,
  -41.3497,
  -41.4724,
  -41.5893,
  -41.6954,
  -41.7877,
  -41.8636,
  -41.9236,
  -41.9702,
  -42.0072,
  -42.0402,
  -42.077,
  -42.1263,
  -42.1942,
  -42.2834,
  -42.3943,
  -42.5228,
  -42.6639,
  -42.8118,
  -42.9601,
  -43.1046,
  -43.2417,
  -43.3708,
  -43.491,
  -43.6036,
  -43.707,
  -43.8001,
  -43.8844,
  -43.9574,
  -44.0214,
  -44.0753,
  -44.1216,
  -44.1611,
  -44.1974,
  -44.2325,
  -44.2692,
  -44.3097,
  -44.3545,
  -44.4036,
  -44.4538,
  -44.505,
  -44.5544,
  -44.5999,
  -44.6405,
  -44.6753,
  -44.7035,
  -44.7252,
  -44.7407,
  -44.7508,
  -44.756,
  -44.7552,
  -44.748,
  -44.7352,
  -44.7151,
  -44.6868,
  -44.6524,
  -44.6085,
  -44.555,
  -44.4928,
  -44.4222,
  -44.3419,
  -44.254,
  -44.1582,
  -44.0563,
  -43.9499,
  -43.8425,
  -43.7368,
  -43.6315,
  -43.5296,
  -43.4303,
  -43.333,
  -43.2351,
  -43.1356,
  -43.0333,
  -42.9267,
  -42.8158,
  -42.7031,
  -42.5941,
  -42.4905,
  -42.3964,
  -42.3172,
  -42.2562,
  -42.2147,
  -42.1939,
  -42.1933,
  -42.2126,
  -42.2497,
  -42.3008,
  -42.3622,
  -42.4306,
  -42.5008,
  -42.5705,
  -42.6365,
  -42.6967,
  -42.7485,
  -42.7898,
  -42.82,
  -42.8386,
  -42.8457,
  -42.8426,
  -42.8306,
  -42.812,
  -42.7881,
  -42.7589,
  -42.725,
  -42.6854,
  -42.6402,
  -42.5885,
  -42.5324,
  -42.4744,
  -42.4173,
  -42.3645,
  -42.319,
  -42.2853,
  -40.2737,
  -40.2946,
  -40.3134,
  -40.3331,
  -40.353,
  -40.3742,
  -40.3961,
  -40.4188,
  -40.4423,
  -40.4656,
  -40.4896,
  -40.5142,
  -40.539,
  -40.5641,
  -40.5901,
  -40.6165,
  -40.6436,
  -40.6706,
  -40.7002,
  -40.7325,
  -40.769,
  -40.8108,
  -40.8595,
  -40.9158,
  -40.9804,
  -41.0535,
  -41.1352,
  -41.2249,
  -41.3225,
  -41.4277,
  -41.5398,
  -41.6578,
  -41.7798,
  -41.9069,
  -42.0366,
  -42.1682,
  -42.3007,
  -42.4322,
  -42.5615,
  -42.6864,
  -42.8053,
  -42.9159,
  -43.0168,
  -43.1075,
  -43.1875,
  -43.257,
  -43.3153,
  -43.3629,
  -43.3986,
  -43.4246,
  -43.441,
  -43.4488,
  -43.4487,
  -43.4425,
  -43.4307,
  -43.4139,
  -43.3929,
  -43.3671,
  -43.3377,
  -43.3045,
  -43.2684,
  -43.2304,
  -43.1915,
  -43.152,
  -43.1114,
  -43.0721,
  -43.0322,
  -42.9913,
  -42.9478,
  -42.9008,
  -42.8501,
  -42.7953,
  -42.7379,
  -42.6795,
  -42.6232,
  -42.5715,
  -42.5274,
  -42.4924,
  -42.4659,
  -42.4472,
  -42.4349,
  -42.4264,
  -42.4184,
  -42.4105,
  -42.3989,
  -42.382,
  -42.3589,
  -42.3308,
  -42.3012,
  -42.2714,
  -42.2429,
  -42.2164,
  -42.1891,
  -42.1589,
  -42.1222,
  -42.0761,
  -42.0201,
  -41.9531,
  -41.8751,
  -41.7879,
  -41.6937,
  -41.5977,
  -41.5032,
  -41.413,
  -41.3288,
  -41.2543,
  -41.1904,
  -41.1364,
  -41.0918,
  -41.0556,
  -41.0258,
  -41.0025,
  -40.9845,
  -40.9716,
  -40.9646,
  -40.9632,
  -40.9666,
  -40.9743,
  -40.9846,
  -40.9959,
  -41.0093,
  -41.0225,
  -41.035,
  -41.0469,
  -41.0581,
  -41.0695,
  -41.0822,
  -41.0972,
  -41.114,
  -41.1333,
  -41.1538,
  -41.1739,
  -41.1914,
  -41.2035,
  -41.209,
  -41.2064,
  -41.1949,
  -41.1751,
  -41.1488,
  -41.1158,
  -41.0775,
  -41.0378,
  -40.9972,
  -40.9561,
  -40.9151,
  -40.8743,
  -40.8334,
  -40.7921,
  -40.7483,
  -40.7045,
  -40.6596,
  -40.614,
  -40.5678,
  -40.5218,
  -40.4764,
  -40.4327,
  -40.3917,
  -40.3538,
  -40.3178,
  -40.2859,
  -40.2563,
  -40.2282,
  -40.2007,
  -40.1724,
  -40.1445,
  -40.1175,
  -40.0933,
  -40.0745,
  -40.0646,
  -40.0651,
  -40.079,
  -40.1078,
  -40.1511,
  -40.2072,
  -40.2744,
  -40.3484,
  -40.4252,
  -40.501,
  -40.5732,
  -40.6405,
  -40.7036,
  -40.7643,
  -40.826,
  -40.893,
  -40.9685,
  -41.0548,
  -41.1527,
  -41.2608,
  -41.3746,
  -41.4906,
  -41.6023,
  -41.7035,
  -41.7906,
  -41.861,
  -41.9152,
  -41.9553,
  -41.9868,
  -42.0169,
  -42.0542,
  -42.1082,
  -42.1836,
  -42.2838,
  -42.4072,
  -42.5483,
  -42.7006,
  -42.857,
  -43.011,
  -43.1585,
  -43.295,
  -43.4203,
  -43.5345,
  -43.6377,
  -43.7315,
  -43.8144,
  -43.8857,
  -43.9465,
  -43.9965,
  -44.0381,
  -44.0714,
  -44.0989,
  -44.1232,
  -44.1475,
  -44.1748,
  -44.2061,
  -44.2428,
  -44.2845,
  -44.3296,
  -44.3759,
  -44.4195,
  -44.4594,
  -44.4938,
  -44.5223,
  -44.5443,
  -44.5587,
  -44.5663,
  -44.5671,
  -44.563,
  -44.5542,
  -44.539,
  -44.5188,
  -44.4921,
  -44.459,
  -44.4175,
  -44.3679,
  -44.3078,
  -44.239,
  -44.1591,
  -44.0713,
  -43.9754,
  -43.8711,
  -43.7633,
  -43.6517,
  -43.5398,
  -43.432,
  -43.3254,
  -43.2236,
  -43.1264,
  -43.0321,
  -42.9382,
  -42.8427,
  -42.7459,
  -42.6455,
  -42.5447,
  -42.4407,
  -42.3417,
  -42.2496,
  -42.1679,
  -42.1002,
  -42.0518,
  -42.024,
  -42.0168,
  -42.0316,
  -42.0655,
  -42.1182,
  -42.1827,
  -42.2564,
  -42.3341,
  -42.4102,
  -42.4825,
  -42.5476,
  -42.6036,
  -42.6489,
  -42.6826,
  -42.7044,
  -42.7142,
  -42.7125,
  -42.7007,
  -42.6801,
  -42.6529,
  -42.6209,
  -42.5851,
  -42.5448,
  -42.5022,
  -42.4561,
  -42.4071,
  -42.3564,
  -42.3059,
  -42.2575,
  -42.2139,
  -42.1771,
  -42.1503,
  -40.3773,
  -40.3982,
  -40.4176,
  -40.4369,
  -40.457,
  -40.4781,
  -40.5002,
  -40.5234,
  -40.5473,
  -40.5724,
  -40.5984,
  -40.6256,
  -40.653,
  -40.6822,
  -40.7125,
  -40.7436,
  -40.7759,
  -40.8086,
  -40.8427,
  -40.8788,
  -40.9185,
  -40.9629,
  -41.0129,
  -41.0696,
  -41.1339,
  -41.2056,
  -41.2849,
  -41.3709,
  -41.4649,
  -41.5654,
  -41.6718,
  -41.7834,
  -41.8992,
  -42.0182,
  -42.1394,
  -42.2621,
  -42.3855,
  -42.5079,
  -42.6283,
  -42.7448,
  -42.8555,
  -42.9585,
  -43.0515,
  -43.1359,
  -43.2106,
  -43.2755,
  -43.3303,
  -43.3751,
  -43.41,
  -43.4348,
  -43.4508,
  -43.4592,
  -43.4604,
  -43.4562,
  -43.4475,
  -43.4351,
  -43.4191,
  -43.3999,
  -43.3776,
  -43.3507,
  -43.3214,
  -43.2895,
  -43.2556,
  -43.2206,
  -43.1847,
  -43.1482,
  -43.1109,
  -43.072,
  -43.0304,
  -42.9853,
  -42.936,
  -42.8828,
  -42.8265,
  -42.7692,
  -42.7134,
  -42.6619,
  -42.6163,
  -42.5803,
  -42.5524,
  -42.5319,
  -42.5182,
  -42.5089,
  -42.5019,
  -42.4954,
  -42.4863,
  -42.4727,
  -42.4531,
  -42.4287,
  -42.4019,
  -42.3747,
  -42.3488,
  -42.3244,
  -42.3006,
  -42.2749,
  -42.2432,
  -42.2055,
  -42.1589,
  -42.1021,
  -42.0347,
  -41.9579,
  -41.8743,
  -41.7867,
  -41.6987,
  -41.6131,
  -41.532,
  -41.4591,
  -41.3953,
  -41.3407,
  -41.2955,
  -41.2585,
  -41.2282,
  -41.2037,
  -41.185,
  -41.1703,
  -41.1626,
  -41.1604,
  -41.1633,
  -41.1703,
  -41.1806,
  -41.193,
  -41.2066,
  -41.2198,
  -41.2318,
  -41.2428,
  -41.2525,
  -41.2619,
  -41.272,
  -41.2835,
  -41.2971,
  -41.3134,
  -41.3316,
  -41.3501,
  -41.3672,
  -41.3794,
  -41.3869,
  -41.387,
  -41.3785,
  -41.3614,
  -41.337,
  -41.3055,
  -41.2689,
  -41.2292,
  -41.1878,
  -41.146,
  -41.1043,
  -41.063,
  -41.0219,
  -40.9804,
  -40.9378,
  -40.8948,
  -40.8508,
  -40.8059,
  -40.7604,
  -40.7153,
  -40.6707,
  -40.6268,
  -40.5863,
  -40.5485,
  -40.5132,
  -40.481,
  -40.4506,
  -40.4213,
  -40.3921,
  -40.3628,
  -40.3331,
  -40.3042,
  -40.2778,
  -40.2566,
  -40.2436,
  -40.2409,
  -40.2514,
  -40.2761,
  -40.315,
  -40.3662,
  -40.4276,
  -40.495,
  -40.5645,
  -40.6321,
  -40.6947,
  -40.7505,
  -40.8015,
  -40.8491,
  -40.8972,
  -40.95,
  -41.0118,
  -41.0851,
  -41.1715,
  -41.2698,
  -41.3767,
  -41.4868,
  -41.5941,
  -41.6923,
  -41.7767,
  -41.8445,
  -41.8958,
  -41.9334,
  -41.9633,
  -41.9939,
  -42.0346,
  -42.0944,
  -42.179,
  -42.2899,
  -42.4235,
  -42.5746,
  -42.735,
  -42.8969,
  -43.0521,
  -43.1977,
  -43.3302,
  -43.4485,
  -43.5535,
  -43.646,
  -43.727,
  -43.7962,
  -43.8544,
  -43.9023,
  -43.9404,
  -43.9694,
  -43.9918,
  -44.0088,
  -44.0236,
  -44.0388,
  -44.0572,
  -44.0811,
  -44.111,
  -44.1466,
  -44.1854,
  -44.2249,
  -44.2627,
  -44.2958,
  -44.3232,
  -44.3437,
  -44.3563,
  -44.3618,
  -44.36,
  -44.3522,
  -44.3383,
  -44.3188,
  -44.2956,
  -44.2673,
  -44.2341,
  -44.1943,
  -44.1467,
  -44.0897,
  -44.0225,
  -43.9456,
  -43.8581,
  -43.7629,
  -43.6587,
  -43.5499,
  -43.4374,
  -43.3227,
  -43.2082,
  -43.1002,
  -42.9939,
  -42.8938,
  -42.7995,
  -42.7095,
  -42.6209,
  -42.5318,
  -42.4428,
  -42.3519,
  -42.2595,
  -42.1681,
  -42.083,
  -42.006,
  -41.9405,
  -41.8901,
  -41.8591,
  -41.8482,
  -41.8592,
  -41.8912,
  -41.9425,
  -42.0103,
  -42.0884,
  -42.1717,
  -42.2563,
  -42.3369,
  -42.4098,
  -42.4726,
  -42.5235,
  -42.5622,
  -42.5885,
  -42.6028,
  -42.6047,
  -42.5952,
  -42.5755,
  -42.547,
  -42.5114,
  -42.4714,
  -42.4285,
  -42.3837,
  -42.3375,
  -42.2908,
  -42.2443,
  -42.199,
  -42.1559,
  -42.1166,
  -42.082,
  -42.0538,
  -42.0338,
  -40.4753,
  -40.4956,
  -40.5143,
  -40.5328,
  -40.5526,
  -40.5736,
  -40.5956,
  -40.618,
  -40.6425,
  -40.6689,
  -40.697,
  -40.7267,
  -40.7579,
  -40.791,
  -40.8257,
  -40.861,
  -40.8981,
  -40.9357,
  -40.9743,
  -41.0146,
  -41.0579,
  -41.1051,
  -41.1563,
  -41.2143,
  -41.2788,
  -41.3499,
  -41.4279,
  -41.5124,
  -41.6033,
  -41.6998,
  -41.8011,
  -41.9068,
  -42.0157,
  -42.1273,
  -42.2405,
  -42.3545,
  -42.4693,
  -42.5819,
  -42.6932,
  -42.8009,
  -42.9034,
  -42.9986,
  -43.0852,
  -43.1633,
  -43.2325,
  -43.2927,
  -43.344,
  -43.3859,
  -43.4188,
  -43.4427,
  -43.4584,
  -43.4672,
  -43.4698,
  -43.4665,
  -43.4606,
  -43.4523,
  -43.4416,
  -43.4284,
  -43.413,
  -43.3942,
  -43.3713,
  -43.3448,
  -43.3155,
  -43.2842,
  -43.251,
  -43.217,
  -43.1818,
  -43.1446,
  -43.1048,
  -43.0617,
  -43.0138,
  -42.9632,
  -42.9103,
  -42.8562,
  -42.8037,
  -42.755,
  -42.7118,
  -42.6765,
  -42.6486,
  -42.627,
  -42.6116,
  -42.6008,
  -42.593,
  -42.5865,
  -42.579,
  -42.568,
  -42.5523,
  -42.5311,
  -42.5079,
  -42.4836,
  -42.4595,
  -42.4366,
  -42.4149,
  -42.3921,
  -42.3659,
  -42.3343,
  -42.2952,
  -42.247,
  -42.1887,
  -42.1215,
  -42.0471,
  -41.9679,
  -41.8871,
  -41.8072,
  -41.7308,
  -41.6602,
  -41.5965,
  -41.5423,
  -41.4967,
  -41.4591,
  -41.4279,
  -41.4025,
  -41.3823,
  -41.3678,
  -41.3589,
  -41.3556,
  -41.3576,
  -41.364,
  -41.3741,
  -41.3865,
  -41.4,
  -41.4132,
  -41.4249,
  -41.4351,
  -41.4437,
  -41.451,
  -41.4573,
  -41.4656,
  -41.4761,
  -41.489,
  -41.5045,
  -41.5211,
  -41.5378,
  -41.552,
  -41.5615,
  -41.5643,
  -41.559,
  -41.5453,
  -41.5235,
  -41.4944,
  -41.4598,
  -41.4217,
  -41.3815,
  -41.3409,
  -41.3003,
  -41.2604,
  -41.2206,
  -41.18,
  -41.1395,
  -41.0984,
  -41.0559,
  -41.0121,
  -40.9673,
  -40.9226,
  -40.8784,
  -40.8353,
  -40.7944,
  -40.7559,
  -40.7198,
  -40.6859,
  -40.6535,
  -40.6219,
  -40.5903,
  -40.5583,
  -40.5262,
  -40.4948,
  -40.466,
  -40.4421,
  -40.4259,
  -40.4198,
  -40.425,
  -40.4448,
  -40.4777,
  -40.522,
  -40.5754,
  -40.6339,
  -40.6936,
  -40.7507,
  -40.8021,
  -40.8465,
  -40.8847,
  -40.919,
  -40.9534,
  -40.9924,
  -41.0406,
  -41.1015,
  -41.1765,
  -41.2655,
  -41.3647,
  -41.4695,
  -41.5737,
  -41.6699,
  -41.7536,
  -41.8213,
  -41.8728,
  -41.9112,
  -41.9415,
  -41.9751,
  -42.0215,
  -42.0886,
  -42.1819,
  -42.3017,
  -42.4427,
  -42.6003,
  -42.7643,
  -42.9265,
  -43.0802,
  -43.2209,
  -43.3463,
  -43.4554,
  -43.5486,
  -43.6279,
  -43.6942,
  -43.7493,
  -43.7936,
  -43.8284,
  -43.8546,
  -43.8736,
  -43.8872,
  -43.8963,
  -43.9039,
  -43.9126,
  -43.9248,
  -43.9428,
  -43.9665,
  -43.9961,
  -44.0273,
  -44.0601,
  -44.0909,
  -44.1165,
  -44.1358,
  -44.1468,
  -44.1493,
  -44.1447,
  -44.1323,
  -44.1137,
  -44.0899,
  -44.0619,
  -44.0299,
  -43.9938,
  -43.9536,
  -43.9071,
  -43.8526,
  -43.7877,
  -43.7127,
  -43.6273,
  -43.5326,
  -43.43,
  -43.32,
  -43.2073,
  -43.0927,
  -42.9769,
  -42.8621,
  -42.7557,
  -42.6508,
  -42.5536,
  -42.4644,
  -42.3798,
  -42.2982,
  -42.2176,
  -42.1384,
  -42.056,
  -41.9777,
  -41.8987,
  -41.8303,
  -41.7721,
  -41.7265,
  -41.6966,
  -41.6862,
  -41.6968,
  -41.729,
  -41.7814,
  -41.8505,
  -41.9331,
  -42.0228,
  -42.1151,
  -42.2041,
  -42.2863,
  -42.3577,
  -42.4163,
  -42.4615,
  -42.4935,
  -42.513,
  -42.5204,
  -42.5157,
  -42.4999,
  -42.4733,
  -42.437,
  -42.3938,
  -42.3451,
  -42.2943,
  -42.2427,
  -42.1918,
  -42.1434,
  -42.0981,
  -42.0572,
  -42.021,
  -41.9894,
  -41.9632,
  -41.9425,
  -41.929,
  -40.5645,
  -40.5846,
  -40.6019,
  -40.6201,
  -40.6393,
  -40.6596,
  -40.6814,
  -40.7049,
  -40.7298,
  -40.7573,
  -40.7868,
  -40.8184,
  -40.8526,
  -40.8893,
  -40.9274,
  -40.9672,
  -41.0083,
  -41.0489,
  -41.0918,
  -41.1362,
  -41.1832,
  -41.2336,
  -41.2887,
  -41.3488,
  -41.4146,
  -41.4863,
  -41.5634,
  -41.6465,
  -41.7348,
  -41.8277,
  -41.9244,
  -42.0245,
  -42.1261,
  -42.2309,
  -42.3367,
  -42.4431,
  -42.549,
  -42.6542,
  -42.7568,
  -42.8558,
  -42.9497,
  -43.0369,
  -43.1163,
  -43.1881,
  -43.2517,
  -43.3075,
  -43.3551,
  -43.3943,
  -43.4244,
  -43.4476,
  -43.4632,
  -43.4729,
  -43.4773,
  -43.4772,
  -43.474,
  -43.4691,
  -43.4629,
  -43.4554,
  -43.4453,
  -43.4321,
  -43.4145,
  -43.3924,
  -43.3668,
  -43.3383,
  -43.3067,
  -43.2748,
  -43.2415,
  -43.2061,
  -43.1682,
  -43.1273,
  -43.0836,
  -43.0372,
  -42.9885,
  -42.9395,
  -42.8918,
  -42.8472,
  -42.8073,
  -42.7737,
  -42.7462,
  -42.7245,
  -42.7079,
  -42.695,
  -42.6862,
  -42.6792,
  -42.6722,
  -42.6629,
  -42.6504,
  -42.6338,
  -42.6139,
  -42.5925,
  -42.5709,
  -42.5498,
  -42.5296,
  -42.5088,
  -42.4861,
  -42.4589,
  -42.4249,
  -42.3831,
  -42.3328,
  -42.2723,
  -42.2057,
  -42.1339,
  -42.06,
  -41.9861,
  -41.9142,
  -41.8468,
  -41.7859,
  -41.7325,
  -41.6869,
  -41.6485,
  -41.6166,
  -41.5904,
  -41.5696,
  -41.5543,
  -41.5446,
  -41.5408,
  -41.5422,
  -41.5486,
  -41.5588,
  -41.5708,
  -41.585,
  -41.5987,
  -41.6109,
  -41.6209,
  -41.6288,
  -41.6349,
  -41.6401,
  -41.6457,
  -41.653,
  -41.6629,
  -41.6758,
  -41.6908,
  -41.7068,
  -41.7216,
  -41.7328,
  -41.7384,
  -41.7361,
  -41.7256,
  -41.707,
  -41.6811,
  -41.6483,
  -41.6129,
  -41.5754,
  -41.5374,
  -41.4996,
  -41.4627,
  -41.4261,
  -41.3895,
  -41.352,
  -41.3133,
  -41.2728,
  -41.2303,
  -41.1861,
  -41.1411,
  -41.096,
  -41.0522,
  -41.0096,
  -40.9692,
  -40.931,
  -40.8946,
  -40.8595,
  -40.8246,
  -40.7889,
  -40.7536,
  -40.7185,
  -40.6844,
  -40.653,
  -40.6265,
  -40.6072,
  -40.5975,
  -40.5994,
  -40.6136,
  -40.6396,
  -40.6761,
  -40.7201,
  -40.7684,
  -40.8173,
  -40.8628,
  -40.9024,
  -40.9346,
  -40.9605,
  -40.9825,
  -41.0044,
  -41.031,
  -41.0671,
  -41.1165,
  -41.181,
  -41.2597,
  -41.3518,
  -41.4519,
  -41.5528,
  -41.6481,
  -41.7322,
  -41.8013,
  -41.855,
  -41.8962,
  -41.9316,
  -41.9702,
  -42.0223,
  -42.0958,
  -42.1947,
  -42.3193,
  -42.4643,
  -42.6229,
  -42.7849,
  -42.9431,
  -43.0905,
  -43.2231,
  -43.3382,
  -43.4354,
  -43.5156,
  -43.5804,
  -43.6325,
  -43.6737,
  -43.7057,
  -43.7289,
  -43.7465,
  -43.7577,
  -43.7653,
  -43.77,
  -43.7735,
  -43.7779,
  -43.7862,
  -43.7995,
  -43.8184,
  -43.8421,
  -43.8676,
  -43.8931,
  -43.9154,
  -43.9323,
  -43.9417,
  -43.9419,
  -43.9335,
  -43.9171,
  -43.8938,
  -43.8646,
  -43.831,
  -43.7951,
  -43.7556,
  -43.7117,
  -43.6633,
  -43.6094,
  -43.5471,
  -43.4737,
  -43.3902,
  -43.2971,
  -43.195,
  -43.0872,
  -42.9724,
  -42.8586,
  -42.7445,
  -42.6304,
  -42.5186,
  -42.4156,
  -42.3123,
  -42.2183,
  -42.1379,
  -42.0648,
  -41.9925,
  -41.9213,
  -41.8525,
  -41.7853,
  -41.7209,
  -41.6572,
  -41.6077,
  -41.5711,
  -41.5472,
  -41.54,
  -41.5538,
  -41.5876,
  -41.6416,
  -41.7135,
  -41.7991,
  -41.894,
  -41.9922,
  -42.0894,
  -42.1794,
  -42.2592,
  -42.3269,
  -42.3798,
  -42.4188,
  -42.4444,
  -42.4579,
  -42.4593,
  -42.4491,
  -42.4274,
  -42.3943,
  -42.3508,
  -42.299,
  -42.2411,
  -42.1801,
  -42.1205,
  -42.0634,
  -42.0116,
  -41.9659,
  -41.9272,
  -41.8957,
  -41.8702,
  -41.8508,
  -41.8369,
  -41.8287,
  -40.644,
  -40.6646,
  -40.6831,
  -40.701,
  -40.7192,
  -40.7389,
  -40.7604,
  -40.7837,
  -40.8094,
  -40.8375,
  -40.868,
  -40.9014,
  -40.9369,
  -40.9762,
  -41.0177,
  -41.0611,
  -41.1055,
  -41.1509,
  -41.1972,
  -41.2455,
  -41.2962,
  -41.3504,
  -41.4086,
  -41.4713,
  -41.5391,
  -41.6117,
  -41.689,
  -41.77,
  -41.8561,
  -41.9457,
  -42.0382,
  -42.1333,
  -42.2305,
  -42.329,
  -42.4281,
  -42.5271,
  -42.6253,
  -42.722,
  -42.8164,
  -42.9069,
  -42.9925,
  -43.0719,
  -43.1435,
  -43.2091,
  -43.2676,
  -43.3188,
  -43.3629,
  -43.3997,
  -43.4294,
  -43.4521,
  -43.4682,
  -43.4787,
  -43.4848,
  -43.4869,
  -43.4863,
  -43.4844,
  -43.4816,
  -43.4777,
  -43.471,
  -43.4621,
  -43.4485,
  -43.4299,
  -43.4068,
  -43.3806,
  -43.3522,
  -43.3218,
  -43.29,
  -43.2562,
  -43.2204,
  -43.1824,
  -43.1423,
  -43.1005,
  -43.0574,
  -43.0145,
  -42.9724,
  -42.9317,
  -42.8958,
  -42.8649,
  -42.8391,
  -42.818,
  -42.8011,
  -42.7884,
  -42.7786,
  -42.771,
  -42.7639,
  -42.7561,
  -42.7458,
  -42.7324,
  -42.716,
  -42.6978,
  -42.6785,
  -42.6594,
  -42.6406,
  -42.6205,
  -42.5996,
  -42.575,
  -42.5447,
  -42.5074,
  -42.4623,
  -42.4091,
  -42.3488,
  -42.2835,
  -42.2152,
  -42.1465,
  -42.0788,
  -42.0144,
  -41.9554,
  -41.9028,
  -41.8571,
  -41.8181,
  -41.7858,
  -41.7593,
  -41.7374,
  -41.7222,
  -41.7127,
  -41.7092,
  -41.7113,
  -41.7185,
  -41.7299,
  -41.7443,
  -41.7601,
  -41.7757,
  -41.7895,
  -41.8011,
  -41.8096,
  -41.8154,
  -41.8197,
  -41.8237,
  -41.8289,
  -41.8364,
  -41.847,
  -41.8604,
  -41.8747,
  -41.8899,
  -41.9024,
  -41.9101,
  -41.9107,
  -41.9033,
  -41.8879,
  -41.8652,
  -41.8368,
  -41.8047,
  -41.7707,
  -41.7365,
  -41.7026,
  -41.6695,
  -41.6368,
  -41.6041,
  -41.5699,
  -41.5338,
  -41.4951,
  -41.4535,
  -41.4094,
  -41.3637,
  -41.316,
  -41.2703,
  -41.2251,
  -41.1819,
  -41.1399,
  -41.1001,
  -41.0611,
  -41.0221,
  -40.9838,
  -40.9456,
  -40.9075,
  -40.8709,
  -40.8372,
  -40.8083,
  -40.7865,
  -40.7739,
  -40.7717,
  -40.7805,
  -40.7997,
  -40.8278,
  -40.8626,
  -40.9006,
  -40.9386,
  -40.9732,
  -41.0006,
  -41.0221,
  -41.0374,
  -41.0491,
  -41.0609,
  -41.0775,
  -41.1036,
  -41.1433,
  -41.1988,
  -41.2704,
  -41.3558,
  -41.4502,
  -41.5476,
  -41.6411,
  -41.725,
  -41.7953,
  -41.8515,
  -41.8958,
  -41.9358,
  -41.9793,
  -42.0356,
  -42.1128,
  -42.2146,
  -42.3397,
  -42.4829,
  -42.637,
  -42.7931,
  -42.9421,
  -43.0799,
  -43.2014,
  -43.3043,
  -43.388,
  -43.4549,
  -43.5063,
  -43.5456,
  -43.5756,
  -43.598,
  -43.6142,
  -43.6254,
  -43.6327,
  -43.6372,
  -43.6395,
  -43.6413,
  -43.6444,
  -43.6505,
  -43.661,
  -43.676,
  -43.6938,
  -43.7129,
  -43.7306,
  -43.7439,
  -43.7506,
  -43.7488,
  -43.7376,
  -43.7175,
  -43.6898,
  -43.6557,
  -43.6169,
  -43.5743,
  -43.5303,
  -43.4839,
  -43.4342,
  -43.3792,
  -43.3173,
  -43.2462,
  -43.1634,
  -43.0712,
  -42.9702,
  -42.8625,
  -42.7501,
  -42.6327,
  -42.5201,
  -42.4087,
  -42.2996,
  -42.1933,
  -42.0935,
  -41.9977,
  -41.9166,
  -41.8485,
  -41.7908,
  -41.7304,
  -41.6697,
  -41.6131,
  -41.5598,
  -41.5111,
  -41.4625,
  -41.4327,
  -41.4162,
  -41.4149,
  -41.4322,
  -41.4702,
  -41.5262,
  -41.6004,
  -41.6891,
  -41.7873,
  -41.8917,
  -41.9937,
  -42.091,
  -42.1792,
  -42.2544,
  -42.3155,
  -42.362,
  -42.3947,
  -42.4146,
  -42.4227,
  -42.4191,
  -42.404,
  -42.3767,
  -42.3371,
  -42.2855,
  -42.224,
  -42.1562,
  -42.0859,
  -42.0169,
  -41.9523,
  -41.8952,
  -41.8473,
  -41.8089,
  -41.7797,
  -41.7586,
  -41.744,
  -41.7351,
  -41.7311,
  -40.7144,
  -40.7362,
  -40.7554,
  -40.7735,
  -40.7916,
  -40.8109,
  -40.8324,
  -40.855,
  -40.8813,
  -40.91,
  -40.9415,
  -40.9764,
  -41.0147,
  -41.0564,
  -41.1004,
  -41.1464,
  -41.1939,
  -41.2423,
  -41.2917,
  -41.3432,
  -41.3974,
  -41.4549,
  -41.5154,
  -41.5809,
  -41.6506,
  -41.7246,
  -41.8025,
  -41.8837,
  -41.9678,
  -42.0543,
  -42.1431,
  -42.2338,
  -42.3262,
  -42.4193,
  -42.5125,
  -42.6051,
  -42.6961,
  -42.7842,
  -42.8704,
  -42.9528,
  -43.0305,
  -43.1026,
  -43.1686,
  -43.2284,
  -43.2817,
  -43.3287,
  -43.3696,
  -43.4043,
  -43.4329,
  -43.4555,
  -43.4724,
  -43.4841,
  -43.4916,
  -43.4947,
  -43.4961,
  -43.4962,
  -43.4958,
  -43.4942,
  -43.4909,
  -43.4845,
  -43.4734,
  -43.457,
  -43.4356,
  -43.4111,
  -43.3844,
  -43.3558,
  -43.3255,
  -43.2933,
  -43.2595,
  -43.2231,
  -43.1869,
  -43.1499,
  -43.1126,
  -43.0759,
  -43.04,
  -43.0061,
  -42.975,
  -42.9475,
  -42.924,
  -42.9042,
  -42.8881,
  -42.8754,
  -42.8654,
  -42.857,
  -42.85,
  -42.8428,
  -42.8344,
  -42.8228,
  -42.8098,
  -42.7947,
  -42.7783,
  -42.7613,
  -42.7442,
  -42.7261,
  -42.7064,
  -42.6832,
  -42.6547,
  -42.6201,
  -42.5784,
  -42.5293,
  -42.4739,
  -42.4134,
  -42.3496,
  -42.2848,
  -42.2205,
  -42.1585,
  -42.0996,
  -42.0474,
  -42.0016,
  -41.9625,
  -41.9303,
  -41.9048,
  -41.8853,
  -41.8714,
  -41.8636,
  -41.8619,
  -41.8662,
  -41.8754,
  -41.8893,
  -41.9064,
  -41.9253,
  -41.9437,
  -41.9606,
  -41.9744,
  -41.9847,
  -41.9908,
  -41.9955,
  -41.999,
  -42.0028,
  -42.0087,
  -42.0177,
  -42.0299,
  -42.0443,
  -42.0595,
  -42.0728,
  -42.082,
  -42.0846,
  -42.0795,
  -42.0666,
  -42.0466,
  -42.0212,
  -41.9927,
  -41.9626,
  -41.9325,
  -41.9029,
  -41.8744,
  -41.8463,
  -41.8166,
  -41.7861,
  -41.7525,
  -41.7155,
  -41.6746,
  -41.6303,
  -41.5837,
  -41.5353,
  -41.4877,
  -41.4399,
  -41.3938,
  -41.3494,
  -41.3058,
  -41.263,
  -41.2206,
  -41.1784,
  -41.1364,
  -41.095,
  -41.0555,
  -41.0191,
  -40.9875,
  -40.9632,
  -40.9477,
  -40.9407,
  -40.9445,
  -40.9574,
  -40.978,
  -41.0042,
  -41.033,
  -41.0617,
  -41.0868,
  -41.1063,
  -41.1195,
  -41.1271,
  -41.1317,
  -41.1362,
  -41.1457,
  -41.164,
  -41.1954,
  -41.2425,
  -41.306,
  -41.384,
  -41.4719,
  -41.5642,
  -41.6543,
  -41.7362,
  -41.8065,
  -41.864,
  -41.9112,
  -41.9531,
  -42.0001,
  -42.0587,
  -42.1375,
  -42.2379,
  -42.359,
  -42.4957,
  -42.6408,
  -42.7864,
  -42.9249,
  -43.0505,
  -43.1588,
  -43.2482,
  -43.3186,
  -43.3725,
  -43.4113,
  -43.4395,
  -43.4616,
  -43.4776,
  -43.4899,
  -43.4984,
  -43.505,
  -43.5093,
  -43.5122,
  -43.5147,
  -43.5179,
  -43.5234,
  -43.5316,
  -43.543,
  -43.5546,
  -43.5673,
  -43.5768,
  -43.5806,
  -43.5769,
  -43.5638,
  -43.5411,
  -43.5097,
  -43.4709,
  -43.4269,
  -43.3803,
  -43.3323,
  -43.2826,
  -43.2312,
  -43.1761,
  -43.1147,
  -43.0441,
  -42.9637,
  -42.8717,
  -42.7708,
  -42.663,
  -42.5496,
  -42.4307,
  -42.3043,
  -42.1984,
  -42.0867,
  -41.9774,
  -41.8747,
  -41.7934,
  -41.7223,
  -41.6565,
  -41.6052,
  -41.5531,
  -41.5018,
  -41.4527,
  -41.4097,
  -41.372,
  -41.3426,
  -41.3153,
  -41.3068,
  -41.312,
  -41.334,
  -41.3738,
  -41.4351,
  -41.5114,
  -41.6026,
  -41.7046,
  -41.8127,
  -41.9221,
  -42.0261,
  -42.1199,
  -42.2018,
  -42.2701,
  -42.3237,
  -42.3634,
  -42.3899,
  -42.4049,
  -42.4086,
  -42.4006,
  -42.3807,
  -42.3477,
  -42.3011,
  -42.241,
  -42.1696,
  -42.0906,
  -42.0087,
  -41.9287,
  -41.8551,
  -41.7913,
  -41.7391,
  -41.6989,
  -41.6698,
  -41.6499,
  -41.6375,
  -41.6313,
  -41.6298,
  -40.777,
  -40.8004,
  -40.8201,
  -40.8387,
  -40.857,
  -40.8765,
  -40.8979,
  -40.9225,
  -40.9491,
  -40.9782,
  -41.0107,
  -41.0466,
  -41.0863,
  -41.1295,
  -41.1754,
  -41.2236,
  -41.2724,
  -41.3232,
  -41.3756,
  -41.4299,
  -41.4868,
  -41.5471,
  -41.6109,
  -41.6787,
  -41.7503,
  -41.8255,
  -41.9036,
  -41.9844,
  -42.0672,
  -42.1514,
  -42.2374,
  -42.3245,
  -42.4117,
  -42.5001,
  -42.5881,
  -42.6747,
  -42.7592,
  -42.8412,
  -42.9199,
  -42.995,
  -43.0654,
  -43.1308,
  -43.1905,
  -43.2444,
  -43.2928,
  -43.3359,
  -43.3738,
  -43.4058,
  -43.4335,
  -43.4561,
  -43.4739,
  -43.4869,
  -43.4956,
  -43.5016,
  -43.5048,
  -43.5064,
  -43.5069,
  -43.5062,
  -43.5038,
  -43.4981,
  -43.488,
  -43.473,
  -43.4533,
  -43.43,
  -43.4036,
  -43.3763,
  -43.3473,
  -43.3166,
  -43.2849,
  -43.2522,
  -43.2194,
  -43.1871,
  -43.1553,
  -43.1244,
  -43.0945,
  -43.0663,
  -43.0401,
  -43.0164,
  -42.9955,
  -42.9777,
  -42.9629,
  -42.9502,
  -42.9402,
  -42.9323,
  -42.9255,
  -42.9191,
  -42.9123,
  -42.9043,
  -42.8944,
  -42.8829,
  -42.8694,
  -42.8548,
  -42.8391,
  -42.8222,
  -42.803,
  -42.7802,
  -42.7527,
  -42.7194,
  -42.6797,
  -42.6325,
  -42.5803,
  -42.5229,
  -42.4624,
  -42.4001,
  -42.3379,
  -42.2771,
  -42.2198,
  -42.1678,
  -42.1222,
  -42.0835,
  -42.0524,
  -42.0283,
  -42.0111,
  -42.0006,
  -41.9961,
  -41.9979,
  -42.0055,
  -42.0188,
  -42.0357,
  -42.057,
  -42.0798,
  -42.1024,
  -42.1233,
  -42.141,
  -42.1546,
  -42.164,
  -42.1701,
  -42.1743,
  -42.1785,
  -42.1838,
  -42.1919,
  -42.2031,
  -42.2167,
  -42.2316,
  -42.2451,
  -42.2547,
  -42.2583,
  -42.2543,
  -42.2432,
  -42.2242,
  -42.2015,
  -42.176,
  -42.1496,
  -42.1235,
  -42.0985,
  -42.0744,
  -42.0504,
  -42.0256,
  -41.9983,
  -41.9673,
  -41.932,
  -41.8916,
  -41.8468,
  -41.799,
  -41.7498,
  -41.6997,
  -41.6503,
  -41.6022,
  -41.5552,
  -41.5089,
  -41.4631,
  -41.4174,
  -41.3706,
  -41.3251,
  -41.2804,
  -41.2378,
  -41.1989,
  -41.1649,
  -41.1381,
  -41.1198,
  -41.1105,
  -41.1102,
  -41.1178,
  -41.1319,
  -41.1508,
  -41.172,
  -41.1932,
  -41.2112,
  -41.2245,
  -41.2324,
  -41.2354,
  -41.2358,
  -41.2362,
  -41.2409,
  -41.2537,
  -41.2785,
  -41.3184,
  -41.3731,
  -41.4429,
  -41.5228,
  -41.6076,
  -41.6913,
  -41.7685,
  -41.8355,
  -41.8916,
  -41.939,
  -41.9827,
  -42.0308,
  -42.0896,
  -42.1651,
  -42.2607,
  -42.3744,
  -42.5012,
  -42.6347,
  -42.7675,
  -42.8925,
  -43.0042,
  -43.0989,
  -43.1752,
  -43.2331,
  -43.2751,
  -43.3047,
  -43.3264,
  -43.3423,
  -43.3558,
  -43.3657,
  -43.3746,
  -43.3816,
  -43.3873,
  -43.3916,
  -43.3949,
  -43.3994,
  -43.4046,
  -43.4112,
  -43.4204,
  -43.4289,
  -43.435,
  -43.4361,
  -43.4314,
  -43.4178,
  -43.3942,
  -43.361,
  -43.3194,
  -43.2718,
  -43.221,
  -43.1691,
  -43.1165,
  -43.0637,
  -43.0087,
  -42.9487,
  -42.8805,
  -42.8021,
  -42.7124,
  -42.6106,
  -42.501,
  -42.387,
  -42.2677,
  -42.134,
  -41.9962,
  -41.884,
  -41.7855,
  -41.7047,
  -41.6259,
  -41.5801,
  -41.5269,
  -41.4676,
  -41.4167,
  -41.3728,
  -41.3309,
  -41.2929,
  -41.2632,
  -41.2402,
  -41.227,
  -41.2214,
  -41.2358,
  -41.2605,
  -41.3075,
  -41.3684,
  -41.4482,
  -41.5397,
  -41.6426,
  -41.754,
  -41.8668,
  -41.9764,
  -42.0771,
  -42.1655,
  -42.2402,
  -42.3004,
  -42.3467,
  -42.3801,
  -42.4019,
  -42.4128,
  -42.4124,
  -42.4001,
  -42.375,
  -42.3356,
  -42.2809,
  -42.2114,
  -42.1291,
  -42.0375,
  -41.9438,
  -41.8526,
  -41.7694,
  -41.6978,
  -41.6399,
  -41.5959,
  -41.5644,
  -41.5437,
  -41.5315,
  -41.526,
  -41.5255,
  -40.8325,
  -40.858,
  -40.8802,
  -40.9001,
  -40.9192,
  -40.9391,
  -40.9611,
  -40.9857,
  -41.0129,
  -41.0431,
  -41.0762,
  -41.1119,
  -41.1526,
  -41.1969,
  -41.2439,
  -41.2935,
  -41.3451,
  -41.398,
  -41.4528,
  -41.5092,
  -41.5682,
  -41.6302,
  -41.6958,
  -41.7649,
  -41.8374,
  -41.9132,
  -41.9905,
  -42.0709,
  -42.1527,
  -42.2352,
  -42.3192,
  -42.4035,
  -42.488,
  -42.5726,
  -42.6556,
  -42.7373,
  -42.8162,
  -42.8918,
  -42.9639,
  -43.032,
  -43.0959,
  -43.1548,
  -43.2075,
  -43.256,
  -43.2998,
  -43.3393,
  -43.3744,
  -43.4057,
  -43.4327,
  -43.4556,
  -43.4741,
  -43.4881,
  -43.4987,
  -43.5061,
  -43.5102,
  -43.5122,
  -43.513,
  -43.5123,
  -43.5083,
  -43.5025,
  -43.4926,
  -43.478,
  -43.4592,
  -43.4371,
  -43.4126,
  -43.3863,
  -43.3588,
  -43.3295,
  -43.2997,
  -43.2697,
  -43.24,
  -43.2114,
  -43.1842,
  -43.1584,
  -43.1338,
  -43.1095,
  -43.0878,
  -43.0678,
  -43.05,
  -43.0346,
  -43.0216,
  -43.0111,
  -43.0023,
  -42.9951,
  -42.9892,
  -42.9842,
  -42.9792,
  -42.9736,
  -42.9666,
  -42.9584,
  -42.9482,
  -42.9361,
  -42.9224,
  -42.9054,
  -42.8865,
  -42.8639,
  -42.8364,
  -42.8036,
  -42.765,
  -42.7206,
  -42.6702,
  -42.6148,
  -42.5556,
  -42.495,
  -42.4333,
  -42.3732,
  -42.3159,
  -42.264,
  -42.2189,
  -42.1816,
  -42.1525,
  -42.1315,
  -42.1172,
  -42.1112,
  -42.1118,
  -42.1187,
  -42.1314,
  -42.1498,
  -42.1728,
  -42.1992,
  -42.227,
  -42.2546,
  -42.2803,
  -42.3027,
  -42.3203,
  -42.333,
  -42.3417,
  -42.3478,
  -42.3529,
  -42.3589,
  -42.3667,
  -42.3771,
  -42.389,
  -42.4032,
  -42.4163,
  -42.4255,
  -42.4289,
  -42.4253,
  -42.4149,
  -42.3983,
  -42.3774,
  -42.3545,
  -42.3312,
  -42.3088,
  -42.2877,
  -42.2676,
  -42.2474,
  -42.2261,
  -42.2017,
  -42.1726,
  -42.1388,
  -42.099,
  -42.0542,
  -42.0061,
  -41.9555,
  -41.905,
  -41.8545,
  -41.8051,
  -41.7568,
  -41.7092,
  -41.6611,
  -41.6128,
  -41.5641,
  -41.5156,
  -41.4681,
  -41.423,
  -41.3814,
  -41.3456,
  -41.3167,
  -41.296,
  -41.2837,
  -41.2795,
  -41.2823,
  -41.2914,
  -41.3043,
  -41.3201,
  -41.3357,
  -41.3491,
  -41.3577,
  -41.363,
  -41.3643,
  -41.3632,
  -41.3621,
  -41.3641,
  -41.3731,
  -41.3924,
  -41.4256,
  -41.4733,
  -41.534,
  -41.6041,
  -41.6787,
  -41.7528,
  -41.8216,
  -41.882,
  -41.9338,
  -41.9784,
  -42.0204,
  -42.0664,
  -42.122,
  -42.193,
  -42.281,
  -42.3846,
  -42.4996,
  -42.6193,
  -42.7379,
  -42.8476,
  -42.9456,
  -43.0272,
  -43.0915,
  -43.1388,
  -43.1722,
  -43.1951,
  -43.2122,
  -43.2263,
  -43.239,
  -43.2505,
  -43.2608,
  -43.2689,
  -43.2759,
  -43.2821,
  -43.2866,
  -43.2913,
  -43.2961,
  -43.3022,
  -43.3088,
  -43.3135,
  -43.314,
  -43.3091,
  -43.2957,
  -43.2734,
  -43.241,
  -43.1993,
  -43.1505,
  -43.0969,
  -43.0416,
  -42.9855,
  -42.9315,
  -42.8767,
  -42.8191,
  -42.7546,
  -42.6804,
  -42.5943,
  -42.4957,
  -42.3858,
  -42.2693,
  -42.1492,
  -42.0216,
  -41.8862,
  -41.7471,
  -41.6445,
  -41.5706,
  -41.519,
  -41.4738,
  -41.4408,
  -41.3966,
  -41.3506,
  -41.2979,
  -41.253,
  -41.2139,
  -41.1901,
  -41.1871,
  -41.1835,
  -41.1897,
  -41.2002,
  -41.23,
  -41.2751,
  -41.3333,
  -41.4088,
  -41.4978,
  -41.5991,
  -41.7102,
  -41.8249,
  -41.9378,
  -42.0438,
  -42.1388,
  -42.2201,
  -42.2874,
  -42.3407,
  -42.3804,
  -42.4086,
  -42.4265,
  -42.434,
  -42.4298,
  -42.4132,
  -42.3825,
  -42.3359,
  -42.2725,
  -42.1928,
  -42.0995,
  -41.9969,
  -41.8913,
  -41.7893,
  -41.696,
  -41.616,
  -41.5512,
  -41.5018,
  -41.4663,
  -41.443,
  -41.4287,
  -41.4223,
  -41.4213,
  -40.8845,
  -40.9125,
  -40.9367,
  -40.958,
  -40.9783,
  -40.9989,
  -41.0215,
  -41.0457,
  -41.0735,
  -41.1044,
  -41.1385,
  -41.1761,
  -41.2172,
  -41.2619,
  -41.3098,
  -41.3603,
  -41.4131,
  -41.4676,
  -41.5239,
  -41.5817,
  -41.6417,
  -41.7036,
  -41.7696,
  -41.839,
  -41.9119,
  -41.9875,
  -42.0654,
  -42.1454,
  -42.2267,
  -42.3082,
  -42.3903,
  -42.4725,
  -42.5543,
  -42.6351,
  -42.7147,
  -42.7915,
  -42.8654,
  -42.9344,
  -43.0005,
  -43.0625,
  -43.1202,
  -43.1733,
  -43.2216,
  -43.2651,
  -43.3048,
  -43.3408,
  -43.3735,
  -43.4031,
  -43.4294,
  -43.4522,
  -43.4714,
  -43.4866,
  -43.4971,
  -43.5055,
  -43.5107,
  -43.513,
  -43.5136,
  -43.5116,
  -43.5073,
  -43.5003,
  -43.4897,
  -43.4753,
  -43.4572,
  -43.4355,
  -43.4118,
  -43.3866,
  -43.3604,
  -43.333,
  -43.3049,
  -43.276,
  -43.2492,
  -43.2233,
  -43.1997,
  -43.1776,
  -43.1571,
  -43.1379,
  -43.1201,
  -43.1035,
  -43.0887,
  -43.0755,
  -43.0645,
  -43.0557,
  -43.0484,
  -43.0428,
  -43.0385,
  -43.035,
  -43.032,
  -43.0278,
  -43.0238,
  -43.0186,
  -43.0117,
  -43.0023,
  -42.9906,
  -42.976,
  -42.9577,
  -42.9352,
  -42.9077,
  -42.8751,
  -42.8369,
  -42.7931,
  -42.7437,
  -42.6895,
  -42.6309,
  -42.57,
  -42.5084,
  -42.4471,
  -42.3901,
  -42.3386,
  -42.2946,
  -42.2594,
  -42.2336,
  -42.2169,
  -42.2092,
  -42.2091,
  -42.2165,
  -42.2299,
  -42.2491,
  -42.2737,
  -42.3026,
  -42.3344,
  -42.3677,
  -42.4006,
  -42.4315,
  -42.4587,
  -42.4807,
  -42.4963,
  -42.5082,
  -42.5165,
  -42.5235,
  -42.5311,
  -42.5392,
  -42.5493,
  -42.5616,
  -42.5748,
  -42.5865,
  -42.5947,
  -42.5973,
  -42.5932,
  -42.5826,
  -42.5666,
  -42.5472,
  -42.5261,
  -42.5054,
  -42.486,
  -42.4682,
  -42.4515,
  -42.4335,
  -42.4149,
  -42.3929,
  -42.3658,
  -42.3331,
  -42.2942,
  -42.2506,
  -42.2034,
  -42.1542,
  -42.1043,
  -42.0542,
  -42.0051,
  -41.957,
  -41.9093,
  -41.8606,
  -41.8109,
  -41.7603,
  -41.7098,
  -41.6602,
  -41.6128,
  -41.5694,
  -41.5314,
  -41.5004,
  -41.4764,
  -41.4619,
  -41.4545,
  -41.4534,
  -41.4578,
  -41.4664,
  -41.4778,
  -41.4901,
  -41.501,
  -41.5091,
  -41.514,
  -41.5156,
  -41.5149,
  -41.5132,
  -41.5141,
  -41.52,
  -41.5348,
  -41.5612,
  -41.6,
  -41.6503,
  -41.7085,
  -41.7705,
  -41.8321,
  -41.8893,
  -41.9404,
  -41.9845,
  -42.0222,
  -42.0604,
  -42.1023,
  -42.1532,
  -42.2177,
  -42.2966,
  -42.3887,
  -42.4909,
  -42.5969,
  -42.7008,
  -42.797,
  -42.8816,
  -42.9513,
  -43.0051,
  -43.0441,
  -43.0712,
  -43.0904,
  -43.1056,
  -43.1195,
  -43.1339,
  -43.1463,
  -43.1577,
  -43.1675,
  -43.1755,
  -43.1819,
  -43.1871,
  -43.1917,
  -43.1964,
  -43.2014,
  -43.2049,
  -43.2063,
  -43.2027,
  -43.1922,
  -43.1726,
  -43.1432,
  -43.1039,
  -43.0563,
  -43.0029,
  -42.9463,
  -42.8894,
  -42.834,
  -42.7806,
  -42.7256,
  -42.6662,
  -42.5968,
  -42.517,
  -42.4235,
  -42.3171,
  -42.2005,
  -42.0793,
  -41.9558,
  -41.827,
  -41.6989,
  -41.5762,
  -41.4913,
  -41.4378,
  -41.3975,
  -41.3655,
  -41.3393,
  -41.3079,
  -41.2733,
  -41.2328,
  -41.1956,
  -41.1743,
  -41.1648,
  -41.1737,
  -41.1879,
  -41.2077,
  -41.2299,
  -41.2733,
  -41.3281,
  -41.3956,
  -41.4769,
  -41.5739,
  -41.6802,
  -41.7932,
  -41.9073,
  -42.017,
  -42.1185,
  -42.2067,
  -42.2809,
  -42.3414,
  -42.3886,
  -42.4238,
  -42.4482,
  -42.4627,
  -42.4671,
  -42.4597,
  -42.4386,
  -42.4017,
  -42.3472,
  -42.2748,
  -42.185,
  -42.0805,
  -41.9669,
  -41.85,
  -41.7371,
  -41.6341,
  -41.5453,
  -41.4731,
  -41.4171,
  -41.3763,
  -41.3483,
  -41.3307,
  -41.3215,
  -41.3189,
  -40.9339,
  -40.9643,
  -40.9896,
  -41.0127,
  -41.034,
  -41.0559,
  -41.0794,
  -41.1052,
  -41.1339,
  -41.1656,
  -41.2004,
  -41.2386,
  -41.2803,
  -41.3251,
  -41.3734,
  -41.4244,
  -41.477,
  -41.5325,
  -41.5894,
  -41.6479,
  -41.7081,
  -41.7705,
  -41.836,
  -41.9049,
  -41.9768,
  -42.0517,
  -42.1287,
  -42.2081,
  -42.2883,
  -42.3696,
  -42.4504,
  -42.5298,
  -42.6095,
  -42.6876,
  -42.7635,
  -42.8363,
  -42.9056,
  -42.9705,
  -43.0311,
  -43.0876,
  -43.1398,
  -43.1878,
  -43.2313,
  -43.2706,
  -43.3066,
  -43.3394,
  -43.3697,
  -43.3965,
  -43.4219,
  -43.4446,
  -43.464,
  -43.4799,
  -43.492,
  -43.501,
  -43.5068,
  -43.5091,
  -43.5087,
  -43.5056,
  -43.4998,
  -43.4912,
  -43.4798,
  -43.4649,
  -43.4467,
  -43.4248,
  -43.4018,
  -43.3777,
  -43.3528,
  -43.3273,
  -43.3014,
  -43.2758,
  -43.2503,
  -43.2266,
  -43.2052,
  -43.1854,
  -43.1678,
  -43.1516,
  -43.1367,
  -43.1232,
  -43.1107,
  -43.0996,
  -43.0905,
  -43.0825,
  -43.0772,
  -43.0735,
  -43.0711,
  -43.0697,
  -43.0689,
  -43.0679,
  -43.0667,
  -43.0646,
  -43.0609,
  -43.0546,
  -43.0452,
  -43.0321,
  -43.0148,
  -42.9927,
  -42.9653,
  -42.9331,
  -42.8952,
  -42.8508,
  -42.8018,
  -42.7475,
  -42.6891,
  -42.6279,
  -42.566,
  -42.5056,
  -42.4488,
  -42.3981,
  -42.3562,
  -42.324,
  -42.3024,
  -42.2914,
  -42.2905,
  -42.298,
  -42.313,
  -42.3342,
  -42.3613,
  -42.3928,
  -42.4268,
  -42.4644,
  -42.5028,
  -42.5406,
  -42.5761,
  -42.6076,
  -42.6339,
  -42.6541,
  -42.6691,
  -42.6803,
  -42.6894,
  -42.6983,
  -42.7074,
  -42.7177,
  -42.7295,
  -42.7414,
  -42.7519,
  -42.7584,
  -42.7596,
  -42.7547,
  -42.7436,
  -42.7268,
  -42.7083,
  -42.6889,
  -42.6702,
  -42.6533,
  -42.6383,
  -42.6244,
  -42.6101,
  -42.5939,
  -42.5738,
  -42.5485,
  -42.5173,
  -42.48,
  -42.4381,
  -42.3922,
  -42.3449,
  -42.2976,
  -42.2498,
  -42.202,
  -42.1558,
  -42.1085,
  -42.0603,
  -42.0098,
  -41.9596,
  -41.9078,
  -41.8568,
  -41.8082,
  -41.7635,
  -41.7239,
  -41.6915,
  -41.6665,
  -41.6491,
  -41.6387,
  -41.6342,
  -41.6348,
  -41.6397,
  -41.6478,
  -41.6576,
  -41.6672,
  -41.6751,
  -41.6807,
  -41.6832,
  -41.6837,
  -41.6827,
  -41.6827,
  -41.6859,
  -41.6964,
  -41.7145,
  -41.7438,
  -41.7821,
  -41.8269,
  -41.8744,
  -41.9213,
  -41.9646,
  -42.0034,
  -42.0381,
  -42.0697,
  -42.1016,
  -42.1382,
  -42.1827,
  -42.2401,
  -42.3099,
  -42.3909,
  -42.4805,
  -42.5728,
  -42.6628,
  -42.746,
  -42.8182,
  -42.8771,
  -42.9222,
  -42.9549,
  -42.9779,
  -42.9953,
  -43.0104,
  -43.0248,
  -43.0392,
  -43.0538,
  -43.0656,
  -43.0759,
  -43.0835,
  -43.0892,
  -43.0936,
  -43.0979,
  -43.102,
  -43.1059,
  -43.1085,
  -43.1073,
  -43.1006,
  -43.0859,
  -43.062,
  -43.0276,
  -42.9841,
  -42.9331,
  -42.878,
  -42.8215,
  -42.7659,
  -42.712,
  -42.6595,
  -42.6047,
  -42.544,
  -42.4716,
  -42.3862,
  -42.2866,
  -42.1736,
  -42.0524,
  -41.9279,
  -41.8041,
  -41.6791,
  -41.5604,
  -41.4637,
  -41.3976,
  -41.3494,
  -41.3132,
  -41.2847,
  -41.265,
  -41.2435,
  -41.2228,
  -41.2016,
  -41.1835,
  -41.179,
  -41.1861,
  -41.2027,
  -41.2274,
  -41.2578,
  -41.292,
  -41.3433,
  -41.4064,
  -41.4795,
  -41.5663,
  -41.6655,
  -41.7726,
  -41.8835,
  -41.9942,
  -42.0984,
  -42.1932,
  -42.2746,
  -42.3428,
  -42.398,
  -42.441,
  -42.4729,
  -42.4948,
  -42.5067,
  -42.5081,
  -42.4972,
  -42.4715,
  -42.4285,
  -42.3665,
  -42.285,
  -42.1857,
  -42.0701,
  -41.9457,
  -41.8186,
  -41.6958,
  -41.5836,
  -41.4865,
  -41.4061,
  -41.3428,
  -41.296,
  -41.2621,
  -41.2393,
  -41.2259,
  -41.2198,
  -40.9803,
  -41.0134,
  -41.0413,
  -41.0662,
  -41.0892,
  -41.1128,
  -41.1371,
  -41.164,
  -41.1936,
  -41.226,
  -41.2615,
  -41.2991,
  -41.341,
  -41.3864,
  -41.435,
  -41.4863,
  -41.5401,
  -41.5956,
  -41.6526,
  -41.7109,
  -41.7703,
  -41.8316,
  -41.8955,
  -41.9627,
  -42.0331,
  -42.1064,
  -42.1814,
  -42.2593,
  -42.339,
  -42.4193,
  -42.4992,
  -42.5781,
  -42.6558,
  -42.7314,
  -42.8041,
  -42.8731,
  -42.9382,
  -42.9986,
  -43.0541,
  -43.1057,
  -43.153,
  -43.1963,
  -43.235,
  -43.2706,
  -43.3033,
  -43.3334,
  -43.3612,
  -43.3873,
  -43.4116,
  -43.4337,
  -43.4531,
  -43.4691,
  -43.4817,
  -43.4908,
  -43.4965,
  -43.4989,
  -43.4977,
  -43.4932,
  -43.4853,
  -43.4756,
  -43.4626,
  -43.4469,
  -43.4287,
  -43.4083,
  -43.386,
  -43.3632,
  -43.34,
  -43.3165,
  -43.2928,
  -43.2689,
  -43.2445,
  -43.2218,
  -43.2013,
  -43.1828,
  -43.1668,
  -43.1516,
  -43.1386,
  -43.1271,
  -43.1165,
  -43.1072,
  -43.0998,
  -43.0947,
  -43.0914,
  -43.0898,
  -43.0897,
  -43.0906,
  -43.0919,
  -43.0935,
  -43.095,
  -43.0956,
  -43.0947,
  -43.0914,
  -43.0834,
  -43.072,
  -43.0564,
  -43.0352,
  -43.0089,
  -42.9773,
  -42.9401,
  -42.8972,
  -42.8485,
  -42.7946,
  -42.7361,
  -42.6747,
  -42.6126,
  -42.5523,
  -42.4963,
  -42.4474,
  -42.4077,
  -42.3795,
  -42.3632,
  -42.3577,
  -42.3643,
  -42.3805,
  -42.4044,
  -42.4344,
  -42.4691,
  -42.5078,
  -42.5492,
  -42.5919,
  -42.6347,
  -42.6766,
  -42.7157,
  -42.7505,
  -42.7799,
  -42.8032,
  -42.821,
  -42.8345,
  -42.8456,
  -42.8558,
  -42.866,
  -42.8765,
  -42.8866,
  -42.8974,
  -42.9061,
  -42.9112,
  -42.9112,
  -42.9052,
  -42.8938,
  -42.8783,
  -42.8605,
  -42.8425,
  -42.8256,
  -42.811,
  -42.7985,
  -42.787,
  -42.7751,
  -42.761,
  -42.7428,
  -42.7194,
  -42.6901,
  -42.6549,
  -42.6153,
  -42.5713,
  -42.5271,
  -42.4824,
  -42.4378,
  -42.3937,
  -42.3497,
  -42.3053,
  -42.2592,
  -42.2113,
  -42.1611,
  -42.1102,
  -42.0597,
  -42.0113,
  -41.9656,
  -41.9253,
  -41.8912,
  -41.8644,
  -41.8447,
  -41.8313,
  -41.8231,
  -41.8201,
  -41.8218,
  -41.8269,
  -41.8346,
  -41.8419,
  -41.8498,
  -41.8562,
  -41.8601,
  -41.8615,
  -41.8608,
  -41.86,
  -41.8612,
  -41.8661,
  -41.8781,
  -41.8966,
  -41.9227,
  -41.9528,
  -41.9848,
  -42.0161,
  -42.0449,
  -42.0706,
  -42.0942,
  -42.1175,
  -42.1423,
  -42.1724,
  -42.211,
  -42.2605,
  -42.3218,
  -42.3932,
  -42.471,
  -42.5513,
  -42.6278,
  -42.6987,
  -42.7597,
  -42.8092,
  -42.8471,
  -42.8751,
  -42.8954,
  -42.9119,
  -42.9272,
  -42.9422,
  -42.9572,
  -42.9715,
  -42.9837,
  -42.9931,
  -42.9996,
  -43.004,
  -43.0074,
  -43.0102,
  -43.0131,
  -43.0158,
  -43.0173,
  -43.014,
  -43.005,
  -42.988,
  -42.9612,
  -42.9241,
  -42.8788,
  -42.8274,
  -42.773,
  -42.7192,
  -42.667,
  -42.6156,
  -42.5653,
  -42.5108,
  -42.4488,
  -42.3735,
  -42.2836,
  -42.179,
  -42.0617,
  -41.9374,
  -41.8117,
  -41.6898,
  -41.574,
  -41.4709,
  -41.3892,
  -41.3329,
  -41.2927,
  -41.2672,
  -41.2474,
  -41.2418,
  -41.2356,
  -41.2297,
  -41.2234,
  -41.2251,
  -41.2329,
  -41.2481,
  -41.2704,
  -41.3003,
  -41.3378,
  -41.3796,
  -41.4348,
  -41.5007,
  -41.5773,
  -41.6645,
  -41.7619,
  -41.8661,
  -41.9733,
  -42.0783,
  -42.1759,
  -42.2638,
  -42.34,
  -42.4033,
  -42.4546,
  -42.4946,
  -42.5245,
  -42.5449,
  -42.5548,
  -42.5537,
  -42.5392,
  -42.5086,
  -42.4599,
  -42.3911,
  -42.302,
  -42.194,
  -42.0704,
  -41.937,
  -41.8007,
  -41.669,
  -41.548,
  -41.4422,
  -41.3535,
  -41.2823,
  -41.2275,
  -41.1869,
  -41.1588,
  -41.14,
  -41.1281,
  -41.0263,
  -41.0603,
  -41.0905,
  -41.1173,
  -41.1425,
  -41.1675,
  -41.1925,
  -41.2204,
  -41.251,
  -41.2841,
  -41.3201,
  -41.3593,
  -41.4019,
  -41.4477,
  -41.4966,
  -41.5479,
  -41.6015,
  -41.6568,
  -41.7133,
  -41.7705,
  -41.8287,
  -41.8873,
  -41.9492,
  -42.014,
  -42.0821,
  -42.1531,
  -42.2272,
  -42.3037,
  -42.3819,
  -42.461,
  -42.5397,
  -42.617,
  -42.6925,
  -42.7658,
  -42.8351,
  -42.9006,
  -42.9605,
  -43.0167,
  -43.068,
  -43.1152,
  -43.1583,
  -43.1979,
  -43.234,
  -43.2666,
  -43.2962,
  -43.3238,
  -43.3496,
  -43.3738,
  -43.3965,
  -43.4178,
  -43.4365,
  -43.4527,
  -43.464,
  -43.4733,
  -43.4791,
  -43.4812,
  -43.4794,
  -43.4739,
  -43.4656,
  -43.4545,
  -43.4409,
  -43.4247,
  -43.4062,
  -43.3863,
  -43.365,
  -43.3436,
  -43.3221,
  -43.3006,
  -43.2787,
  -43.2551,
  -43.2321,
  -43.2099,
  -43.1891,
  -43.171,
  -43.1552,
  -43.1416,
  -43.1298,
  -43.1193,
  -43.1101,
  -43.1025,
  -43.0967,
  -43.0932,
  -43.092,
  -43.0925,
  -43.0945,
  -43.0975,
  -43.1,
  -43.1043,
  -43.1083,
  -43.1117,
  -43.1135,
  -43.1125,
  -43.1077,
  -43.0988,
  -43.0849,
  -43.0655,
  -43.041,
  -43.0111,
  -42.9752,
  -42.9334,
  -42.8856,
  -42.8324,
  -42.7743,
  -42.7135,
  -42.6522,
  -42.5918,
  -42.5373,
  -42.4907,
  -42.4541,
  -42.4303,
  -42.4197,
  -42.4223,
  -42.4372,
  -42.4625,
  -42.4957,
  -42.5345,
  -42.5772,
  -42.6226,
  -42.6696,
  -42.7168,
  -42.7631,
  -42.8073,
  -42.8484,
  -42.8852,
  -42.9167,
  -42.9409,
  -42.9606,
  -42.976,
  -42.9887,
  -43.0001,
  -43.011,
  -43.0217,
  -43.0322,
  -43.0416,
  -43.0491,
  -43.0531,
  -43.0522,
  -43.0456,
  -43.0342,
  -43.0192,
  -43.0026,
  -42.9861,
  -42.9712,
  -42.9587,
  -42.9483,
  -42.939,
  -42.9281,
  -42.916,
  -42.9001,
  -42.8785,
  -42.851,
  -42.8182,
  -42.781,
  -42.7415,
  -42.7009,
  -42.6603,
  -42.6193,
  -42.5797,
  -42.5398,
  -42.4982,
  -42.4551,
  -42.4095,
  -42.3618,
  -42.3129,
  -42.2639,
  -42.2165,
  -42.1715,
  -42.1309,
  -42.0963,
  -42.0673,
  -42.0452,
  -42.0285,
  -42.0172,
  -42.0102,
  -42.0082,
  -42.0106,
  -42.0156,
  -42.0227,
  -42.0301,
  -42.0367,
  -42.0412,
  -42.0433,
  -42.043,
  -42.0408,
  -42.0387,
  -42.0388,
  -42.0428,
  -42.0513,
  -42.0638,
  -42.0797,
  -42.096,
  -42.1115,
  -42.1258,
  -42.1389,
  -42.1516,
  -42.1648,
  -42.1823,
  -42.2059,
  -42.2386,
  -42.2817,
  -42.3351,
  -42.3977,
  -42.4658,
  -42.5353,
  -42.602,
  -42.662,
  -42.7132,
  -42.7544,
  -42.7861,
  -42.8098,
  -42.8283,
  -42.8437,
  -42.8582,
  -42.8728,
  -42.8867,
  -42.8992,
  -42.9098,
  -42.9173,
  -42.922,
  -42.9246,
  -42.9263,
  -42.9275,
  -42.9304,
  -42.9321,
  -42.93,
  -42.9253,
  -42.9152,
  -42.8968,
  -42.8686,
  -42.8312,
  -42.7863,
  -42.7368,
  -42.6858,
  -42.6364,
  -42.5885,
  -42.5421,
  -42.4942,
  -42.4406,
  -42.3772,
  -42.2994,
  -42.2066,
  -42.0989,
  -41.9795,
  -41.8544,
  -41.7297,
  -41.611,
  -41.5038,
  -41.4134,
  -41.3403,
  -41.2934,
  -41.2627,
  -41.247,
  -41.2423,
  -41.2472,
  -41.2526,
  -41.2592,
  -41.268,
  -41.2804,
  -41.3012,
  -41.3233,
  -41.353,
  -41.389,
  -41.4314,
  -41.4775,
  -41.5349,
  -41.6005,
  -41.6761,
  -41.7605,
  -41.8536,
  -41.9533,
  -42.056,
  -42.1555,
  -42.2479,
  -42.3312,
  -42.403,
  -42.4632,
  -42.5121,
  -42.5504,
  -42.579,
  -42.598,
  -42.6065,
  -42.603,
  -42.585,
  -42.5504,
  -42.4966,
  -42.4221,
  -42.3269,
  -42.2121,
  -42.0815,
  -41.9408,
  -41.797,
  -41.6573,
  -41.5279,
  -41.4136,
  -41.3162,
  -41.2362,
  -41.1727,
  -41.1242,
  -41.0888,
  -41.0637,
  -41.0463,
  -41.07,
  -41.1049,
  -41.1349,
  -41.1639,
  -41.1914,
  -41.2184,
  -41.2461,
  -41.2756,
  -41.3073,
  -41.3413,
  -41.378,
  -41.418,
  -41.4612,
  -41.5075,
  -41.5568,
  -41.6081,
  -41.6602,
  -41.7149,
  -41.7703,
  -41.8262,
  -41.8829,
  -41.9405,
  -41.9998,
  -42.0622,
  -42.1275,
  -42.1958,
  -42.267,
  -42.3413,
  -42.4176,
  -42.4949,
  -42.572,
  -42.6465,
  -42.7195,
  -42.7899,
  -42.8557,
  -42.9173,
  -42.9744,
  -43.0269,
  -43.0747,
  -43.1186,
  -43.1587,
  -43.1951,
  -43.2282,
  -43.2581,
  -43.2854,
  -43.3104,
  -43.3338,
  -43.3549,
  -43.3759,
  -43.3956,
  -43.4136,
  -43.4289,
  -43.4416,
  -43.4506,
  -43.4563,
  -43.4581,
  -43.4562,
  -43.4501,
  -43.4407,
  -43.4286,
  -43.4141,
  -43.3976,
  -43.3795,
  -43.3591,
  -43.3392,
  -43.319,
  -43.2995,
  -43.2797,
  -43.2595,
  -43.2382,
  -43.2158,
  -43.1936,
  -43.1724,
  -43.1535,
  -43.1374,
  -43.1235,
  -43.1116,
  -43.1015,
  -43.0933,
  -43.087,
  -43.0818,
  -43.0799,
  -43.0805,
  -43.083,
  -43.0867,
  -43.0917,
  -43.0973,
  -43.1038,
  -43.1103,
  -43.1163,
  -43.1206,
  -43.1218,
  -43.1195,
  -43.1127,
  -43.1013,
  -43.0847,
  -43.0627,
  -43.0351,
  -43.0003,
  -42.9605,
  -42.9143,
  -42.8626,
  -42.8062,
  -42.7469,
  -42.6873,
  -42.6296,
  -42.5776,
  -42.534,
  -42.5018,
  -42.4827,
  -42.4782,
  -42.4881,
  -42.5114,
  -42.5455,
  -42.5874,
  -42.6345,
  -42.6844,
  -42.7357,
  -42.7861,
  -42.8365,
  -42.8846,
  -42.9299,
  -42.9715,
  -43.0086,
  -43.0406,
  -43.0668,
  -43.0875,
  -43.104,
  -43.1179,
  -43.1303,
  -43.1416,
  -43.1523,
  -43.162,
  -43.1704,
  -43.1768,
  -43.1801,
  -43.179,
  -43.1727,
  -43.1613,
  -43.1477,
  -43.1325,
  -43.1178,
  -43.105,
  -43.0945,
  -43.086,
  -43.0786,
  -43.0705,
  -43.0602,
  -43.046,
  -43.0266,
  -43.0009,
  -42.9702,
  -42.9362,
  -42.9005,
  -42.8637,
  -42.8269,
  -42.7905,
  -42.7546,
  -42.7183,
  -42.681,
  -42.6413,
  -42.5982,
  -42.554,
  -42.5083,
  -42.4622,
  -42.417,
  -42.3739,
  -42.3348,
  -42.3003,
  -42.2715,
  -42.2478,
  -42.2283,
  -42.213,
  -42.2027,
  -42.1969,
  -42.1956,
  -42.198,
  -42.2031,
  -42.2092,
  -42.2151,
  -42.2195,
  -42.2212,
  -42.2199,
  -42.2167,
  -42.2112,
  -42.2062,
  -42.2019,
  -42.2006,
  -42.2009,
  -42.203,
  -42.2048,
  -42.2063,
  -42.2073,
  -42.2084,
  -42.211,
  -42.2167,
  -42.2272,
  -42.2448,
  -42.2717,
  -42.3088,
  -42.3557,
  -42.4106,
  -42.4702,
  -42.5303,
  -42.5872,
  -42.6376,
  -42.6802,
  -42.7142,
  -42.7403,
  -42.7604,
  -42.7763,
  -42.7898,
  -42.8024,
  -42.8134,
  -42.8249,
  -42.835,
  -42.8431,
  -42.8481,
  -42.8506,
  -42.8515,
  -42.852,
  -42.8526,
  -42.8542,
  -42.8544,
  -42.8526,
  -42.8464,
  -42.8347,
  -42.8158,
  -42.7877,
  -42.7514,
  -42.7088,
  -42.6632,
  -42.6174,
  -42.5729,
  -42.5297,
  -42.4871,
  -42.4416,
  -42.3885,
  -42.3243,
  -42.245,
  -42.1509,
  -42.0423,
  -41.9234,
  -41.7997,
  -41.6776,
  -41.5633,
  -41.4615,
  -41.3789,
  -41.3137,
  -41.2729,
  -41.2514,
  -41.2456,
  -41.2513,
  -41.2663,
  -41.2833,
  -41.3024,
  -41.3239,
  -41.348,
  -41.3789,
  -41.4101,
  -41.446,
  -41.4859,
  -41.5314,
  -41.5794,
  -41.6365,
  -41.6996,
  -41.7719,
  -41.8523,
  -41.9415,
  -42.0362,
  -42.1336,
  -42.228,
  -42.3159,
  -42.3954,
  -42.4642,
  -42.5221,
  -42.5696,
  -42.6074,
  -42.6352,
  -42.6525,
  -42.6593,
  -42.6535,
  -42.6326,
  -42.5942,
  -42.5367,
  -42.458,
  -42.3583,
  -42.238,
  -42.103,
  -41.9572,
  -41.8075,
  -41.661,
  -41.5239,
  -41.401,
  -41.2944,
  -41.2048,
  -41.1316,
  -41.0744,
  -41.0304,
  -40.9977,
  -40.9737,
  -41.1088,
  -41.1444,
  -41.177,
  -41.2076,
  -41.2369,
  -41.2662,
  -41.2963,
  -41.3274,
  -41.3606,
  -41.3957,
  -41.4336,
  -41.4733,
  -41.5171,
  -41.5643,
  -41.6137,
  -41.6648,
  -41.7177,
  -41.7713,
  -41.8257,
  -41.8801,
  -41.9348,
  -41.9903,
  -42.0472,
  -42.1066,
  -42.1686,
  -42.2338,
  -42.3012,
  -42.3724,
  -42.4461,
  -42.5213,
  -42.5962,
  -42.6694,
  -42.7394,
  -42.806,
  -42.8681,
  -42.926,
  -42.9794,
  -43.0284,
  -43.074,
  -43.1155,
  -43.1532,
  -43.1861,
  -43.2169,
  -43.2446,
  -43.2695,
  -43.2921,
  -43.3132,
  -43.333,
  -43.3518,
  -43.3696,
  -43.386,
  -43.4007,
  -43.4124,
  -43.4214,
  -43.4274,
  -43.4291,
  -43.4269,
  -43.4194,
  -43.4095,
  -43.397,
  -43.3821,
  -43.3658,
  -43.3481,
  -43.3298,
  -43.3112,
  -43.2924,
  -43.2745,
  -43.2564,
  -43.2373,
  -43.217,
  -43.1951,
  -43.1728,
  -43.1511,
  -43.1314,
  -43.113,
  -43.0981,
  -43.0856,
  -43.0756,
  -43.068,
  -43.0627,
  -43.0599,
  -43.0595,
  -43.0617,
  -43.0659,
  -43.0713,
  -43.0778,
  -43.085,
  -43.0933,
  -43.1022,
  -43.1107,
  -43.1173,
  -43.1208,
  -43.1198,
  -43.1158,
  -43.1073,
  -43.0938,
  -43.0747,
  -43.0501,
  -43.0192,
  -42.982,
  -42.9387,
  -42.8898,
  -42.8362,
  -42.7799,
  -42.7234,
  -42.6691,
  -42.6204,
  -42.5809,
  -42.5529,
  -42.5387,
  -42.5403,
  -42.5567,
  -42.5875,
  -42.6298,
  -42.6797,
  -42.7338,
  -42.7896,
  -42.8453,
  -42.8997,
  -42.9518,
  -43.0003,
  -43.0451,
  -43.0858,
  -43.1221,
  -43.1535,
  -43.1794,
  -43.2005,
  -43.2177,
  -43.2321,
  -43.2451,
  -43.2566,
  -43.2659,
  -43.275,
  -43.2826,
  -43.2885,
  -43.2916,
  -43.2909,
  -43.2858,
  -43.2769,
  -43.2654,
  -43.2525,
  -43.24,
  -43.2292,
  -43.2206,
  -43.2139,
  -43.208,
  -43.2014,
  -43.1925,
  -43.1799,
  -43.162,
  -43.1383,
  -43.11,
  -43.0789,
  -43.0456,
  -43.013,
  -42.9804,
  -42.9479,
  -42.9156,
  -42.8831,
  -42.8491,
  -42.8131,
  -42.775,
  -42.7351,
  -42.6936,
  -42.6514,
  -42.61,
  -42.5701,
  -42.5331,
  -42.5001,
  -42.4714,
  -42.4461,
  -42.4243,
  -42.4064,
  -42.3922,
  -42.3827,
  -42.3778,
  -42.3767,
  -42.3779,
  -42.3819,
  -42.3863,
  -42.3898,
  -42.3908,
  -42.3887,
  -42.3834,
  -42.3753,
  -42.3657,
  -42.3555,
  -42.3452,
  -42.3351,
  -42.325,
  -42.3146,
  -42.304,
  -42.2939,
  -42.285,
  -42.2785,
  -42.2766,
  -42.2805,
  -42.2923,
  -42.3137,
  -42.3452,
  -42.3861,
  -42.434,
  -42.4857,
  -42.5374,
  -42.5849,
  -42.6268,
  -42.6616,
  -42.6888,
  -42.7097,
  -42.7256,
  -42.7382,
  -42.7487,
  -42.7581,
  -42.7668,
  -42.7744,
  -42.7811,
  -42.7861,
  -42.7889,
  -42.7901,
  -42.7897,
  -42.7892,
  -42.7892,
  -42.7894,
  -42.7889,
  -42.7856,
  -42.7787,
  -42.7663,
  -42.7469,
  -42.7195,
  -42.6852,
  -42.6465,
  -42.6057,
  -42.565,
  -42.5258,
  -42.4863,
  -42.4466,
  -42.4028,
  -42.3506,
  -42.286,
  -42.207,
  -42.1131,
  -42.0062,
  -41.8897,
  -41.77,
  -41.6516,
  -41.5429,
  -41.448,
  -41.3721,
  -41.3146,
  -41.28,
  -41.2656,
  -41.2681,
  -41.2823,
  -41.3053,
  -41.3318,
  -41.3609,
  -41.3929,
  -41.4264,
  -41.4648,
  -41.5021,
  -41.5419,
  -41.5846,
  -41.6312,
  -41.679,
  -41.7334,
  -41.7957,
  -41.863,
  -41.9395,
  -42.0237,
  -42.1137,
  -42.2062,
  -42.2965,
  -42.3802,
  -42.4572,
  -42.524,
  -42.5804,
  -42.6271,
  -42.6638,
  -42.6906,
  -42.7067,
  -42.7117,
  -42.7037,
  -42.68,
  -42.6389,
  -42.5783,
  -42.4971,
  -42.395,
  -42.2734,
  -42.1361,
  -41.9876,
  -41.8342,
  -41.6827,
  -41.5387,
  -41.4071,
  -41.2915,
  -41.1912,
  -41.1078,
  -41.0402,
  -40.9867,
  -40.9447,
  -40.913,
  -41.1444,
  -41.1806,
  -41.2143,
  -41.2465,
  -41.2781,
  -41.3098,
  -41.341,
  -41.3743,
  -41.4091,
  -41.4457,
  -41.4848,
  -41.5265,
  -41.571,
  -41.6182,
  -41.6677,
  -41.7189,
  -41.771,
  -41.8238,
  -41.8769,
  -41.9298,
  -41.9826,
  -42.0348,
  -42.0893,
  -42.1457,
  -42.2047,
  -42.2664,
  -42.331,
  -42.3992,
  -42.4702,
  -42.5424,
  -42.6145,
  -42.6847,
  -42.7515,
  -42.8142,
  -42.8723,
  -42.9263,
  -42.9757,
  -43.0224,
  -43.0658,
  -43.1054,
  -43.1412,
  -43.1734,
  -43.202,
  -43.2278,
  -43.2506,
  -43.2711,
  -43.2897,
  -43.3072,
  -43.3239,
  -43.3396,
  -43.3542,
  -43.3674,
  -43.3776,
  -43.3862,
  -43.3917,
  -43.3931,
  -43.3907,
  -43.3842,
  -43.3741,
  -43.3615,
  -43.3469,
  -43.3309,
  -43.3144,
  -43.2972,
  -43.2799,
  -43.2627,
  -43.2459,
  -43.2291,
  -43.2113,
  -43.1904,
  -43.1693,
  -43.147,
  -43.1249,
  -43.1042,
  -43.0855,
  -43.0695,
  -43.0562,
  -43.046,
  -43.0387,
  -43.0343,
  -43.0328,
  -43.0339,
  -43.0374,
  -43.043,
  -43.0497,
  -43.0574,
  -43.0651,
  -43.0749,
  -43.0857,
  -43.096,
  -43.1048,
  -43.1106,
  -43.1133,
  -43.1122,
  -43.1068,
  -43.0967,
  -43.0809,
  -43.0594,
  -43.0322,
  -42.999,
  -42.9596,
  -42.9149,
  -42.8659,
  -42.8144,
  -42.7624,
  -42.7116,
  -42.6674,
  -42.6325,
  -42.6094,
  -42.6006,
  -42.6079,
  -42.6313,
  -42.6689,
  -42.7178,
  -42.7738,
  -42.8332,
  -42.8933,
  -42.9519,
  -43.0077,
  -43.06,
  -43.1076,
  -43.1509,
  -43.1899,
  -43.2245,
  -43.2532,
  -43.2785,
  -43.2993,
  -43.3167,
  -43.3316,
  -43.3448,
  -43.3562,
  -43.366,
  -43.3746,
  -43.3816,
  -43.3871,
  -43.3905,
  -43.3906,
  -43.3873,
  -43.3806,
  -43.3716,
  -43.3614,
  -43.3513,
  -43.3427,
  -43.336,
  -43.3308,
  -43.325,
  -43.3193,
  -43.3115,
  -43.2996,
  -43.2828,
  -43.261,
  -43.2349,
  -43.2066,
  -43.1778,
  -43.149,
  -43.1204,
  -43.0916,
  -43.063,
  -43.0338,
  -43.0034,
  -42.9708,
  -42.9368,
  -42.9014,
  -42.8643,
  -42.8269,
  -42.7897,
  -42.7538,
  -42.7201,
  -42.6891,
  -42.6601,
  -42.6345,
  -42.6114,
  -42.5909,
  -42.5737,
  -42.5607,
  -42.5519,
  -42.5474,
  -42.5462,
  -42.5474,
  -42.5498,
  -42.5516,
  -42.5516,
  -42.5486,
  -42.542,
  -42.5317,
  -42.5181,
  -42.5021,
  -42.4846,
  -42.4659,
  -42.4464,
  -42.4262,
  -42.406,
  -42.3868,
  -42.3699,
  -42.3548,
  -42.3456,
  -42.344,
  -42.3504,
  -42.3665,
  -42.3922,
  -42.4271,
  -42.4681,
  -42.5126,
  -42.5567,
  -42.5972,
  -42.6316,
  -42.6592,
  -42.68,
  -42.6955,
  -42.7068,
  -42.7152,
  -42.722,
  -42.7277,
  -42.7323,
  -42.7357,
  -42.7384,
  -42.7405,
  -42.7416,
  -42.7416,
  -42.7408,
  -42.74,
  -42.7397,
  -42.7393,
  -42.7368,
  -42.7328,
  -42.7253,
  -42.7125,
  -42.6929,
  -42.6668,
  -42.6353,
  -42.6003,
  -42.5642,
  -42.5285,
  -42.4936,
  -42.4586,
  -42.4214,
  -42.3792,
  -42.3276,
  -42.2635,
  -42.1856,
  -42.0939,
  -41.9906,
  -41.8792,
  -41.765,
  -41.6529,
  -41.5508,
  -41.4639,
  -41.395,
  -41.3446,
  -41.3168,
  -41.3084,
  -41.317,
  -41.3372,
  -41.3658,
  -41.3986,
  -41.4358,
  -41.474,
  -41.5142,
  -41.5556,
  -41.5968,
  -41.6386,
  -41.6823,
  -41.7278,
  -41.7758,
  -41.828,
  -41.8862,
  -41.9509,
  -42.0234,
  -42.1031,
  -42.1885,
  -42.2763,
  -42.3626,
  -42.4446,
  -42.5189,
  -42.5836,
  -42.6389,
  -42.6845,
  -42.7207,
  -42.7464,
  -42.7614,
  -42.765,
  -42.7547,
  -42.7288,
  -42.6854,
  -42.6229,
  -42.5402,
  -42.4374,
  -42.3158,
  -42.1785,
  -42.03,
  -41.8755,
  -41.7209,
  -41.5716,
  -41.4325,
  -41.3073,
  -41.1971,
  -41.1019,
  -41.0229,
  -40.9577,
  -40.9058,
  -40.8648,
  -41.1749,
  -41.2111,
  -41.2461,
  -41.28,
  -41.3136,
  -41.3476,
  -41.3823,
  -41.4179,
  -41.4544,
  -41.4926,
  -41.5327,
  -41.575,
  -41.62,
  -41.6676,
  -41.717,
  -41.7678,
  -41.8182,
  -41.8701,
  -41.9218,
  -41.9731,
  -42.024,
  -42.0753,
  -42.1273,
  -42.1808,
  -42.2367,
  -42.2952,
  -42.3564,
  -42.4211,
  -42.4885,
  -42.5573,
  -42.626,
  -42.6919,
  -42.7554,
  -42.8145,
  -42.8693,
  -42.9201,
  -42.9674,
  -43.0117,
  -43.0532,
  -43.0913,
  -43.1254,
  -43.1558,
  -43.1827,
  -43.2065,
  -43.2275,
  -43.246,
  -43.2615,
  -43.2769,
  -43.2912,
  -43.3049,
  -43.3175,
  -43.329,
  -43.339,
  -43.3467,
  -43.3514,
  -43.3522,
  -43.3496,
  -43.3432,
  -43.3333,
  -43.3211,
  -43.3074,
  -43.2925,
  -43.277,
  -43.2601,
  -43.244,
  -43.2283,
  -43.2123,
  -43.1963,
  -43.1791,
  -43.1601,
  -43.1398,
  -43.118,
  -43.0957,
  -43.0744,
  -43.055,
  -43.0381,
  -43.0244,
  -43.0139,
  -43.007,
  -43.0034,
  -43.0017,
  -43.0041,
  -43.009,
  -43.0156,
  -43.0234,
  -43.0322,
  -43.042,
  -43.0532,
  -43.0653,
  -43.0772,
  -43.0878,
  -43.0962,
  -43.1015,
  -43.1033,
  -43.1008,
  -43.0937,
  -43.0814,
  -43.0637,
  -43.0396,
  -43.0112,
  -42.9773,
  -42.9384,
  -42.8957,
  -42.8502,
  -42.8044,
  -42.7605,
  -42.7218,
  -42.6917,
  -42.6737,
  -42.6702,
  -42.6824,
  -42.7108,
  -42.7534,
  -42.8068,
  -42.8669,
  -42.9298,
  -42.9922,
  -43.051,
  -43.1068,
  -43.1582,
  -43.2044,
  -43.2454,
  -43.2819,
  -43.3143,
  -43.3426,
  -43.3668,
  -43.3873,
  -43.4047,
  -43.4198,
  -43.433,
  -43.4441,
  -43.4535,
  -43.4613,
  -43.4681,
  -43.4736,
  -43.4774,
  -43.4786,
  -43.4771,
  -43.4718,
  -43.4657,
  -43.4582,
  -43.4507,
  -43.4442,
  -43.439,
  -43.4349,
  -43.4309,
  -43.4258,
  -43.4182,
  -43.4068,
  -43.3909,
  -43.3707,
  -43.3471,
  -43.3216,
  -43.2959,
  -43.2708,
  -43.2456,
  -43.2201,
  -43.1947,
  -43.1686,
  -43.1415,
  -43.1128,
  -43.0816,
  -43.0503,
  -43.018,
  -42.9852,
  -42.9526,
  -42.9208,
  -42.8907,
  -42.8623,
  -42.8358,
  -42.8107,
  -42.787,
  -42.765,
  -42.7458,
  -42.7298,
  -42.7178,
  -42.7098,
  -42.7054,
  -42.7036,
  -42.7036,
  -42.7037,
  -42.7022,
  -42.6982,
  -42.6901,
  -42.6781,
  -42.6606,
  -42.6406,
  -42.6179,
  -42.5931,
  -42.5669,
  -42.5397,
  -42.5128,
  -42.4871,
  -42.4637,
  -42.4438,
  -42.4291,
  -42.4214,
  -42.4224,
  -42.433,
  -42.4532,
  -42.4817,
  -42.516,
  -42.5533,
  -42.59,
  -42.6231,
  -42.6505,
  -42.6713,
  -42.6861,
  -42.6961,
  -42.7025,
  -42.7064,
  -42.7085,
  -42.7099,
  -42.7089,
  -42.7086,
  -42.708,
  -42.7076,
  -42.7071,
  -42.7069,
  -42.7063,
  -42.7061,
  -42.706,
  -42.7052,
  -42.7032,
  -42.6987,
  -42.6908,
  -42.6775,
  -42.6583,
  -42.6333,
  -42.6041,
  -42.5725,
  -42.5404,
  -42.5087,
  -42.4774,
  -42.4452,
  -42.4098,
  -42.3686,
  -42.3179,
  -42.2555,
  -42.1797,
  -42.0916,
  -41.9932,
  -41.8882,
  -41.7815,
  -41.6774,
  -41.5824,
  -41.502,
  -41.4397,
  -41.3961,
  -41.3738,
  -41.3696,
  -41.3806,
  -41.4047,
  -41.4366,
  -41.4739,
  -41.5155,
  -41.5592,
  -41.604,
  -41.6497,
  -41.6938,
  -41.7373,
  -41.7805,
  -41.8251,
  -41.8714,
  -41.9227,
  -41.9785,
  -42.0405,
  -42.1094,
  -42.1846,
  -42.2653,
  -42.3485,
  -42.431,
  -42.5092,
  -42.5808,
  -42.6437,
  -42.6976,
  -42.742,
  -42.7768,
  -42.8014,
  -42.8153,
  -42.8173,
  -42.8052,
  -42.7773,
  -42.732,
  -42.6683,
  -42.5854,
  -42.4824,
  -42.3624,
  -42.2272,
  -42.0806,
  -41.927,
  -41.7715,
  -41.6189,
  -41.4738,
  -41.3398,
  -41.2189,
  -41.1124,
  -41.0208,
  -40.9434,
  -40.8794,
  -40.8276,
  -41.1989,
  -41.2372,
  -41.2734,
  -41.3091,
  -41.3451,
  -41.3817,
  -41.4189,
  -41.4567,
  -41.4951,
  -41.5345,
  -41.5753,
  -41.6172,
  -41.6625,
  -41.71,
  -41.7592,
  -41.8093,
  -41.8599,
  -41.9104,
  -41.961,
  -42.0108,
  -42.0601,
  -42.1095,
  -42.1597,
  -42.2107,
  -42.2636,
  -42.3189,
  -42.3762,
  -42.4374,
  -42.5013,
  -42.5665,
  -42.6315,
  -42.6946,
  -42.7545,
  -42.8105,
  -42.8622,
  -42.91,
  -42.9548,
  -42.9967,
  -43.0359,
  -43.072,
  -43.1044,
  -43.1319,
  -43.1571,
  -43.179,
  -43.1986,
  -43.2153,
  -43.2303,
  -43.2437,
  -43.256,
  -43.2676,
  -43.2781,
  -43.2876,
  -43.2959,
  -43.3021,
  -43.3058,
  -43.306,
  -43.303,
  -43.2957,
  -43.2865,
  -43.2753,
  -43.2629,
  -43.2494,
  -43.2351,
  -43.2204,
  -43.2054,
  -43.1901,
  -43.1744,
  -43.1586,
  -43.142,
  -43.1241,
  -43.1044,
  -43.0839,
  -43.0623,
  -43.0413,
  -43.0208,
  -43.0039,
  -42.9902,
  -42.98,
  -42.9735,
  -42.9707,
  -42.9711,
  -42.9744,
  -42.9799,
  -42.9873,
  -42.9959,
  -43.0059,
  -43.0169,
  -43.029,
  -43.0421,
  -43.0555,
  -43.0679,
  -43.0784,
  -43.0855,
  -43.09,
  -43.0906,
  -43.0862,
  -43.077,
  -43.063,
  -43.0446,
  -43.0218,
  -42.9945,
  -42.9628,
  -42.9275,
  -42.8898,
  -42.8516,
  -42.8145,
  -42.7818,
  -42.757,
  -42.7438,
  -42.745,
  -42.7614,
  -42.7919,
  -42.8374,
  -42.8931,
  -42.9552,
  -43.0194,
  -43.0823,
  -43.142,
  -43.197,
  -43.2467,
  -43.2908,
  -43.3295,
  -43.3634,
  -43.3935,
  -43.4203,
  -43.4436,
  -43.4639,
  -43.4815,
  -43.4968,
  -43.5098,
  -43.5207,
  -43.5286,
  -43.5361,
  -43.5424,
  -43.5479,
  -43.5521,
  -43.5545,
  -43.5547,
  -43.553,
  -43.5496,
  -43.545,
  -43.5398,
  -43.5351,
  -43.5312,
  -43.5279,
  -43.5241,
  -43.5189,
  -43.5112,
  -43.5001,
  -43.485,
  -43.4663,
  -43.445,
  -43.4225,
  -43.3989,
  -43.3767,
  -43.3547,
  -43.3323,
  -43.3094,
  -43.2859,
  -43.2616,
  -43.2364,
  -43.2098,
  -43.1825,
  -43.1546,
  -43.1264,
  -43.0984,
  -43.071,
  -43.0445,
  -43.0193,
  -42.9951,
  -42.9713,
  -42.9481,
  -42.9258,
  -42.9053,
  -42.8873,
  -42.8729,
  -42.8619,
  -42.8535,
  -42.8491,
  -42.8465,
  -42.8447,
  -42.8419,
  -42.8366,
  -42.8276,
  -42.8144,
  -42.7965,
  -42.7742,
  -42.7487,
  -42.7204,
  -42.6901,
  -42.659,
  -42.6282,
  -42.5985,
  -42.5706,
  -42.546,
  -42.5264,
  -42.5132,
  -42.5084,
  -42.5132,
  -42.5272,
  -42.5488,
  -42.5761,
  -42.606,
  -42.6343,
  -42.6604,
  -42.6811,
  -42.6955,
  -42.7042,
  -42.7085,
  -42.7098,
  -42.7091,
  -42.7072,
  -42.704,
  -42.6999,
  -42.6957,
  -42.6923,
  -42.6904,
  -42.6894,
  -42.6894,
  -42.6904,
  -42.6913,
  -42.6919,
  -42.6913,
  -42.6891,
  -42.6845,
  -42.6758,
  -42.6624,
  -42.643,
  -42.6186,
  -42.5913,
  -42.5624,
  -42.5334,
  -42.5046,
  -42.4758,
  -42.4442,
  -42.41,
  -42.3695,
  -42.3199,
  -42.2595,
  -42.187,
  -42.1041,
  -42.0124,
  -41.9152,
  -41.8171,
  -41.7232,
  -41.6379,
  -41.5655,
  -41.5101,
  -41.4718,
  -41.4533,
  -41.4521,
  -41.4651,
  -41.49,
  -41.5232,
  -41.563,
  -41.608,
  -41.6543,
  -41.7007,
  -41.7482,
  -41.7938,
  -41.8377,
  -41.8806,
  -41.9241,
  -41.969,
  -42.0181,
  -42.0722,
  -42.1318,
  -42.1975,
  -42.2692,
  -42.3453,
  -42.4241,
  -42.5011,
  -42.5756,
  -42.6436,
  -42.704,
  -42.7557,
  -42.7983,
  -42.8314,
  -42.8543,
  -42.867,
  -42.867,
  -42.853,
  -42.823,
  -42.7761,
  -42.7118,
  -42.6295,
  -42.5294,
  -42.4126,
  -42.2812,
  -42.1384,
  -41.9879,
  -41.8334,
  -41.6794,
  -41.5296,
  -41.3878,
  -41.2568,
  -41.1384,
  -41.0339,
  -40.9432,
  -40.8662,
  -40.8025,
  -41.2191,
  -41.2585,
  -41.2966,
  -41.334,
  -41.3721,
  -41.4109,
  -41.4492,
  -41.489,
  -41.5288,
  -41.5692,
  -41.6108,
  -41.6543,
  -41.7,
  -41.7475,
  -41.7963,
  -41.8456,
  -41.8953,
  -41.9449,
  -41.9934,
  -42.042,
  -42.0902,
  -42.1372,
  -42.1848,
  -42.2337,
  -42.2843,
  -42.3368,
  -42.3921,
  -42.4503,
  -42.5105,
  -42.5721,
  -42.6332,
  -42.6928,
  -42.7493,
  -42.8023,
  -42.8514,
  -42.8967,
  -42.9378,
  -42.9768,
  -43.0133,
  -43.047,
  -43.0773,
  -43.1039,
  -43.1273,
  -43.1477,
  -43.1657,
  -43.181,
  -43.1948,
  -43.2066,
  -43.2172,
  -43.2267,
  -43.2352,
  -43.2424,
  -43.2478,
  -43.2525,
  -43.2548,
  -43.2543,
  -43.2509,
  -43.2446,
  -43.2363,
  -43.2261,
  -43.2147,
  -43.2024,
  -43.1893,
  -43.1755,
  -43.1611,
  -43.1463,
  -43.1312,
  -43.1155,
  -43.0984,
  -43.0811,
  -43.0628,
  -43.0434,
  -43.0235,
  -43.0037,
  -42.9853,
  -42.9691,
  -42.9562,
  -42.9468,
  -42.9413,
  -42.9396,
  -42.941,
  -42.9451,
  -42.9515,
  -42.9597,
  -42.9692,
  -42.98,
  -42.9907,
  -43.0037,
  -43.0175,
  -43.032,
  -43.0459,
  -43.0586,
  -43.0689,
  -43.0759,
  -43.0788,
  -43.0772,
  -43.0711,
  -43.0612,
  -43.0477,
  -43.031,
  -43.0108,
  -42.987,
  -42.9601,
  -42.931,
  -42.8998,
  -42.8703,
  -42.8441,
  -42.8251,
  -42.8168,
  -42.8219,
  -42.8409,
  -42.8742,
  -42.9206,
  -42.9766,
  -43.0385,
  -43.1021,
  -43.1642,
  -43.2225,
  -43.276,
  -43.3239,
  -43.3659,
  -43.4022,
  -43.434,
  -43.4624,
  -43.4868,
  -43.5096,
  -43.5299,
  -43.5477,
  -43.5632,
  -43.5764,
  -43.5872,
  -43.5957,
  -43.6028,
  -43.609,
  -43.6146,
  -43.6194,
  -43.623,
  -43.6251,
  -43.6256,
  -43.6246,
  -43.6222,
  -43.6191,
  -43.6158,
  -43.6125,
  -43.6092,
  -43.604,
  -43.5983,
  -43.5903,
  -43.5791,
  -43.5652,
  -43.5483,
  -43.5293,
  -43.5095,
  -43.4898,
  -43.4704,
  -43.4513,
  -43.4314,
  -43.411,
  -43.3898,
  -43.3681,
  -43.3456,
  -43.3227,
  -43.299,
  -43.2752,
  -43.2513,
  -43.2274,
  -43.204,
  -43.1813,
  -43.1583,
  -43.1369,
  -43.1149,
  -43.0931,
  -43.0712,
  -43.0505,
  -43.0315,
  -43.0156,
  -43.0029,
  -42.9938,
  -42.9872,
  -42.9822,
  -42.9782,
  -42.9737,
  -42.967,
  -42.957,
  -42.9431,
  -42.9247,
  -42.9018,
  -42.8752,
  -42.8455,
  -42.814,
  -42.7813,
  -42.7488,
  -42.7171,
  -42.6867,
  -42.6579,
  -42.6342,
  -42.6163,
  -42.6061,
  -42.6046,
  -42.6116,
  -42.626,
  -42.6456,
  -42.668,
  -42.69,
  -42.7092,
  -42.7234,
  -42.7319,
  -42.7352,
  -42.7345,
  -42.731,
  -42.726,
  -42.72,
  -42.7132,
  -42.7058,
  -42.6987,
  -42.6931,
  -42.6899,
  -42.6888,
  -42.69,
  -42.6923,
  -42.6947,
  -42.6961,
  -42.6962,
  -42.693,
  -42.6878,
  -42.6786,
  -42.6644,
  -42.6453,
  -42.6215,
  -42.595,
  -42.5671,
  -42.5399,
  -42.5134,
  -42.4862,
  -42.4567,
  -42.4236,
  -42.3842,
  -42.3363,
  -42.2785,
  -42.21,
  -42.1325,
  -42.0482,
  -41.9597,
  -41.8715,
  -41.7872,
  -41.7116,
  -41.6481,
  -41.5992,
  -41.5662,
  -41.5503,
  -41.5504,
  -41.5644,
  -41.5895,
  -41.6227,
  -41.6633,
  -41.7082,
  -41.7557,
  -41.8029,
  -41.851,
  -41.8967,
  -41.9409,
  -41.9834,
  -42.0256,
  -42.0695,
  -42.1169,
  -42.1691,
  -42.2261,
  -42.2885,
  -42.3562,
  -42.428,
  -42.5013,
  -42.5747,
  -42.6446,
  -42.7086,
  -42.7656,
  -42.8145,
  -42.8547,
  -42.8855,
  -42.9064,
  -42.9172,
  -42.9151,
  -42.8985,
  -42.8666,
  -42.8186,
  -42.7541,
  -42.6727,
  -42.5753,
  -42.4624,
  -42.3358,
  -42.198,
  -42.0517,
  -41.9001,
  -41.7464,
  -41.5935,
  -41.4456,
  -41.3053,
  -41.176,
  -41.0591,
  -40.9551,
  -40.8649,
  -40.7886,
  -41.2351,
  -41.275,
  -41.3145,
  -41.3539,
  -41.3939,
  -41.4345,
  -41.4754,
  -41.5166,
  -41.5576,
  -41.5989,
  -41.6413,
  -41.6852,
  -41.731,
  -41.7786,
  -41.8268,
  -41.8759,
  -41.9235,
  -41.9717,
  -42.0191,
  -42.0664,
  -42.1131,
  -42.1593,
  -42.2054,
  -42.2526,
  -42.3008,
  -42.351,
  -42.4037,
  -42.4588,
  -42.5156,
  -42.5733,
  -42.6309,
  -42.6859,
  -42.7396,
  -42.7899,
  -42.8362,
  -42.8787,
  -42.9178,
  -42.9541,
  -42.9879,
  -43.019,
  -43.047,
  -43.0713,
  -43.0928,
  -43.1117,
  -43.1278,
  -43.1421,
  -43.1537,
  -43.1643,
  -43.1734,
  -43.1811,
  -43.1874,
  -43.1926,
  -43.197,
  -43.2,
  -43.2007,
  -43.1992,
  -43.1952,
  -43.1893,
  -43.1817,
  -43.1725,
  -43.1621,
  -43.1507,
  -43.1383,
  -43.1242,
  -43.1105,
  -43.096,
  -43.0812,
  -43.0656,
  -43.0501,
  -43.0341,
  -43.0173,
  -42.9997,
  -42.9818,
  -42.964,
  -42.9476,
  -42.9331,
  -42.9216,
  -42.9139,
  -42.9096,
  -42.909,
  -42.9105,
  -42.9159,
  -42.9234,
  -42.9324,
  -42.9431,
  -42.9547,
  -42.9671,
  -42.9804,
  -42.9949,
  -43.01,
  -43.0253,
  -43.0396,
  -43.0518,
  -43.0606,
  -43.0657,
  -43.0666,
  -43.0638,
  -43.058,
  -43.0487,
  -43.0381,
  -43.025,
  -43.0091,
  -42.9908,
  -42.9704,
  -42.9483,
  -42.9268,
  -42.9079,
  -42.8947,
  -42.8907,
  -42.8987,
  -42.92,
  -42.9534,
  -42.9985,
  -43.0529,
  -43.113,
  -43.1748,
  -43.2349,
  -43.2903,
  -43.3417,
  -43.3875,
  -43.4274,
  -43.4621,
  -43.4924,
  -43.5194,
  -43.5441,
  -43.5667,
  -43.5872,
  -43.6055,
  -43.6214,
  -43.6348,
  -43.6456,
  -43.6542,
  -43.6613,
  -43.6675,
  -43.6736,
  -43.6791,
  -43.6838,
  -43.6875,
  -43.6887,
  -43.6897,
  -43.6892,
  -43.6875,
  -43.6849,
  -43.6817,
  -43.6778,
  -43.6728,
  -43.6663,
  -43.6578,
  -43.647,
  -43.6343,
  -43.6193,
  -43.6028,
  -43.5856,
  -43.5687,
  -43.552,
  -43.5352,
  -43.5177,
  -43.4997,
  -43.4808,
  -43.4615,
  -43.4406,
  -43.4205,
  -43.4003,
  -43.3798,
  -43.3597,
  -43.3398,
  -43.3203,
  -43.3013,
  -43.2827,
  -43.2639,
  -43.2446,
  -43.2246,
  -43.2041,
  -43.1838,
  -43.1652,
  -43.1487,
  -43.1353,
  -43.1245,
  -43.1167,
  -43.1103,
  -43.1043,
  -43.0977,
  -43.0895,
  -43.0788,
  -43.0645,
  -43.045,
  -43.0225,
  -42.9965,
  -42.9671,
  -42.9365,
  -42.9041,
  -42.8719,
  -42.8398,
  -42.8084,
  -42.7786,
  -42.752,
  -42.7299,
  -42.7146,
  -42.7068,
  -42.7067,
  -42.7131,
  -42.725,
  -42.7394,
  -42.754,
  -42.7663,
  -42.7745,
  -42.7777,
  -42.7762,
  -42.7714,
  -42.764,
  -42.7556,
  -42.7463,
  -42.7355,
  -42.7255,
  -42.7166,
  -42.7098,
  -42.7056,
  -42.705,
  -42.7071,
  -42.7104,
  -42.7142,
  -42.7161,
  -42.7169,
  -42.7145,
  -42.709,
  -42.6991,
  -42.6841,
  -42.6642,
  -42.6402,
  -42.6136,
  -42.5867,
  -42.5604,
  -42.5348,
  -42.5086,
  -42.4805,
  -42.4485,
  -42.4106,
  -42.3651,
  -42.3103,
  -42.2465,
  -42.1751,
  -42.0984,
  -42.0189,
  -41.9407,
  -41.867,
  -41.8003,
  -41.7452,
  -41.7032,
  -41.675,
  -41.6614,
  -41.6622,
  -41.6761,
  -41.7001,
  -41.7324,
  -41.7721,
  -41.8165,
  -41.8636,
  -41.9117,
  -41.9594,
  -42.0049,
  -42.0487,
  -42.0903,
  -42.1313,
  -42.1741,
  -42.2199,
  -42.2705,
  -42.3247,
  -42.3838,
  -42.4477,
  -42.5141,
  -42.5822,
  -42.6499,
  -42.7146,
  -42.7741,
  -42.827,
  -42.8727,
  -42.9096,
  -42.9372,
  -42.9559,
  -42.9636,
  -42.9592,
  -42.9406,
  -42.9067,
  -42.8578,
  -42.7933,
  -42.7133,
  -42.6175,
  -42.5086,
  -42.3868,
  -42.2543,
  -42.1129,
  -41.9648,
  -41.8125,
  -41.6588,
  -41.506,
  -41.3589,
  -41.2206,
  -41.0919,
  -40.9755,
  -40.8725,
  -40.7837,
  -41.2463,
  -41.289,
  -41.3304,
  -41.3714,
  -41.413,
  -41.4548,
  -41.4971,
  -41.5392,
  -41.5809,
  -41.6229,
  -41.6656,
  -41.7087,
  -41.7545,
  -41.8018,
  -41.8497,
  -41.8978,
  -41.9456,
  -41.9927,
  -42.0391,
  -42.085,
  -42.1304,
  -42.1753,
  -42.2202,
  -42.2655,
  -42.312,
  -42.3602,
  -42.4096,
  -42.4618,
  -42.5155,
  -42.5696,
  -42.6239,
  -42.6768,
  -42.7273,
  -42.775,
  -42.8186,
  -42.8584,
  -42.8948,
  -42.928,
  -42.9588,
  -42.9868,
  -43.0121,
  -43.0332,
  -43.0526,
  -43.0696,
  -43.0841,
  -43.0973,
  -43.1086,
  -43.1185,
  -43.1264,
  -43.1326,
  -43.1373,
  -43.1407,
  -43.1429,
  -43.1438,
  -43.1433,
  -43.1405,
  -43.1362,
  -43.1294,
  -43.1223,
  -43.1137,
  -43.1039,
  -43.093,
  -43.0813,
  -43.0687,
  -43.0554,
  -43.0413,
  -43.0269,
  -43.0121,
  -42.9971,
  -42.9825,
  -42.9675,
  -42.9522,
  -42.9368,
  -42.9219,
  -42.9069,
  -42.8949,
  -42.8855,
  -42.8796,
  -42.877,
  -42.8778,
  -42.8819,
  -42.8887,
  -42.8975,
  -42.9079,
  -42.9195,
  -42.932,
  -42.9451,
  -42.959,
  -42.9738,
  -42.9897,
  -43.006,
  -43.0214,
  -43.034,
  -43.0445,
  -43.0513,
  -43.0546,
  -43.055,
  -43.0533,
  -43.05,
  -43.0453,
  -43.0389,
  -43.0307,
  -43.0205,
  -43.0083,
  -42.9946,
  -42.9808,
  -42.969,
  -42.9616,
  -42.9617,
  -42.9721,
  -42.9936,
  -43.0254,
  -43.0684,
  -43.1198,
  -43.1768,
  -43.2355,
  -43.2928,
  -43.3467,
  -43.3958,
  -43.4396,
  -43.4781,
  -43.5113,
  -43.5408,
  -43.5673,
  -43.5916,
  -43.6144,
  -43.6354,
  -43.6542,
  -43.6706,
  -43.6844,
  -43.6956,
  -43.7034,
  -43.7108,
  -43.7174,
  -43.7239,
  -43.7302,
  -43.736,
  -43.741,
  -43.7448,
  -43.7473,
  -43.7483,
  -43.7472,
  -43.7449,
  -43.7413,
  -43.7367,
  -43.7305,
  -43.723,
  -43.7141,
  -43.7039,
  -43.6924,
  -43.6795,
  -43.6655,
  -43.6501,
  -43.6358,
  -43.6216,
  -43.6073,
  -43.5923,
  -43.5765,
  -43.56,
  -43.5429,
  -43.5257,
  -43.5079,
  -43.4904,
  -43.4732,
  -43.4564,
  -43.4401,
  -43.4241,
  -43.4085,
  -43.3931,
  -43.3773,
  -43.3605,
  -43.3427,
  -43.3238,
  -43.3051,
  -43.2874,
  -43.2715,
  -43.257,
  -43.246,
  -43.237,
  -43.2294,
  -43.2218,
  -43.2135,
  -43.2038,
  -43.192,
  -43.1775,
  -43.1594,
  -43.1379,
  -43.1134,
  -43.0859,
  -43.057,
  -43.0267,
  -42.9956,
  -42.9643,
  -42.9331,
  -42.9027,
  -42.874,
  -42.8488,
  -42.8289,
  -42.8152,
  -42.808,
  -42.8068,
  -42.8104,
  -42.8172,
  -42.8236,
  -42.8291,
  -42.8317,
  -42.8301,
  -42.8248,
  -42.8166,
  -42.8065,
  -42.7954,
  -42.7839,
  -42.7722,
  -42.7609,
  -42.7508,
  -42.7433,
  -42.7394,
  -42.7387,
  -42.7411,
  -42.7451,
  -42.7495,
  -42.7525,
  -42.7533,
  -42.7512,
  -42.7447,
  -42.7335,
  -42.7174,
  -42.6963,
  -42.6716,
  -42.6448,
  -42.6176,
  -42.5915,
  -42.5662,
  -42.5399,
  -42.5128,
  -42.4824,
  -42.4467,
  -42.4039,
  -42.353,
  -42.2942,
  -42.2293,
  -42.1602,
  -42.0896,
  -42.0211,
  -41.9574,
  -41.9014,
  -41.8547,
  -41.8191,
  -41.7957,
  -41.7847,
  -41.7857,
  -41.7989,
  -41.8216,
  -41.8526,
  -41.8911,
  -41.9345,
  -41.9805,
  -42.0277,
  -42.0745,
  -42.1192,
  -42.1615,
  -42.2019,
  -42.2418,
  -42.2823,
  -42.3258,
  -42.3734,
  -42.4253,
  -42.4805,
  -42.5393,
  -42.6004,
  -42.6619,
  -42.7238,
  -42.7828,
  -42.8373,
  -42.8856,
  -42.9268,
  -42.9599,
  -42.9846,
  -43,
  -43.005,
  -42.9979,
  -42.9771,
  -42.9418,
  -42.8919,
  -42.8273,
  -42.7483,
  -42.6559,
  -42.5505,
  -42.4335,
  -42.3057,
  -42.169,
  -42.0248,
  -41.875,
  -41.7214,
  -41.567,
  -41.4153,
  -41.2697,
  -41.132,
  -41.0051,
  -40.8905,
  -40.7899,
  -41.2552,
  -41.2999,
  -41.3432,
  -41.386,
  -41.429,
  -41.4721,
  -41.514,
  -41.5565,
  -41.5986,
  -41.6409,
  -41.6837,
  -41.7277,
  -41.7734,
  -41.82,
  -41.8675,
  -41.9148,
  -41.9617,
  -42.0079,
  -42.0533,
  -42.0983,
  -42.1415,
  -42.1854,
  -42.2292,
  -42.273,
  -42.3175,
  -42.3639,
  -42.4119,
  -42.4615,
  -42.5123,
  -42.5634,
  -42.6142,
  -42.664,
  -42.7117,
  -42.7566,
  -42.7978,
  -42.8347,
  -42.8673,
  -42.8976,
  -42.9253,
  -42.95,
  -42.9723,
  -42.992,
  -43.0091,
  -43.0242,
  -43.0373,
  -43.0493,
  -43.0596,
  -43.0685,
  -43.0756,
  -43.0809,
  -43.0843,
  -43.086,
  -43.0851,
  -43.0841,
  -43.0818,
  -43.0779,
  -43.073,
  -43.067,
  -43.0602,
  -43.0521,
  -43.0425,
  -43.0317,
  -43.0207,
  -43.0086,
  -42.9957,
  -42.9822,
  -42.9685,
  -42.9549,
  -42.9402,
  -42.9271,
  -42.9141,
  -42.9014,
  -42.8888,
  -42.8771,
  -42.866,
  -42.8567,
  -42.8497,
  -42.8457,
  -42.845,
  -42.8478,
  -42.8534,
  -42.8618,
  -42.8725,
  -42.8844,
  -42.8975,
  -42.9112,
  -42.9239,
  -42.9384,
  -42.954,
  -42.9703,
  -42.9871,
  -43.0036,
  -43.0181,
  -43.0296,
  -43.038,
  -43.0435,
  -43.0468,
  -43.049,
  -43.0506,
  -43.0511,
  -43.0508,
  -43.0493,
  -43.0463,
  -43.0415,
  -43.0346,
  -43.0284,
  -43.0234,
  -43.0217,
  -43.0258,
  -43.0378,
  -43.0593,
  -43.0904,
  -43.1306,
  -43.1785,
  -43.2316,
  -43.2866,
  -43.3405,
  -43.3915,
  -43.4383,
  -43.4804,
  -43.5173,
  -43.5501,
  -43.5789,
  -43.6055,
  -43.629,
  -43.6521,
  -43.6735,
  -43.6928,
  -43.7099,
  -43.7243,
  -43.7358,
  -43.7452,
  -43.7534,
  -43.7607,
  -43.768,
  -43.775,
  -43.7816,
  -43.7876,
  -43.7926,
  -43.7961,
  -43.7979,
  -43.7975,
  -43.795,
  -43.7909,
  -43.7853,
  -43.7771,
  -43.7688,
  -43.7598,
  -43.7501,
  -43.74,
  -43.7295,
  -43.7183,
  -43.7066,
  -43.6949,
  -43.6832,
  -43.6713,
  -43.6587,
  -43.6453,
  -43.6312,
  -43.6161,
  -43.6008,
  -43.5857,
  -43.5706,
  -43.5562,
  -43.5425,
  -43.5293,
  -43.5164,
  -43.504,
  -43.4906,
  -43.4774,
  -43.4633,
  -43.4475,
  -43.4309,
  -43.4139,
  -43.3979,
  -43.3831,
  -43.3704,
  -43.3595,
  -43.35,
  -43.3416,
  -43.3327,
  -43.3229,
  -43.312,
  -43.2992,
  -43.2844,
  -43.2669,
  -43.2466,
  -43.2238,
  -43.1987,
  -43.1718,
  -43.1442,
  -43.1154,
  -43.0855,
  -43.0544,
  -43.0237,
  -42.9939,
  -42.9668,
  -42.9432,
  -42.9244,
  -42.9111,
  -42.9028,
  -42.8989,
  -42.8981,
  -42.8985,
  -42.898,
  -42.8952,
  -42.8899,
  -42.8817,
  -42.8712,
  -42.8592,
  -42.8467,
  -42.8337,
  -42.8209,
  -42.8092,
  -42.7993,
  -42.7915,
  -42.7877,
  -42.7868,
  -42.7891,
  -42.7931,
  -42.7973,
  -42.8004,
  -42.8001,
  -42.7971,
  -42.7895,
  -42.7769,
  -42.7595,
  -42.7373,
  -42.7116,
  -42.6841,
  -42.6563,
  -42.6298,
  -42.6047,
  -42.5802,
  -42.5545,
  -42.526,
  -42.4929,
  -42.4532,
  -42.4066,
  -42.3533,
  -42.2948,
  -42.2332,
  -42.1713,
  -42.1118,
  -42.0572,
  -42.0101,
  -41.972,
  -41.9429,
  -41.9235,
  -41.915,
  -41.9169,
  -41.9287,
  -41.9488,
  -41.9789,
  -42.0146,
  -42.0556,
  -42.0997,
  -42.144,
  -42.1889,
  -42.2321,
  -42.2733,
  -42.3123,
  -42.3506,
  -42.3893,
  -42.4301,
  -42.4747,
  -42.523,
  -42.574,
  -42.6279,
  -42.6834,
  -42.7399,
  -42.7958,
  -42.8489,
  -42.8978,
  -42.9412,
  -42.9776,
  -43.0068,
  -43.0283,
  -43.0406,
  -43.0427,
  -43.033,
  -43.0103,
  -42.9738,
  -42.9231,
  -42.8585,
  -42.7801,
  -42.6892,
  -42.5862,
  -42.4723,
  -42.3483,
  -42.2155,
  -42.075,
  -41.9285,
  -41.7768,
  -41.6228,
  -41.4693,
  -41.3198,
  -41.1758,
  -41.0409,
  -40.9168,
  -40.8057,
  -41.2611,
  -41.3067,
  -41.352,
  -41.3968,
  -41.4411,
  -41.4851,
  -41.5286,
  -41.5715,
  -41.614,
  -41.6564,
  -41.6992,
  -41.743,
  -41.7879,
  -41.8339,
  -41.8805,
  -41.9261,
  -41.9723,
  -42.0175,
  -42.0619,
  -42.1058,
  -42.1489,
  -42.1918,
  -42.2346,
  -42.2771,
  -42.3202,
  -42.3645,
  -42.4102,
  -42.4573,
  -42.5051,
  -42.5532,
  -42.6,
  -42.6468,
  -42.6917,
  -42.7338,
  -42.772,
  -42.8065,
  -42.8372,
  -42.8648,
  -42.8895,
  -42.9119,
  -42.931,
  -42.948,
  -42.9627,
  -42.9758,
  -42.9875,
  -42.9979,
  -43.0062,
  -43.0143,
  -43.0206,
  -43.0252,
  -43.0276,
  -43.0279,
  -43.0266,
  -43.0237,
  -43.0198,
  -43.0149,
  -43.009,
  -43.0025,
  -42.9951,
  -42.9871,
  -42.9779,
  -42.9674,
  -42.9556,
  -42.944,
  -42.932,
  -42.9196,
  -42.9072,
  -42.8949,
  -42.8831,
  -42.8721,
  -42.8616,
  -42.8515,
  -42.8419,
  -42.8327,
  -42.8247,
  -42.818,
  -42.8134,
  -42.8116,
  -42.813,
  -42.8177,
  -42.8242,
  -42.8344,
  -42.8469,
  -42.8605,
  -42.8749,
  -42.8897,
  -42.9047,
  -42.9202,
  -42.9367,
  -42.9536,
  -42.9711,
  -42.9879,
  -43.0027,
  -43.0151,
  -43.0249,
  -43.0323,
  -43.0386,
  -43.0441,
  -43.0487,
  -43.0538,
  -43.0585,
  -43.0628,
  -43.0661,
  -43.0677,
  -43.0689,
  -43.0698,
  -43.0711,
  -43.0745,
  -43.0824,
  -43.096,
  -43.1172,
  -43.1465,
  -43.1839,
  -43.2279,
  -43.2766,
  -43.3275,
  -43.3779,
  -43.4248,
  -43.4692,
  -43.5095,
  -43.5457,
  -43.5781,
  -43.6073,
  -43.6339,
  -43.6589,
  -43.6825,
  -43.7043,
  -43.7241,
  -43.7415,
  -43.7564,
  -43.7686,
  -43.7789,
  -43.7878,
  -43.796,
  -43.804,
  -43.8117,
  -43.8191,
  -43.8258,
  -43.8305,
  -43.8348,
  -43.8371,
  -43.8369,
  -43.8344,
  -43.8297,
  -43.8234,
  -43.8154,
  -43.8067,
  -43.7978,
  -43.7892,
  -43.7808,
  -43.7724,
  -43.7638,
  -43.7549,
  -43.7459,
  -43.7369,
  -43.7273,
  -43.717,
  -43.7058,
  -43.6937,
  -43.6808,
  -43.6665,
  -43.6535,
  -43.6409,
  -43.629,
  -43.6178,
  -43.6074,
  -43.5972,
  -43.5877,
  -43.578,
  -43.5674,
  -43.5555,
  -43.542,
  -43.5275,
  -43.5128,
  -43.4988,
  -43.4858,
  -43.4741,
  -43.4637,
  -43.4542,
  -43.4452,
  -43.4356,
  -43.4249,
  -43.4129,
  -43.3994,
  -43.3834,
  -43.3663,
  -43.3468,
  -43.3253,
  -43.3023,
  -43.2784,
  -43.253,
  -43.2267,
  -43.199,
  -43.1699,
  -43.14,
  -43.1099,
  -43.0812,
  -43.0551,
  -43.0326,
  -43.0142,
  -43,
  -42.9896,
  -42.9821,
  -42.9763,
  -42.9705,
  -42.9637,
  -42.9551,
  -42.9446,
  -42.9324,
  -42.9196,
  -42.906,
  -42.8929,
  -42.8791,
  -42.8676,
  -42.8582,
  -42.8506,
  -42.8464,
  -42.8451,
  -42.8463,
  -42.8492,
  -42.8523,
  -42.855,
  -42.8545,
  -42.8505,
  -42.8418,
  -42.8279,
  -42.809,
  -42.7855,
  -42.7591,
  -42.7308,
  -42.7028,
  -42.6762,
  -42.6513,
  -42.6275,
  -42.6033,
  -42.5769,
  -42.5463,
  -42.5103,
  -42.4681,
  -42.4202,
  -42.368,
  -42.3137,
  -42.2598,
  -42.209,
  -42.1622,
  -42.1231,
  -42.092,
  -42.0694,
  -42.0546,
  -42.0481,
  -42.0501,
  -42.0608,
  -42.0799,
  -42.1069,
  -42.14,
  -42.178,
  -42.2193,
  -42.2618,
  -42.3044,
  -42.3454,
  -42.3845,
  -42.422,
  -42.4578,
  -42.4939,
  -42.5323,
  -42.5731,
  -42.6168,
  -42.6635,
  -42.712,
  -42.7621,
  -42.8127,
  -42.8629,
  -42.91,
  -42.9536,
  -42.9914,
  -43.0232,
  -43.0484,
  -43.0666,
  -43.076,
  -43.0755,
  -43.0638,
  -43.0395,
  -43.0018,
  -42.9504,
  -42.8853,
  -42.8062,
  -42.7158,
  -42.6138,
  -42.5016,
  -42.3799,
  -42.2499,
  -42.1124,
  -41.9689,
  -41.8206,
  -41.6691,
  -41.5167,
  -41.366,
  -41.2195,
  -41.0797,
  -40.9492,
  -40.8299,
  -41.2633,
  -41.3115,
  -41.3586,
  -41.4052,
  -41.4508,
  -41.4958,
  -41.5399,
  -41.5835,
  -41.6264,
  -41.669,
  -41.7118,
  -41.7542,
  -41.7984,
  -41.8435,
  -41.8893,
  -41.935,
  -41.98,
  -42.0245,
  -42.0676,
  -42.1107,
  -42.1529,
  -42.1948,
  -42.2362,
  -42.2775,
  -42.3192,
  -42.3608,
  -42.4043,
  -42.4487,
  -42.4935,
  -42.5386,
  -42.5834,
  -42.6274,
  -42.6694,
  -42.7085,
  -42.7442,
  -42.7763,
  -42.8048,
  -42.8301,
  -42.8522,
  -42.8713,
  -42.8879,
  -42.901,
  -42.9137,
  -42.9247,
  -42.9346,
  -42.9435,
  -42.9517,
  -42.9589,
  -42.9646,
  -42.9686,
  -42.9702,
  -42.9696,
  -42.9671,
  -42.9628,
  -42.9573,
  -42.9512,
  -42.9442,
  -42.9358,
  -42.9279,
  -42.9195,
  -42.9101,
  -42.8997,
  -42.8893,
  -42.8788,
  -42.8681,
  -42.8572,
  -42.8467,
  -42.8367,
  -42.8275,
  -42.8188,
  -42.8106,
  -42.8032,
  -42.7965,
  -42.79,
  -42.7834,
  -42.7793,
  -42.7768,
  -42.777,
  -42.7804,
  -42.7867,
  -42.7963,
  -42.8084,
  -42.8225,
  -42.8375,
  -42.8533,
  -42.8694,
  -42.8861,
  -42.903,
  -42.9203,
  -42.9382,
  -42.9561,
  -42.9718,
  -42.9869,
  -43.0001,
  -43.011,
  -43.0204,
  -43.0291,
  -43.0376,
  -43.0464,
  -43.0554,
  -43.0644,
  -43.0731,
  -43.0815,
  -43.0892,
  -43.0962,
  -43.1032,
  -43.1101,
  -43.1183,
  -43.1296,
  -43.145,
  -43.1648,
  -43.1925,
  -43.2272,
  -43.2677,
  -43.3123,
  -43.359,
  -43.4055,
  -43.4505,
  -43.4928,
  -43.5314,
  -43.5668,
  -43.599,
  -43.6286,
  -43.6559,
  -43.6816,
  -43.7052,
  -43.7273,
  -43.7473,
  -43.7651,
  -43.7804,
  -43.7924,
  -43.8034,
  -43.8132,
  -43.8224,
  -43.8312,
  -43.8396,
  -43.8475,
  -43.8549,
  -43.8612,
  -43.866,
  -43.8686,
  -43.8685,
  -43.866,
  -43.8612,
  -43.8544,
  -43.8464,
  -43.8376,
  -43.8293,
  -43.8218,
  -43.815,
  -43.8089,
  -43.8028,
  -43.7958,
  -43.7896,
  -43.7831,
  -43.7757,
  -43.7676,
  -43.7584,
  -43.7481,
  -43.7371,
  -43.7258,
  -43.7147,
  -43.7042,
  -43.6946,
  -43.6857,
  -43.6775,
  -43.6702,
  -43.6629,
  -43.6556,
  -43.6472,
  -43.6373,
  -43.6258,
  -43.6138,
  -43.6015,
  -43.5898,
  -43.5786,
  -43.5673,
  -43.5579,
  -43.5487,
  -43.5392,
  -43.5293,
  -43.5181,
  -43.5056,
  -43.4916,
  -43.4763,
  -43.4592,
  -43.4401,
  -43.42,
  -43.3989,
  -43.3772,
  -43.3545,
  -43.3303,
  -43.3045,
  -43.2766,
  -43.2473,
  -43.2174,
  -43.188,
  -43.1604,
  -43.1354,
  -43.1135,
  -43.0951,
  -43.0799,
  -43.0661,
  -43.0552,
  -43.0451,
  -43.0345,
  -43.0233,
  -43.0109,
  -42.9979,
  -42.9844,
  -42.9707,
  -42.9575,
  -42.9453,
  -42.9345,
  -42.9257,
  -42.9187,
  -42.9138,
  -42.9116,
  -42.9114,
  -42.9122,
  -42.9136,
  -42.9148,
  -42.9134,
  -42.9076,
  -42.8975,
  -42.8821,
  -42.8623,
  -42.8381,
  -42.8109,
  -42.7828,
  -42.755,
  -42.7286,
  -42.7042,
  -42.6803,
  -42.6574,
  -42.6329,
  -42.605,
  -42.5723,
  -42.5343,
  -42.4915,
  -42.4452,
  -42.398,
  -42.3515,
  -42.3083,
  -42.2702,
  -42.2385,
  -42.2138,
  -42.1962,
  -42.1854,
  -42.1809,
  -42.1837,
  -42.1938,
  -42.211,
  -42.2346,
  -42.2644,
  -42.2992,
  -42.3375,
  -42.377,
  -42.4166,
  -42.455,
  -42.4917,
  -42.5265,
  -42.56,
  -42.5935,
  -42.6282,
  -42.6649,
  -42.704,
  -42.7454,
  -42.789,
  -42.8338,
  -42.8779,
  -42.9218,
  -42.9637,
  -43.0017,
  -43.0346,
  -43.062,
  -43.0836,
  -43.0985,
  -43.1049,
  -43.1023,
  -43.089,
  -43.0636,
  -43.0252,
  -42.9731,
  -42.9075,
  -42.8288,
  -42.7379,
  -42.6356,
  -42.5229,
  -42.4018,
  -42.2727,
  -42.1376,
  -41.9975,
  -41.8532,
  -41.7059,
  -41.5571,
  -41.4088,
  -41.263,
  -41.1221,
  -40.9887,
  -40.8643,
  -41.2643,
  -41.3132,
  -41.3618,
  -41.4099,
  -41.4569,
  -41.5028,
  -41.5469,
  -41.5912,
  -41.6345,
  -41.6771,
  -41.7199,
  -41.7631,
  -41.8064,
  -41.8506,
  -41.8952,
  -41.9396,
  -41.9835,
  -42.0266,
  -42.0688,
  -42.1112,
  -42.151,
  -42.1925,
  -42.2327,
  -42.2735,
  -42.314,
  -42.3551,
  -42.3965,
  -42.4384,
  -42.4805,
  -42.5225,
  -42.5642,
  -42.605,
  -42.6441,
  -42.6807,
  -42.7139,
  -42.7436,
  -42.7689,
  -42.7918,
  -42.8112,
  -42.8275,
  -42.8415,
  -42.8531,
  -42.8631,
  -42.8719,
  -42.8805,
  -42.8881,
  -42.8952,
  -42.9018,
  -42.9073,
  -42.9106,
  -42.9118,
  -42.9096,
  -42.9063,
  -42.9009,
  -42.8941,
  -42.8868,
  -42.8789,
  -42.8706,
  -42.8617,
  -42.8528,
  -42.8428,
  -42.8332,
  -42.8236,
  -42.8141,
  -42.8049,
  -42.7965,
  -42.7885,
  -42.7812,
  -42.7734,
  -42.7676,
  -42.7622,
  -42.7577,
  -42.7536,
  -42.7498,
  -42.7466,
  -42.7446,
  -42.7441,
  -42.7461,
  -42.7508,
  -42.7589,
  -42.7701,
  -42.7834,
  -42.7986,
  -42.815,
  -42.8319,
  -42.8483,
  -42.8661,
  -42.8845,
  -42.9028,
  -42.9217,
  -42.9394,
  -42.9567,
  -42.972,
  -42.9856,
  -42.9978,
  -43.009,
  -43.0197,
  -43.0309,
  -43.0425,
  -43.0546,
  -43.0673,
  -43.0802,
  -43.0932,
  -43.1059,
  -43.1171,
  -43.1289,
  -43.1408,
  -43.1532,
  -43.1677,
  -43.1846,
  -43.2055,
  -43.2317,
  -43.2639,
  -43.3011,
  -43.3419,
  -43.3847,
  -43.428,
  -43.4701,
  -43.51,
  -43.5473,
  -43.5818,
  -43.6136,
  -43.6432,
  -43.6696,
  -43.6954,
  -43.7194,
  -43.7416,
  -43.7618,
  -43.7798,
  -43.7955,
  -43.8092,
  -43.821,
  -43.8316,
  -43.8416,
  -43.8512,
  -43.8603,
  -43.8689,
  -43.8767,
  -43.8835,
  -43.8887,
  -43.8915,
  -43.8917,
  -43.8894,
  -43.8848,
  -43.8784,
  -43.8697,
  -43.8615,
  -43.8541,
  -43.8478,
  -43.843,
  -43.839,
  -43.8352,
  -43.8318,
  -43.8283,
  -43.8241,
  -43.819,
  -43.8126,
  -43.8051,
  -43.7965,
  -43.787,
  -43.7777,
  -43.7684,
  -43.7597,
  -43.7517,
  -43.7454,
  -43.7393,
  -43.7341,
  -43.7289,
  -43.7227,
  -43.7161,
  -43.7081,
  -43.6986,
  -43.6886,
  -43.6787,
  -43.6692,
  -43.66,
  -43.6513,
  -43.6428,
  -43.6343,
  -43.6253,
  -43.6148,
  -43.6031,
  -43.5903,
  -43.5762,
  -43.5611,
  -43.5443,
  -43.5255,
  -43.5064,
  -43.4868,
  -43.4668,
  -43.4461,
  -43.4239,
  -43.3993,
  -43.3717,
  -43.3431,
  -43.3138,
  -43.2844,
  -43.2561,
  -43.2298,
  -43.206,
  -43.1851,
  -43.1667,
  -43.1506,
  -43.1361,
  -43.1224,
  -43.109,
  -43.0952,
  -43.0814,
  -43.0674,
  -43.0535,
  -43.0398,
  -43.0273,
  -43.0159,
  -43.006,
  -42.9977,
  -42.9908,
  -42.9856,
  -42.9823,
  -42.9802,
  -42.9791,
  -42.9784,
  -42.9776,
  -42.9731,
  -42.9659,
  -42.9543,
  -42.9375,
  -42.917,
  -42.8927,
  -42.8658,
  -42.8381,
  -42.8112,
  -42.7857,
  -42.7621,
  -42.74,
  -42.7185,
  -42.6956,
  -42.6698,
  -42.64,
  -42.6056,
  -42.5673,
  -42.5269,
  -42.4858,
  -42.446,
  -42.4094,
  -42.3781,
  -42.3525,
  -42.3332,
  -42.3199,
  -42.3121,
  -42.3098,
  -42.3134,
  -42.3229,
  -42.3381,
  -42.359,
  -42.3854,
  -42.4163,
  -42.4498,
  -42.4857,
  -42.5214,
  -42.5568,
  -42.5905,
  -42.6225,
  -42.6531,
  -42.6839,
  -42.715,
  -42.7476,
  -42.7821,
  -42.8187,
  -42.8572,
  -42.8967,
  -42.9366,
  -42.9752,
  -43.0115,
  -43.0443,
  -43.0726,
  -43.0961,
  -43.1142,
  -43.1261,
  -43.13,
  -43.1254,
  -43.1108,
  -43.0842,
  -43.0449,
  -42.992,
  -42.9258,
  -42.8466,
  -42.7544,
  -42.6502,
  -42.5362,
  -42.414,
  -42.285,
  -42.1512,
  -42.0142,
  -41.8743,
  -41.7322,
  -41.5888,
  -41.4455,
  -41.304,
  -41.1655,
  -41.0327,
  -40.9066,
  -41.2627,
  -41.3114,
  -41.3607,
  -41.4097,
  -41.4574,
  -41.5045,
  -41.5505,
  -41.5954,
  -41.6391,
  -41.6821,
  -41.7248,
  -41.7677,
  -41.8109,
  -41.8543,
  -41.8977,
  -41.9398,
  -41.9825,
  -42.0242,
  -42.0655,
  -42.1068,
  -42.1472,
  -42.1876,
  -42.2276,
  -42.2674,
  -42.307,
  -42.3468,
  -42.3867,
  -42.4263,
  -42.4658,
  -42.5049,
  -42.5426,
  -42.5801,
  -42.6161,
  -42.6498,
  -42.6806,
  -42.7081,
  -42.7323,
  -42.7529,
  -42.7698,
  -42.7835,
  -42.7946,
  -42.8035,
  -42.8107,
  -42.8177,
  -42.8251,
  -42.8319,
  -42.8373,
  -42.8431,
  -42.8481,
  -42.8513,
  -42.8522,
  -42.8507,
  -42.8469,
  -42.8411,
  -42.8336,
  -42.8249,
  -42.8159,
  -42.8063,
  -42.7965,
  -42.7868,
  -42.7773,
  -42.7681,
  -42.7586,
  -42.7508,
  -42.7438,
  -42.7382,
  -42.7328,
  -42.7284,
  -42.7249,
  -42.7221,
  -42.7197,
  -42.7176,
  -42.716,
  -42.715,
  -42.7141,
  -42.7138,
  -42.7149,
  -42.7182,
  -42.7242,
  -42.7324,
  -42.7446,
  -42.7592,
  -42.7752,
  -42.7923,
  -42.8101,
  -42.8285,
  -42.8474,
  -42.8666,
  -42.8862,
  -42.9051,
  -42.9235,
  -42.9409,
  -42.9565,
  -42.9706,
  -42.984,
  -42.9967,
  -43.0097,
  -43.0231,
  -43.0359,
  -43.0508,
  -43.0666,
  -43.083,
  -43.0997,
  -43.1165,
  -43.1328,
  -43.1492,
  -43.1653,
  -43.1818,
  -43.1988,
  -43.2176,
  -43.239,
  -43.2641,
  -43.2939,
  -43.3282,
  -43.366,
  -43.4056,
  -43.4454,
  -43.4841,
  -43.5219,
  -43.5578,
  -43.5912,
  -43.6222,
  -43.6509,
  -43.6782,
  -43.7038,
  -43.7277,
  -43.7496,
  -43.7698,
  -43.7879,
  -43.8041,
  -43.8182,
  -43.8307,
  -43.8422,
  -43.853,
  -43.8632,
  -43.8731,
  -43.8824,
  -43.89,
  -43.8973,
  -43.9029,
  -43.9061,
  -43.9067,
  -43.905,
  -43.901,
  -43.8955,
  -43.8887,
  -43.8818,
  -43.8755,
  -43.8707,
  -43.8675,
  -43.8655,
  -43.8641,
  -43.863,
  -43.8615,
  -43.8594,
  -43.856,
  -43.851,
  -43.8449,
  -43.8376,
  -43.8298,
  -43.8208,
  -43.8129,
  -43.8059,
  -43.8,
  -43.7955,
  -43.7914,
  -43.7878,
  -43.7844,
  -43.7809,
  -43.7763,
  -43.77,
  -43.7624,
  -43.7544,
  -43.7467,
  -43.7393,
  -43.7322,
  -43.7253,
  -43.718,
  -43.7098,
  -43.7011,
  -43.6907,
  -43.679,
  -43.6664,
  -43.6524,
  -43.6366,
  -43.6199,
  -43.6024,
  -43.5838,
  -43.5655,
  -43.5469,
  -43.5275,
  -43.5063,
  -43.4828,
  -43.457,
  -43.4295,
  -43.4008,
  -43.3719,
  -43.3436,
  -43.3172,
  -43.293,
  -43.2711,
  -43.2515,
  -43.2334,
  -43.2165,
  -43.2004,
  -43.1845,
  -43.1688,
  -43.1536,
  -43.1387,
  -43.1245,
  -43.1111,
  -43.0991,
  -43.0874,
  -43.078,
  -43.0701,
  -43.0633,
  -43.0574,
  -43.0526,
  -43.0487,
  -43.0456,
  -43.043,
  -43.0395,
  -43.0338,
  -43.0247,
  -43.0117,
  -42.9945,
  -42.9737,
  -42.95,
  -42.9243,
  -42.8981,
  -42.8727,
  -42.8487,
  -42.8261,
  -42.805,
  -42.7842,
  -42.7626,
  -42.7384,
  -42.711,
  -42.6798,
  -42.6455,
  -42.6098,
  -42.574,
  -42.5397,
  -42.5091,
  -42.4823,
  -42.4619,
  -42.4468,
  -42.4368,
  -42.4314,
  -42.4306,
  -42.4346,
  -42.4433,
  -42.4567,
  -42.4749,
  -42.4977,
  -42.5247,
  -42.5548,
  -42.5866,
  -42.6188,
  -42.6505,
  -42.681,
  -42.7102,
  -42.7381,
  -42.7659,
  -42.7938,
  -42.8226,
  -42.853,
  -42.8848,
  -42.9184,
  -42.9531,
  -42.9877,
  -43.0213,
  -43.0525,
  -43.0807,
  -43.1052,
  -43.1252,
  -43.1402,
  -43.1492,
  -43.1509,
  -43.1448,
  -43.1288,
  -43.1011,
  -43.0612,
  -43.0077,
  -42.9396,
  -42.8587,
  -42.7649,
  -42.6585,
  -42.5416,
  -42.417,
  -42.2867,
  -42.1532,
  -42.0185,
  -41.8825,
  -41.7464,
  -41.61,
  -41.4739,
  -41.3391,
  -41.2065,
  -41.0773,
  -40.9526,
  -41.2576,
  -41.3076,
  -41.357,
  -41.4062,
  -41.4545,
  -41.5021,
  -41.5487,
  -41.5939,
  -41.6382,
  -41.6815,
  -41.7236,
  -41.7666,
  -41.8096,
  -41.8524,
  -41.8947,
  -41.9365,
  -41.9778,
  -42.0187,
  -42.0592,
  -42.0995,
  -42.1398,
  -42.1797,
  -42.2192,
  -42.2586,
  -42.2978,
  -42.3358,
  -42.3744,
  -42.4123,
  -42.4493,
  -42.4856,
  -42.5212,
  -42.5557,
  -42.5887,
  -42.6198,
  -42.6482,
  -42.6732,
  -42.6949,
  -42.7129,
  -42.7271,
  -42.7377,
  -42.7457,
  -42.7508,
  -42.7562,
  -42.7615,
  -42.7669,
  -42.7727,
  -42.7787,
  -42.7845,
  -42.7894,
  -42.7925,
  -42.7935,
  -42.7918,
  -42.7879,
  -42.7817,
  -42.7738,
  -42.7642,
  -42.7541,
  -42.7426,
  -42.7324,
  -42.7228,
  -42.7138,
  -42.7057,
  -42.6988,
  -42.693,
  -42.6883,
  -42.6851,
  -42.6827,
  -42.6814,
  -42.6809,
  -42.681,
  -42.6815,
  -42.6822,
  -42.6833,
  -42.6843,
  -42.6847,
  -42.6861,
  -42.6887,
  -42.6932,
  -42.7002,
  -42.7104,
  -42.7233,
  -42.7385,
  -42.7548,
  -42.7722,
  -42.7905,
  -42.8095,
  -42.8288,
  -42.8485,
  -42.8681,
  -42.8873,
  -42.9057,
  -42.9223,
  -42.9385,
  -42.9537,
  -42.9681,
  -42.9824,
  -42.9972,
  -43.0124,
  -43.0287,
  -43.0462,
  -43.0649,
  -43.0844,
  -43.1041,
  -43.1244,
  -43.1445,
  -43.1645,
  -43.1842,
  -43.2038,
  -43.2234,
  -43.2439,
  -43.265,
  -43.2895,
  -43.3176,
  -43.3495,
  -43.3848,
  -43.4218,
  -43.4589,
  -43.4961,
  -43.5322,
  -43.5663,
  -43.598,
  -43.6276,
  -43.6551,
  -43.6813,
  -43.7061,
  -43.7294,
  -43.751,
  -43.771,
  -43.7891,
  -43.8054,
  -43.819,
  -43.8323,
  -43.8444,
  -43.8558,
  -43.8668,
  -43.8775,
  -43.8876,
  -43.897,
  -43.9049,
  -43.9111,
  -43.9149,
  -43.9162,
  -43.9154,
  -43.9126,
  -43.9083,
  -43.9032,
  -43.8979,
  -43.8932,
  -43.8901,
  -43.8886,
  -43.8883,
  -43.8887,
  -43.8883,
  -43.8886,
  -43.8879,
  -43.8857,
  -43.8819,
  -43.8771,
  -43.8711,
  -43.8646,
  -43.8577,
  -43.8515,
  -43.8461,
  -43.8417,
  -43.8383,
  -43.8358,
  -43.8341,
  -43.8325,
  -43.8304,
  -43.8273,
  -43.8227,
  -43.8167,
  -43.8105,
  -43.8045,
  -43.7987,
  -43.7933,
  -43.7868,
  -43.7807,
  -43.7734,
  -43.765,
  -43.755,
  -43.7436,
  -43.7313,
  -43.7179,
  -43.7036,
  -43.6882,
  -43.6711,
  -43.6539,
  -43.6358,
  -43.6182,
  -43.5994,
  -43.5785,
  -43.5564,
  -43.5316,
  -43.505,
  -43.4772,
  -43.4493,
  -43.4221,
  -43.3962,
  -43.3728,
  -43.3514,
  -43.3316,
  -43.312,
  -43.2939,
  -43.276,
  -43.2583,
  -43.2412,
  -43.225,
  -43.2094,
  -43.195,
  -43.1817,
  -43.17,
  -43.1597,
  -43.1505,
  -43.1426,
  -43.1353,
  -43.1287,
  -43.1227,
  -43.1173,
  -43.1124,
  -43.1075,
  -43.1015,
  -43.0937,
  -43.083,
  -43.0688,
  -43.0515,
  -43.0313,
  -43.0087,
  -42.9847,
  -42.9606,
  -42.9369,
  -42.9144,
  -42.8918,
  -42.8717,
  -42.8516,
  -42.8306,
  -42.8079,
  -42.7824,
  -42.754,
  -42.7233,
  -42.6913,
  -42.6599,
  -42.6305,
  -42.6047,
  -42.5833,
  -42.5669,
  -42.555,
  -42.547,
  -42.5434,
  -42.544,
  -42.5484,
  -42.5565,
  -42.5682,
  -42.5836,
  -42.6031,
  -42.6261,
  -42.6519,
  -42.6795,
  -42.708,
  -42.7359,
  -42.7631,
  -42.7887,
  -42.8139,
  -42.8388,
  -42.8638,
  -42.8892,
  -42.9157,
  -42.9432,
  -42.9723,
  -43.0012,
  -43.031,
  -43.0598,
  -43.0862,
  -43.1103,
  -43.1314,
  -43.1484,
  -43.1604,
  -43.1672,
  -43.1671,
  -43.1596,
  -43.1422,
  -43.1137,
  -43.0728,
  -43.0185,
  -42.9503,
  -42.8678,
  -42.7713,
  -42.6623,
  -42.5423,
  -42.4143,
  -42.2818,
  -42.1478,
  -42.0143,
  -41.8823,
  -41.7521,
  -41.6231,
  -41.4953,
  -41.3688,
  -41.244,
  -41.1211,
  -41.0003,
  -41.2508,
  -41.3,
  -41.3492,
  -41.3981,
  -41.4464,
  -41.4943,
  -41.5402,
  -41.586,
  -41.6307,
  -41.6747,
  -41.7183,
  -41.7615,
  -41.8044,
  -41.8468,
  -41.8884,
  -41.9292,
  -41.9695,
  -42.0095,
  -42.0493,
  -42.0893,
  -42.1284,
  -42.1684,
  -42.208,
  -42.2473,
  -42.2861,
  -42.3244,
  -42.3617,
  -42.398,
  -42.433,
  -42.4669,
  -42.4998,
  -42.5315,
  -42.5618,
  -42.59,
  -42.6158,
  -42.6374,
  -42.6565,
  -42.6715,
  -42.6827,
  -42.6902,
  -42.695,
  -42.6985,
  -42.7015,
  -42.7049,
  -42.7091,
  -42.7141,
  -42.7198,
  -42.7257,
  -42.7307,
  -42.7341,
  -42.7355,
  -42.733,
  -42.7289,
  -42.7224,
  -42.7141,
  -42.7042,
  -42.6932,
  -42.6826,
  -42.6724,
  -42.6632,
  -42.6552,
  -42.6487,
  -42.6439,
  -42.6403,
  -42.638,
  -42.6371,
  -42.6376,
  -42.639,
  -42.6403,
  -42.6432,
  -42.6465,
  -42.6499,
  -42.6534,
  -42.6568,
  -42.6601,
  -42.6634,
  -42.6673,
  -42.6729,
  -42.6808,
  -42.6917,
  -42.705,
  -42.7204,
  -42.737,
  -42.7543,
  -42.7723,
  -42.7903,
  -42.8096,
  -42.8291,
  -42.8485,
  -42.8676,
  -42.886,
  -42.9037,
  -42.9208,
  -42.9368,
  -42.9525,
  -42.9683,
  -42.9846,
  -43.0018,
  -43.0201,
  -43.0399,
  -43.0611,
  -43.0832,
  -43.1061,
  -43.1292,
  -43.1514,
  -43.1744,
  -43.197,
  -43.2191,
  -43.2409,
  -43.263,
  -43.2859,
  -43.3105,
  -43.3376,
  -43.3677,
  -43.4006,
  -43.4353,
  -43.4705,
  -43.5054,
  -43.5393,
  -43.5718,
  -43.6017,
  -43.6297,
  -43.6556,
  -43.6792,
  -43.7027,
  -43.7248,
  -43.7454,
  -43.7649,
  -43.7827,
  -43.7992,
  -43.8142,
  -43.8281,
  -43.841,
  -43.8532,
  -43.865,
  -43.8764,
  -43.8873,
  -43.8974,
  -43.9061,
  -43.913,
  -43.9176,
  -43.92,
  -43.9203,
  -43.9191,
  -43.9154,
  -43.9122,
  -43.9086,
  -43.906,
  -43.9045,
  -43.9047,
  -43.906,
  -43.9077,
  -43.9094,
  -43.9108,
  -43.9112,
  -43.91,
  -43.9072,
  -43.9033,
  -43.8984,
  -43.8932,
  -43.8878,
  -43.8828,
  -43.8788,
  -43.8758,
  -43.8738,
  -43.8728,
  -43.8723,
  -43.871,
  -43.8703,
  -43.8685,
  -43.8652,
  -43.8607,
  -43.8558,
  -43.8513,
  -43.847,
  -43.8427,
  -43.8384,
  -43.8335,
  -43.8272,
  -43.8194,
  -43.8099,
  -43.7991,
  -43.7871,
  -43.7744,
  -43.7611,
  -43.7467,
  -43.7312,
  -43.7144,
  -43.6973,
  -43.68,
  -43.6617,
  -43.6417,
  -43.6199,
  -43.595,
  -43.5695,
  -43.543,
  -43.5165,
  -43.4907,
  -43.4665,
  -43.4442,
  -43.424,
  -43.4049,
  -43.3865,
  -43.3681,
  -43.3496,
  -43.3309,
  -43.313,
  -43.2958,
  -43.2798,
  -43.2652,
  -43.2519,
  -43.2402,
  -43.23,
  -43.2207,
  -43.2122,
  -43.2042,
  -43.1969,
  -43.1897,
  -43.1827,
  -43.1761,
  -43.1691,
  -43.1611,
  -43.1501,
  -43.1381,
  -43.1234,
  -43.1066,
  -43.0874,
  -43.0666,
  -43.0446,
  -43.0224,
  -43.0006,
  -42.9794,
  -42.959,
  -42.9392,
  -42.9197,
  -42.8994,
  -42.8779,
  -42.8541,
  -42.8282,
  -42.8005,
  -42.772,
  -42.7443,
  -42.7189,
  -42.697,
  -42.679,
  -42.6651,
  -42.6555,
  -42.6495,
  -42.6471,
  -42.6483,
  -42.6528,
  -42.6602,
  -42.6699,
  -42.6828,
  -42.6992,
  -42.7186,
  -42.7395,
  -42.7635,
  -42.7879,
  -42.8123,
  -42.8356,
  -42.8586,
  -42.8808,
  -42.9026,
  -42.9245,
  -42.9467,
  -42.9696,
  -42.9933,
  -43.0183,
  -43.0439,
  -43.0692,
  -43.0934,
  -43.1159,
  -43.1364,
  -43.154,
  -43.168,
  -43.1777,
  -43.1823,
  -43.1808,
  -43.1717,
  -43.1532,
  -43.1236,
  -43.0818,
  -43.0264,
  -42.9569,
  -42.8728,
  -42.774,
  -42.6617,
  -42.5379,
  -42.4064,
  -42.2713,
  -42.1358,
  -42.0029,
  -41.8738,
  -41.7487,
  -41.6269,
  -41.5076,
  -41.3902,
  -41.2741,
  -41.1589,
  -41.0439,
  -41.2405,
  -41.2874,
  -41.3357,
  -41.384,
  -41.4318,
  -41.4797,
  -41.5269,
  -41.5731,
  -41.6187,
  -41.6635,
  -41.7081,
  -41.7519,
  -41.7949,
  -41.8371,
  -41.8779,
  -41.9168,
  -41.9563,
  -41.9958,
  -42.0356,
  -42.0756,
  -42.1161,
  -42.1563,
  -42.1962,
  -42.2353,
  -42.2738,
  -42.3111,
  -42.3474,
  -42.3823,
  -42.4158,
  -42.4478,
  -42.4774,
  -42.5065,
  -42.534,
  -42.5596,
  -42.5827,
  -42.6026,
  -42.6187,
  -42.6308,
  -42.6388,
  -42.6433,
  -42.6449,
  -42.6457,
  -42.6465,
  -42.6484,
  -42.6516,
  -42.6561,
  -42.6606,
  -42.6665,
  -42.6718,
  -42.6758,
  -42.6771,
  -42.676,
  -42.672,
  -42.6655,
  -42.657,
  -42.6471,
  -42.6363,
  -42.6258,
  -42.6164,
  -42.6082,
  -42.6019,
  -42.5972,
  -42.5935,
  -42.5922,
  -42.5922,
  -42.5932,
  -42.5958,
  -42.5997,
  -42.6045,
  -42.6103,
  -42.6163,
  -42.6223,
  -42.628,
  -42.6335,
  -42.6388,
  -42.6439,
  -42.6494,
  -42.6563,
  -42.6648,
  -42.6752,
  -42.6889,
  -42.7042,
  -42.7204,
  -42.7373,
  -42.7547,
  -42.7728,
  -42.7916,
  -42.8106,
  -42.8297,
  -42.8483,
  -42.8665,
  -42.8845,
  -42.9022,
  -42.9195,
  -42.9365,
  -42.9536,
  -42.9714,
  -42.9894,
  -43.0094,
  -43.031,
  -43.0544,
  -43.0792,
  -43.1045,
  -43.1303,
  -43.1559,
  -43.1814,
  -43.2061,
  -43.2302,
  -43.2539,
  -43.2774,
  -43.3012,
  -43.3262,
  -43.3527,
  -43.3814,
  -43.4124,
  -43.445,
  -43.4782,
  -43.5101,
  -43.542,
  -43.5722,
  -43.6003,
  -43.6264,
  -43.6502,
  -43.673,
  -43.6948,
  -43.7154,
  -43.735,
  -43.7534,
  -43.7709,
  -43.7876,
  -43.803,
  -43.8174,
  -43.831,
  -43.8441,
  -43.8567,
  -43.8689,
  -43.8806,
  -43.8905,
  -43.9,
  -43.9077,
  -43.9133,
  -43.9168,
  -43.9185,
  -43.9188,
  -43.9181,
  -43.9168,
  -43.9155,
  -43.9149,
  -43.9152,
  -43.9169,
  -43.9192,
  -43.922,
  -43.9247,
  -43.9268,
  -43.9278,
  -43.9273,
  -43.9254,
  -43.9226,
  -43.9188,
  -43.9137,
  -43.9095,
  -43.9058,
  -43.9029,
  -43.9013,
  -43.9007,
  -43.901,
  -43.9017,
  -43.9026,
  -43.9028,
  -43.9024,
  -43.9005,
  -43.897,
  -43.8933,
  -43.8897,
  -43.8864,
  -43.8832,
  -43.8798,
  -43.8758,
  -43.8704,
  -43.8635,
  -43.8548,
  -43.8444,
  -43.8331,
  -43.8212,
  -43.808,
  -43.7952,
  -43.7811,
  -43.7658,
  -43.7497,
  -43.7327,
  -43.7147,
  -43.6951,
  -43.6738,
  -43.6507,
  -43.6264,
  -43.6013,
  -43.5763,
  -43.5522,
  -43.5298,
  -43.5093,
  -43.4904,
  -43.4725,
  -43.4547,
  -43.4367,
  -43.418,
  -43.3992,
  -43.3807,
  -43.363,
  -43.3468,
  -43.332,
  -43.3187,
  -43.3057,
  -43.2949,
  -43.285,
  -43.276,
  -43.2672,
  -43.2586,
  -43.2504,
  -43.2425,
  -43.2346,
  -43.2259,
  -43.2159,
  -43.2045,
  -43.1912,
  -43.1765,
  -43.1604,
  -43.1427,
  -43.1236,
  -43.1039,
  -43.0838,
  -43.0637,
  -43.0437,
  -43.024,
  -43.0049,
  -42.9857,
  -42.9662,
  -42.9457,
  -42.9235,
  -42.8996,
  -42.8746,
  -42.8492,
  -42.8247,
  -42.8029,
  -42.784,
  -42.7679,
  -42.7563,
  -42.748,
  -42.7431,
  -42.7417,
  -42.7432,
  -42.7473,
  -42.7535,
  -42.7618,
  -42.7722,
  -42.7855,
  -42.8013,
  -42.8197,
  -42.8399,
  -42.8608,
  -42.8816,
  -42.9016,
  -42.9212,
  -42.9404,
  -42.9594,
  -42.9786,
  -42.9979,
  -43.0177,
  -43.038,
  -43.0592,
  -43.0807,
  -43.1022,
  -43.1226,
  -43.1417,
  -43.1589,
  -43.1735,
  -43.1847,
  -43.1919,
  -43.1944,
  -43.1909,
  -43.1802,
  -43.1604,
  -43.1295,
  -43.0867,
  -43.0305,
  -42.9586,
  -42.8727,
  -42.7719,
  -42.6567,
  -42.5296,
  -42.3945,
  -42.2561,
  -42.1185,
  -41.9851,
  -41.8577,
  -41.7366,
  -41.6208,
  -41.5092,
  -41.4004,
  -41.293,
  -41.186,
  -41.078,
  -41.2246,
  -41.2711,
  -41.3182,
  -41.3656,
  -41.4132,
  -41.4608,
  -41.5083,
  -41.5553,
  -41.6016,
  -41.6474,
  -41.6916,
  -41.7363,
  -41.7796,
  -41.8216,
  -41.8621,
  -41.9017,
  -41.9407,
  -41.9799,
  -42.0198,
  -42.0602,
  -42.101,
  -42.1414,
  -42.1814,
  -42.2207,
  -42.259,
  -42.295,
  -42.3305,
  -42.3642,
  -42.3962,
  -42.4266,
  -42.4551,
  -42.4819,
  -42.507,
  -42.5301,
  -42.5505,
  -42.5679,
  -42.5812,
  -42.5902,
  -42.5954,
  -42.5969,
  -42.5958,
  -42.593,
  -42.5918,
  -42.5921,
  -42.5945,
  -42.5986,
  -42.604,
  -42.6098,
  -42.6155,
  -42.6194,
  -42.6212,
  -42.6204,
  -42.6168,
  -42.6104,
  -42.6022,
  -42.5926,
  -42.5825,
  -42.5715,
  -42.5632,
  -42.5568,
  -42.5526,
  -42.5501,
  -42.5492,
  -42.5501,
  -42.552,
  -42.555,
  -42.5594,
  -42.5651,
  -42.5722,
  -42.5803,
  -42.5888,
  -42.5971,
  -42.605,
  -42.6112,
  -42.6184,
  -42.6252,
  -42.6323,
  -42.6401,
  -42.6497,
  -42.6617,
  -42.6756,
  -42.6907,
  -42.7065,
  -42.7228,
  -42.7392,
  -42.7562,
  -42.7738,
  -42.792,
  -42.8106,
  -42.8289,
  -42.847,
  -42.8642,
  -42.8824,
  -42.9008,
  -42.919,
  -42.9373,
  -42.9566,
  -42.9768,
  -42.9987,
  -43.0218,
  -43.047,
  -43.0735,
  -43.1011,
  -43.129,
  -43.1567,
  -43.1841,
  -43.2105,
  -43.2362,
  -43.2614,
  -43.2861,
  -43.3098,
  -43.335,
  -43.3614,
  -43.3891,
  -43.4184,
  -43.4488,
  -43.4801,
  -43.5112,
  -43.541,
  -43.5691,
  -43.5952,
  -43.6191,
  -43.6414,
  -43.6622,
  -43.682,
  -43.7009,
  -43.7191,
  -43.7365,
  -43.7535,
  -43.77,
  -43.7847,
  -43.7997,
  -43.8141,
  -43.8279,
  -43.8413,
  -43.8543,
  -43.8666,
  -43.8782,
  -43.8883,
  -43.8968,
  -43.9034,
  -43.9081,
  -43.9114,
  -43.9135,
  -43.9149,
  -43.9156,
  -43.9165,
  -43.9178,
  -43.9199,
  -43.9227,
  -43.926,
  -43.9295,
  -43.9318,
  -43.9344,
  -43.9361,
  -43.9363,
  -43.9352,
  -43.9333,
  -43.9309,
  -43.9279,
  -43.9248,
  -43.9221,
  -43.9208,
  -43.9204,
  -43.9211,
  -43.9225,
  -43.924,
  -43.9257,
  -43.9269,
  -43.9275,
  -43.9266,
  -43.924,
  -43.9213,
  -43.9184,
  -43.9159,
  -43.9128,
  -43.9102,
  -43.907,
  -43.9025,
  -43.8967,
  -43.8888,
  -43.8791,
  -43.8686,
  -43.8577,
  -43.8466,
  -43.8351,
  -43.8225,
  -43.8085,
  -43.7935,
  -43.7773,
  -43.7596,
  -43.7407,
  -43.7199,
  -43.6979,
  -43.6749,
  -43.6513,
  -43.628,
  -43.6057,
  -43.5851,
  -43.5662,
  -43.5487,
  -43.5316,
  -43.5139,
  -43.4963,
  -43.4782,
  -43.4596,
  -43.4411,
  -43.4234,
  -43.4072,
  -43.3926,
  -43.3794,
  -43.3673,
  -43.3559,
  -43.3452,
  -43.3351,
  -43.3253,
  -43.3155,
  -43.3061,
  -43.2971,
  -43.2878,
  -43.2778,
  -43.2664,
  -43.2541,
  -43.2403,
  -43.2258,
  -43.2106,
  -43.1942,
  -43.177,
  -43.159,
  -43.1405,
  -43.1218,
  -43.1028,
  -43.0829,
  -43.0643,
  -43.0459,
  -43.0276,
  -43.0084,
  -42.9882,
  -42.9665,
  -42.9438,
  -42.9212,
  -42.8998,
  -42.8807,
  -42.8645,
  -42.8512,
  -42.8411,
  -42.834,
  -42.8301,
  -42.8289,
  -42.8303,
  -42.8339,
  -42.8389,
  -42.8456,
  -42.854,
  -42.8644,
  -42.8772,
  -42.8922,
  -42.9087,
  -42.9263,
  -42.9437,
  -42.9607,
  -42.9773,
  -42.9935,
  -43.0097,
  -43.0261,
  -43.0424,
  -43.0592,
  -43.0767,
  -43.0943,
  -43.1111,
  -43.1291,
  -43.1463,
  -43.1624,
  -43.1768,
  -43.1883,
  -43.1969,
  -43.2015,
  -43.2017,
  -43.196,
  -43.1834,
  -43.162,
  -43.13,
  -43.0861,
  -43.0291,
  -42.9575,
  -42.8703,
  -42.7678,
  -42.6503,
  -42.5205,
  -42.3822,
  -42.2404,
  -42.1001,
  -41.9651,
  -41.8379,
  -41.7191,
  -41.6077,
  -41.5022,
  -41.4007,
  -41.3013,
  -41.2022,
  -41.1015,
  -41.2035,
  -41.2489,
  -41.2951,
  -41.3418,
  -41.3892,
  -41.4359,
  -41.4836,
  -41.5313,
  -41.5784,
  -41.625,
  -41.6711,
  -41.7163,
  -41.7601,
  -41.8023,
  -41.8428,
  -41.8823,
  -41.9212,
  -41.9607,
  -42.0007,
  -42.0413,
  -42.0813,
  -42.1221,
  -42.1623,
  -42.2019,
  -42.2402,
  -42.2768,
  -42.3115,
  -42.3442,
  -42.3751,
  -42.4038,
  -42.4307,
  -42.4555,
  -42.4782,
  -42.499,
  -42.517,
  -42.5308,
  -42.5416,
  -42.5481,
  -42.5506,
  -42.5498,
  -42.5466,
  -42.5429,
  -42.5399,
  -42.5392,
  -42.5405,
  -42.5443,
  -42.5493,
  -42.555,
  -42.5605,
  -42.5647,
  -42.5668,
  -42.5655,
  -42.5624,
  -42.5565,
  -42.5487,
  -42.5398,
  -42.5308,
  -42.5224,
  -42.5154,
  -42.5108,
  -42.5082,
  -42.5079,
  -42.5089,
  -42.5116,
  -42.5154,
  -42.5202,
  -42.5264,
  -42.534,
  -42.5421,
  -42.5519,
  -42.5619,
  -42.5722,
  -42.5818,
  -42.5908,
  -42.5993,
  -42.6077,
  -42.6161,
  -42.6254,
  -42.636,
  -42.6481,
  -42.6621,
  -42.6772,
  -42.6929,
  -42.7084,
  -42.7239,
  -42.7383,
  -42.7549,
  -42.7723,
  -42.7898,
  -42.8079,
  -42.8259,
  -42.8444,
  -42.8629,
  -42.8821,
  -42.9017,
  -42.9212,
  -42.9413,
  -42.9629,
  -42.986,
  -43.0108,
  -43.0371,
  -43.0653,
  -43.0945,
  -43.1241,
  -43.1524,
  -43.1812,
  -43.209,
  -43.236,
  -43.2623,
  -43.288,
  -43.3133,
  -43.3385,
  -43.3644,
  -43.3912,
  -43.4188,
  -43.4473,
  -43.4765,
  -43.5056,
  -43.5336,
  -43.5597,
  -43.584,
  -43.6063,
  -43.6269,
  -43.645,
  -43.6631,
  -43.6801,
  -43.6967,
  -43.7131,
  -43.7293,
  -43.7455,
  -43.7613,
  -43.7766,
  -43.7914,
  -43.8061,
  -43.82,
  -43.8335,
  -43.8466,
  -43.8586,
  -43.8693,
  -43.8783,
  -43.8858,
  -43.892,
  -43.897,
  -43.901,
  -43.9034,
  -43.9064,
  -43.9093,
  -43.9125,
  -43.916,
  -43.9198,
  -43.9239,
  -43.9279,
  -43.9319,
  -43.9351,
  -43.9372,
  -43.9384,
  -43.9383,
  -43.9375,
  -43.9359,
  -43.9342,
  -43.9326,
  -43.9312,
  -43.9309,
  -43.9314,
  -43.933,
  -43.9355,
  -43.938,
  -43.9392,
  -43.9412,
  -43.9422,
  -43.9419,
  -43.9404,
  -43.9386,
  -43.9365,
  -43.935,
  -43.9337,
  -43.932,
  -43.9297,
  -43.926,
  -43.9207,
  -43.9135,
  -43.9052,
  -43.8958,
  -43.8858,
  -43.876,
  -43.8656,
  -43.8544,
  -43.8418,
  -43.8278,
  -43.8124,
  -43.7955,
  -43.7771,
  -43.7568,
  -43.7357,
  -43.714,
  -43.6919,
  -43.6702,
  -43.6495,
  -43.6304,
  -43.6128,
  -43.5963,
  -43.5803,
  -43.5642,
  -43.5474,
  -43.5299,
  -43.5118,
  -43.4939,
  -43.4767,
  -43.461,
  -43.4467,
  -43.4337,
  -43.4215,
  -43.41,
  -43.3986,
  -43.3875,
  -43.3764,
  -43.3656,
  -43.355,
  -43.3446,
  -43.3342,
  -43.3231,
  -43.31,
  -43.2969,
  -43.283,
  -43.2688,
  -43.2544,
  -43.2392,
  -43.2234,
  -43.2067,
  -43.1895,
  -43.1715,
  -43.1535,
  -43.1352,
  -43.1179,
  -43.1007,
  -43.0838,
  -43.0665,
  -43.0484,
  -43.0289,
  -43.0086,
  -42.9886,
  -42.9702,
  -42.9533,
  -42.9393,
  -42.9275,
  -42.9186,
  -42.9126,
  -42.9093,
  -42.9083,
  -42.9095,
  -42.9121,
  -42.9161,
  -42.9212,
  -42.9276,
  -42.9357,
  -42.9454,
  -42.9562,
  -42.9696,
  -42.9838,
  -42.9982,
  -43.0123,
  -43.0259,
  -43.0393,
  -43.0528,
  -43.0663,
  -43.08,
  -43.094,
  -43.1083,
  -43.1228,
  -43.1374,
  -43.1522,
  -43.1668,
  -43.1804,
  -43.192,
  -43.2011,
  -43.207,
  -43.2089,
  -43.2062,
  -43.1979,
  -43.183,
  -43.16,
  -43.127,
  -43.0824,
  -43.0249,
  -42.9528,
  -42.8653,
  -42.7619,
  -42.643,
  -42.5111,
  -42.37,
  -42.225,
  -42.0815,
  -41.944,
  -41.8155,
  -41.6972,
  -41.5882,
  -41.4866,
  -41.3905,
  -41.2977,
  -41.2058,
  -41.1114,
  -41.1768,
  -41.2202,
  -41.2659,
  -41.3124,
  -41.3594,
  -41.4071,
  -41.4551,
  -41.503,
  -41.5507,
  -41.598,
  -41.6448,
  -41.6904,
  -41.7347,
  -41.7772,
  -41.8181,
  -41.8569,
  -41.8963,
  -41.9358,
  -41.9761,
  -42.017,
  -42.0579,
  -42.099,
  -42.1395,
  -42.1793,
  -42.2176,
  -42.254,
  -42.2881,
  -42.32,
  -42.3497,
  -42.3771,
  -42.4014,
  -42.4244,
  -42.4452,
  -42.4638,
  -42.4796,
  -42.4923,
  -42.5008,
  -42.5051,
  -42.5057,
  -42.5033,
  -42.4989,
  -42.4939,
  -42.4897,
  -42.4878,
  -42.4886,
  -42.4917,
  -42.4956,
  -42.501,
  -42.5064,
  -42.5107,
  -42.513,
  -42.5132,
  -42.5104,
  -42.5052,
  -42.4986,
  -42.4909,
  -42.4832,
  -42.4767,
  -42.4715,
  -42.4687,
  -42.4681,
  -42.4693,
  -42.4711,
  -42.4752,
  -42.4805,
  -42.487,
  -42.4947,
  -42.5038,
  -42.5143,
  -42.5255,
  -42.537,
  -42.5483,
  -42.5589,
  -42.5691,
  -42.579,
  -42.5888,
  -42.5987,
  -42.6091,
  -42.6207,
  -42.6324,
  -42.6463,
  -42.6612,
  -42.6767,
  -42.6916,
  -42.7061,
  -42.7208,
  -42.7361,
  -42.7522,
  -42.7691,
  -42.7867,
  -42.8043,
  -42.8227,
  -42.8424,
  -42.8621,
  -42.8823,
  -42.9034,
  -42.9247,
  -42.9461,
  -42.97,
  -42.9958,
  -43.0233,
  -43.0525,
  -43.0829,
  -43.1138,
  -43.1444,
  -43.1745,
  -43.2035,
  -43.2314,
  -43.2583,
  -43.2844,
  -43.3098,
  -43.3349,
  -43.3601,
  -43.3858,
  -43.4119,
  -43.4385,
  -43.4643,
  -43.4915,
  -43.5176,
  -43.5421,
  -43.5646,
  -43.5855,
  -43.6047,
  -43.6222,
  -43.6387,
  -43.6542,
  -43.6694,
  -43.6846,
  -43.7001,
  -43.7159,
  -43.7315,
  -43.7471,
  -43.7623,
  -43.7771,
  -43.7915,
  -43.8056,
  -43.8188,
  -43.83,
  -43.841,
  -43.8507,
  -43.8591,
  -43.8666,
  -43.8731,
  -43.8792,
  -43.8846,
  -43.8898,
  -43.8948,
  -43.8997,
  -43.9046,
  -43.9093,
  -43.9139,
  -43.9186,
  -43.9232,
  -43.9272,
  -43.9302,
  -43.9327,
  -43.9338,
  -43.9342,
  -43.9339,
  -43.9325,
  -43.9318,
  -43.9316,
  -43.9324,
  -43.9339,
  -43.9366,
  -43.939,
  -43.9422,
  -43.9451,
  -43.9474,
  -43.9487,
  -43.949,
  -43.9483,
  -43.9471,
  -43.9462,
  -43.9457,
  -43.9452,
  -43.9444,
  -43.9426,
  -43.9395,
  -43.9347,
  -43.9285,
  -43.9208,
  -43.9126,
  -43.9036,
  -43.8938,
  -43.8845,
  -43.8745,
  -43.8632,
  -43.8503,
  -43.8359,
  -43.8204,
  -43.8031,
  -43.7848,
  -43.7651,
  -43.7442,
  -43.7238,
  -43.7038,
  -43.6848,
  -43.667,
  -43.6503,
  -43.6345,
  -43.6191,
  -43.6035,
  -43.5875,
  -43.5706,
  -43.5533,
  -43.5362,
  -43.5199,
  -43.5049,
  -43.4913,
  -43.4787,
  -43.4661,
  -43.4545,
  -43.4427,
  -43.4307,
  -43.4186,
  -43.4065,
  -43.3947,
  -43.3832,
  -43.3719,
  -43.3599,
  -43.3471,
  -43.3337,
  -43.3202,
  -43.3064,
  -43.2924,
  -43.278,
  -43.2628,
  -43.247,
  -43.2305,
  -43.2131,
  -43.1958,
  -43.1791,
  -43.1627,
  -43.1472,
  -43.1323,
  -43.1173,
  -43.1015,
  -43.0847,
  -43.0669,
  -43.0495,
  -43.0333,
  -43.0187,
  -43.0052,
  -42.9948,
  -42.987,
  -42.9819,
  -42.9792,
  -42.9782,
  -42.979,
  -42.9808,
  -42.9838,
  -42.9877,
  -42.9921,
  -42.9979,
  -43.0052,
  -43.014,
  -43.0244,
  -43.0355,
  -43.0471,
  -43.0586,
  -43.0695,
  -43.0802,
  -43.091,
  -43.1018,
  -43.113,
  -43.1245,
  -43.1357,
  -43.1471,
  -43.1589,
  -43.1711,
  -43.1831,
  -43.1942,
  -43.2037,
  -43.2106,
  -43.214,
  -43.213,
  -43.2073,
  -43.1964,
  -43.179,
  -43.1538,
  -43.1196,
  -43.0744,
  -43.0158,
  -42.944,
  -42.8567,
  -42.7533,
  -42.6342,
  -42.5014,
  -42.3584,
  -42.2105,
  -42.0637,
  -41.9228,
  -41.7918,
  -41.6721,
  -41.5633,
  -41.4635,
  -41.3708,
  -41.2825,
  -41.1962,
  -41.1094,
  -41.1425,
  -41.1867,
  -41.2322,
  -41.2789,
  -41.3262,
  -41.3737,
  -41.4217,
  -41.4696,
  -41.5175,
  -41.5651,
  -41.6112,
  -41.6572,
  -41.702,
  -41.7452,
  -41.7868,
  -41.8271,
  -41.8668,
  -41.9068,
  -41.947,
  -41.9879,
  -42.0289,
  -42.07,
  -42.1106,
  -42.1503,
  -42.1885,
  -42.2236,
  -42.2572,
  -42.2884,
  -42.3172,
  -42.3435,
  -42.3676,
  -42.3892,
  -42.4082,
  -42.4249,
  -42.439,
  -42.4496,
  -42.4563,
  -42.4592,
  -42.4588,
  -42.4555,
  -42.4494,
  -42.4438,
  -42.4392,
  -42.4367,
  -42.4368,
  -42.4397,
  -42.4441,
  -42.4496,
  -42.455,
  -42.4592,
  -42.4619,
  -42.4621,
  -42.46,
  -42.4559,
  -42.4499,
  -42.444,
  -42.437,
  -42.4325,
  -42.4295,
  -42.4283,
  -42.4292,
  -42.432,
  -42.436,
  -42.4413,
  -42.4478,
  -42.4559,
  -42.4652,
  -42.4755,
  -42.4869,
  -42.4989,
  -42.5111,
  -42.5229,
  -42.5342,
  -42.5443,
  -42.555,
  -42.5661,
  -42.5772,
  -42.5889,
  -42.6012,
  -42.6145,
  -42.6287,
  -42.6434,
  -42.6586,
  -42.6732,
  -42.6873,
  -42.7012,
  -42.7156,
  -42.7307,
  -42.7469,
  -42.7639,
  -42.7814,
  -42.7989,
  -42.8183,
  -42.8386,
  -42.8597,
  -42.8818,
  -42.9044,
  -42.9276,
  -42.9522,
  -42.9783,
  -43.0064,
  -43.0362,
  -43.0674,
  -43.0991,
  -43.1309,
  -43.162,
  -43.1918,
  -43.2202,
  -43.2473,
  -43.2732,
  -43.2973,
  -43.3218,
  -43.3459,
  -43.3701,
  -43.3947,
  -43.4195,
  -43.4443,
  -43.4692,
  -43.4937,
  -43.5168,
  -43.5382,
  -43.5575,
  -43.5755,
  -43.592,
  -43.6071,
  -43.6214,
  -43.6355,
  -43.6496,
  -43.6644,
  -43.6797,
  -43.694,
  -43.7095,
  -43.7247,
  -43.7394,
  -43.754,
  -43.768,
  -43.7813,
  -43.7935,
  -43.8048,
  -43.8149,
  -43.8241,
  -43.8329,
  -43.8411,
  -43.8489,
  -43.8564,
  -43.8636,
  -43.8705,
  -43.8772,
  -43.8834,
  -43.8891,
  -43.8947,
  -43.899,
  -43.9042,
  -43.9092,
  -43.9137,
  -43.9173,
  -43.9199,
  -43.9217,
  -43.9226,
  -43.9231,
  -43.9237,
  -43.9246,
  -43.9264,
  -43.9289,
  -43.9319,
  -43.9351,
  -43.9383,
  -43.9412,
  -43.9436,
  -43.9453,
  -43.9461,
  -43.9459,
  -43.9457,
  -43.9459,
  -43.9466,
  -43.946,
  -43.9459,
  -43.9446,
  -43.9419,
  -43.9376,
  -43.9318,
  -43.9252,
  -43.9177,
  -43.9099,
  -43.9021,
  -43.8937,
  -43.8847,
  -43.8746,
  -43.863,
  -43.8497,
  -43.8352,
  -43.8193,
  -43.8021,
  -43.7836,
  -43.7647,
  -43.7454,
  -43.7269,
  -43.7092,
  -43.6927,
  -43.6766,
  -43.6611,
  -43.645,
  -43.6299,
  -43.6145,
  -43.5984,
  -43.5819,
  -43.5658,
  -43.5507,
  -43.5368,
  -43.524,
  -43.5122,
  -43.5008,
  -43.4895,
  -43.478,
  -43.4652,
  -43.4524,
  -43.4392,
  -43.4264,
  -43.4142,
  -43.4017,
  -43.3891,
  -43.3759,
  -43.3625,
  -43.3491,
  -43.3355,
  -43.3217,
  -43.3073,
  -43.2924,
  -43.277,
  -43.2609,
  -43.2444,
  -43.2285,
  -43.2117,
  -43.1972,
  -43.1838,
  -43.171,
  -43.1585,
  -43.1452,
  -43.131,
  -43.1162,
  -43.1016,
  -43.0878,
  -43.0749,
  -43.0637,
  -43.0544,
  -43.0475,
  -43.0431,
  -43.0407,
  -43.0399,
  -43.0401,
  -43.0412,
  -43.0434,
  -43.046,
  -43.0489,
  -43.0527,
  -43.0576,
  -43.0641,
  -43.0717,
  -43.0803,
  -43.0895,
  -43.0984,
  -43.1071,
  -43.1153,
  -43.1236,
  -43.1323,
  -43.1409,
  -43.1495,
  -43.158,
  -43.1668,
  -43.1751,
  -43.1848,
  -43.1944,
  -43.2035,
  -43.2109,
  -43.2155,
  -43.2162,
  -43.2125,
  -43.204,
  -43.1903,
  -43.1705,
  -43.1434,
  -43.1078,
  -43.0621,
  -43.0047,
  -42.9334,
  -42.847,
  -42.7446,
  -42.6262,
  -42.4935,
  -42.3497,
  -42.1998,
  -42.0493,
  -41.9049,
  -41.7703,
  -41.6478,
  -41.5371,
  -41.4372,
  -41.3459,
  -41.2606,
  -41.1785,
  -41.0966,
  -41.1029,
  -41.1475,
  -41.1932,
  -41.2401,
  -41.2877,
  -41.3341,
  -41.3817,
  -41.4293,
  -41.477,
  -41.5245,
  -41.5716,
  -41.6179,
  -41.6633,
  -41.7073,
  -41.7496,
  -41.7907,
  -41.831,
  -41.871,
  -41.9111,
  -41.9518,
  -41.9919,
  -42.0328,
  -42.0733,
  -42.1128,
  -42.1507,
  -42.1864,
  -42.2195,
  -42.2502,
  -42.2782,
  -42.3038,
  -42.3271,
  -42.3475,
  -42.3653,
  -42.3804,
  -42.3927,
  -42.4007,
  -42.4063,
  -42.4083,
  -42.4074,
  -42.4039,
  -42.3989,
  -42.3937,
  -42.3894,
  -42.3869,
  -42.3867,
  -42.389,
  -42.3932,
  -42.3987,
  -42.404,
  -42.4084,
  -42.4109,
  -42.4105,
  -42.4089,
  -42.4056,
  -42.4012,
  -42.3967,
  -42.3931,
  -42.3908,
  -42.39,
  -42.3907,
  -42.3928,
  -42.3967,
  -42.4015,
  -42.408,
  -42.4154,
  -42.4248,
  -42.4355,
  -42.447,
  -42.458,
  -42.4703,
  -42.4823,
  -42.494,
  -42.5054,
  -42.5167,
  -42.5281,
  -42.5402,
  -42.5525,
  -42.5653,
  -42.5784,
  -42.5924,
  -42.6071,
  -42.6221,
  -42.6369,
  -42.6515,
  -42.6653,
  -42.6781,
  -42.6917,
  -42.706,
  -42.7214,
  -42.7378,
  -42.755,
  -42.7732,
  -42.7926,
  -42.8135,
  -42.835,
  -42.8579,
  -42.8814,
  -42.9055,
  -42.9303,
  -42.9565,
  -42.9844,
  -43.0143,
  -43.0456,
  -43.0769,
  -43.1093,
  -43.1409,
  -43.1714,
  -43.2001,
  -43.2269,
  -43.2523,
  -43.2763,
  -43.2997,
  -43.3225,
  -43.3451,
  -43.3679,
  -43.391,
  -43.4141,
  -43.4373,
  -43.4601,
  -43.4822,
  -43.5024,
  -43.5209,
  -43.5376,
  -43.5522,
  -43.5665,
  -43.5801,
  -43.5932,
  -43.6066,
  -43.6206,
  -43.6351,
  -43.65,
  -43.6652,
  -43.6799,
  -43.6946,
  -43.7087,
  -43.7224,
  -43.7354,
  -43.7476,
  -43.759,
  -43.7697,
  -43.7797,
  -43.7894,
  -43.7991,
  -43.8088,
  -43.8172,
  -43.8263,
  -43.835,
  -43.8431,
  -43.8507,
  -43.8577,
  -43.8642,
  -43.8706,
  -43.8768,
  -43.8829,
  -43.8885,
  -43.8934,
  -43.8975,
  -43.9005,
  -43.9028,
  -43.9046,
  -43.9064,
  -43.9086,
  -43.9112,
  -43.9143,
  -43.9178,
  -43.9214,
  -43.9246,
  -43.9265,
  -43.9286,
  -43.9305,
  -43.9318,
  -43.9327,
  -43.9336,
  -43.9351,
  -43.9367,
  -43.9382,
  -43.9387,
  -43.9378,
  -43.9353,
  -43.9314,
  -43.9263,
  -43.9203,
  -43.9138,
  -43.9071,
  -43.9002,
  -43.8928,
  -43.8847,
  -43.8752,
  -43.8644,
  -43.8522,
  -43.8389,
  -43.8242,
  -43.8072,
  -43.7903,
  -43.7726,
  -43.7548,
  -43.7375,
  -43.7209,
  -43.7051,
  -43.6898,
  -43.6746,
  -43.6598,
  -43.6449,
  -43.6299,
  -43.6145,
  -43.5993,
  -43.5845,
  -43.5705,
  -43.5577,
  -43.546,
  -43.5348,
  -43.524,
  -43.5132,
  -43.5016,
  -43.489,
  -43.4757,
  -43.462,
  -43.4485,
  -43.4353,
  -43.4221,
  -43.4089,
  -43.3945,
  -43.3812,
  -43.3678,
  -43.3541,
  -43.34,
  -43.3254,
  -43.3105,
  -43.2952,
  -43.2797,
  -43.2642,
  -43.2495,
  -43.2356,
  -43.2233,
  -43.2121,
  -43.2019,
  -43.1917,
  -43.1809,
  -43.1696,
  -43.1578,
  -43.1458,
  -43.1339,
  -43.1227,
  -43.1128,
  -43.1045,
  -43.0983,
  -43.0942,
  -43.0921,
  -43.0909,
  -43.0909,
  -43.0914,
  -43.0928,
  -43.0941,
  -43.0959,
  -43.098,
  -43.1002,
  -43.1045,
  -43.11,
  -43.1166,
  -43.1237,
  -43.1308,
  -43.1373,
  -43.1437,
  -43.15,
  -43.1563,
  -43.1623,
  -43.1682,
  -43.1743,
  -43.1807,
  -43.1876,
  -43.195,
  -43.2026,
  -43.2098,
  -43.2152,
  -43.2175,
  -43.2157,
  -43.2094,
  -43.1981,
  -43.1818,
  -43.16,
  -43.1315,
  -43.0947,
  -43.0483,
  -42.9912,
  -42.9207,
  -42.8354,
  -42.7345,
  -42.6175,
  -42.4857,
  -42.3417,
  -42.1903,
  -42.0377,
  -41.8894,
  -41.7507,
  -41.6242,
  -41.5105,
  -41.4088,
  -41.3173,
  -41.2331,
  -41.1534,
  -41.0742,
  -41.0563,
  -41.1004,
  -41.1467,
  -41.194,
  -41.2416,
  -41.2889,
  -41.3363,
  -41.3835,
  -41.4308,
  -41.478,
  -41.525,
  -41.5716,
  -41.6174,
  -41.662,
  -41.7052,
  -41.7458,
  -41.7864,
  -41.8264,
  -41.8666,
  -41.9071,
  -41.9481,
  -41.9889,
  -42.029,
  -42.0681,
  -42.1054,
  -42.1405,
  -42.173,
  -42.2032,
  -42.2309,
  -42.2561,
  -42.2775,
  -42.2973,
  -42.3141,
  -42.328,
  -42.339,
  -42.3469,
  -42.3516,
  -42.3536,
  -42.3526,
  -42.3495,
  -42.3453,
  -42.341,
  -42.3374,
  -42.3354,
  -42.3354,
  -42.3375,
  -42.3405,
  -42.3457,
  -42.3511,
  -42.3556,
  -42.3581,
  -42.359,
  -42.3582,
  -42.356,
  -42.3532,
  -42.3508,
  -42.3494,
  -42.3494,
  -42.3509,
  -42.3534,
  -42.3569,
  -42.3614,
  -42.3661,
  -42.3732,
  -42.3819,
  -42.3921,
  -42.4037,
  -42.4159,
  -42.4282,
  -42.4402,
  -42.4519,
  -42.4632,
  -42.4741,
  -42.4853,
  -42.4973,
  -42.5099,
  -42.5231,
  -42.5368,
  -42.551,
  -42.5647,
  -42.5797,
  -42.595,
  -42.6099,
  -42.6243,
  -42.6382,
  -42.6517,
  -42.6651,
  -42.6791,
  -42.6936,
  -42.7094,
  -42.7263,
  -42.7443,
  -42.7637,
  -42.7846,
  -42.8068,
  -42.8299,
  -42.8541,
  -42.8775,
  -42.9023,
  -42.9281,
  -42.9555,
  -42.9848,
  -43.0158,
  -43.0478,
  -43.0803,
  -43.1121,
  -43.1427,
  -43.1714,
  -43.198,
  -43.2224,
  -43.2454,
  -43.2672,
  -43.2885,
  -43.3094,
  -43.3303,
  -43.3516,
  -43.3724,
  -43.3942,
  -43.4156,
  -43.4364,
  -43.4559,
  -43.4738,
  -43.4899,
  -43.5045,
  -43.5184,
  -43.5313,
  -43.5441,
  -43.5567,
  -43.5699,
  -43.5838,
  -43.5981,
  -43.6125,
  -43.6267,
  -43.6406,
  -43.6544,
  -43.6673,
  -43.6801,
  -43.6913,
  -43.7029,
  -43.7141,
  -43.725,
  -43.7359,
  -43.7469,
  -43.7581,
  -43.7691,
  -43.7797,
  -43.7898,
  -43.7993,
  -43.8083,
  -43.8166,
  -43.8244,
  -43.8319,
  -43.8393,
  -43.8465,
  -43.8532,
  -43.8596,
  -43.8648,
  -43.8693,
  -43.8729,
  -43.8751,
  -43.8784,
  -43.8817,
  -43.8853,
  -43.8888,
  -43.893,
  -43.8969,
  -43.9001,
  -43.9028,
  -43.9053,
  -43.9077,
  -43.9093,
  -43.9114,
  -43.9134,
  -43.9158,
  -43.9185,
  -43.9207,
  -43.922,
  -43.9216,
  -43.9196,
  -43.9161,
  -43.9115,
  -43.906,
  -43.9004,
  -43.8936,
  -43.8877,
  -43.8808,
  -43.8733,
  -43.8647,
  -43.8546,
  -43.8435,
  -43.831,
  -43.8173,
  -43.8026,
  -43.7868,
  -43.7703,
  -43.7535,
  -43.7374,
  -43.722,
  -43.707,
  -43.692,
  -43.6772,
  -43.6626,
  -43.6483,
  -43.6337,
  -43.6193,
  -43.6052,
  -43.5917,
  -43.579,
  -43.5674,
  -43.5563,
  -43.5457,
  -43.5345,
  -43.5241,
  -43.5127,
  -43.5002,
  -43.4869,
  -43.4731,
  -43.4593,
  -43.4453,
  -43.4316,
  -43.418,
  -43.4047,
  -43.3913,
  -43.3776,
  -43.3637,
  -43.3491,
  -43.3343,
  -43.3192,
  -43.3043,
  -43.2897,
  -43.2756,
  -43.2626,
  -43.2509,
  -43.2409,
  -43.2325,
  -43.2245,
  -43.2166,
  -43.2083,
  -43.1997,
  -43.1905,
  -43.1806,
  -43.1706,
  -43.1609,
  -43.1511,
  -43.1437,
  -43.1381,
  -43.1343,
  -43.1319,
  -43.1304,
  -43.1298,
  -43.1299,
  -43.1303,
  -43.1307,
  -43.1314,
  -43.1322,
  -43.134,
  -43.1368,
  -43.1409,
  -43.1459,
  -43.1515,
  -43.1569,
  -43.1622,
  -43.167,
  -43.1715,
  -43.1754,
  -43.1792,
  -43.1828,
  -43.1866,
  -43.1907,
  -43.1952,
  -43.2007,
  -43.2064,
  -43.2116,
  -43.2149,
  -43.215,
  -43.2108,
  -43.2021,
  -43.1889,
  -43.1707,
  -43.1474,
  -43.1172,
  -43.0794,
  -43.0327,
  -42.9743,
  -42.9045,
  -42.8205,
  -42.7211,
  -42.606,
  -42.4757,
  -42.3326,
  -42.1808,
  -42.0259,
  -41.8746,
  -41.7319,
  -41.6013,
  -41.4838,
  -41.3793,
  -41.286,
  -41.2015,
  -41.1227,
  -41.0466,
  -41.001,
  -41.0471,
  -41.0941,
  -41.1416,
  -41.1891,
  -41.2365,
  -41.2834,
  -41.3304,
  -41.3771,
  -41.424,
  -41.4699,
  -41.5166,
  -41.5628,
  -41.6079,
  -41.6516,
  -41.6936,
  -41.7344,
  -41.7749,
  -41.8151,
  -41.8557,
  -41.8964,
  -41.9368,
  -41.9763,
  -42.0146,
  -42.0509,
  -42.0842,
  -42.1163,
  -42.1461,
  -42.1735,
  -42.1986,
  -42.2209,
  -42.2402,
  -42.2564,
  -42.2694,
  -42.2796,
  -42.2868,
  -42.2914,
  -42.2933,
  -42.2929,
  -42.2908,
  -42.2868,
  -42.2837,
  -42.2813,
  -42.2803,
  -42.2807,
  -42.2828,
  -42.2867,
  -42.2916,
  -42.2969,
  -42.3014,
  -42.3042,
  -42.3056,
  -42.3056,
  -42.3047,
  -42.304,
  -42.3037,
  -42.3037,
  -42.306,
  -42.3095,
  -42.3138,
  -42.3186,
  -42.3238,
  -42.3302,
  -42.338,
  -42.3475,
  -42.3584,
  -42.3704,
  -42.3829,
  -42.3952,
  -42.4067,
  -42.4176,
  -42.4281,
  -42.4385,
  -42.4483,
  -42.4604,
  -42.4734,
  -42.4874,
  -42.5018,
  -42.5166,
  -42.5321,
  -42.5476,
  -42.5632,
  -42.5784,
  -42.5927,
  -42.6066,
  -42.6202,
  -42.6337,
  -42.6471,
  -42.6611,
  -42.6762,
  -42.6928,
  -42.7099,
  -42.7294,
  -42.7503,
  -42.7726,
  -42.7958,
  -42.8199,
  -42.8443,
  -42.869,
  -42.8942,
  -42.9205,
  -42.9486,
  -42.9788,
  -43.01,
  -43.0417,
  -43.0734,
  -43.1038,
  -43.1324,
  -43.1584,
  -43.1819,
  -43.2024,
  -43.2226,
  -43.2421,
  -43.2615,
  -43.2812,
  -43.3012,
  -43.3215,
  -43.3423,
  -43.3627,
  -43.3825,
  -43.4012,
  -43.4185,
  -43.4342,
  -43.4486,
  -43.4618,
  -43.4745,
  -43.4867,
  -43.4988,
  -43.5114,
  -43.5244,
  -43.5369,
  -43.5504,
  -43.5638,
  -43.577,
  -43.5899,
  -43.6025,
  -43.6148,
  -43.6271,
  -43.639,
  -43.6507,
  -43.6625,
  -43.6744,
  -43.6867,
  -43.699,
  -43.7113,
  -43.7232,
  -43.7345,
  -43.7452,
  -43.7555,
  -43.7652,
  -43.7743,
  -43.782,
  -43.7908,
  -43.7992,
  -43.8071,
  -43.8146,
  -43.8212,
  -43.8269,
  -43.832,
  -43.8365,
  -43.8409,
  -43.8454,
  -43.8498,
  -43.8544,
  -43.8587,
  -43.8627,
  -43.8665,
  -43.8695,
  -43.8723,
  -43.8749,
  -43.8775,
  -43.8804,
  -43.8836,
  -43.887,
  -43.8907,
  -43.8928,
  -43.8948,
  -43.8951,
  -43.8937,
  -43.8909,
  -43.8871,
  -43.8824,
  -43.8776,
  -43.8728,
  -43.8671,
  -43.8609,
  -43.8538,
  -43.8458,
  -43.8363,
  -43.8259,
  -43.8142,
  -43.8017,
  -43.7878,
  -43.7728,
  -43.7574,
  -43.7418,
  -43.7266,
  -43.712,
  -43.6975,
  -43.683,
  -43.6687,
  -43.6536,
  -43.6397,
  -43.6259,
  -43.6126,
  -43.5998,
  -43.5876,
  -43.5762,
  -43.5651,
  -43.5548,
  -43.5448,
  -43.535,
  -43.5247,
  -43.5134,
  -43.5014,
  -43.4882,
  -43.4745,
  -43.4606,
  -43.4464,
  -43.4321,
  -43.4183,
  -43.4049,
  -43.3913,
  -43.3774,
  -43.3633,
  -43.3485,
  -43.3334,
  -43.3186,
  -43.3043,
  -43.2909,
  -43.2785,
  -43.2676,
  -43.2575,
  -43.25,
  -43.2438,
  -43.2382,
  -43.2327,
  -43.2268,
  -43.2205,
  -43.2132,
  -43.2054,
  -43.1974,
  -43.189,
  -43.1812,
  -43.1745,
  -43.1693,
  -43.1654,
  -43.1624,
  -43.1605,
  -43.1595,
  -43.1588,
  -43.1583,
  -43.1577,
  -43.1575,
  -43.1574,
  -43.1582,
  -43.1601,
  -43.1633,
  -43.1673,
  -43.1716,
  -43.176,
  -43.1802,
  -43.1839,
  -43.1867,
  -43.1889,
  -43.1906,
  -43.1923,
  -43.1939,
  -43.1945,
  -43.197,
  -43.2006,
  -43.2045,
  -43.2076,
  -43.2089,
  -43.2068,
  -43.2009,
  -43.1906,
  -43.1758,
  -43.1564,
  -43.1317,
  -43.1008,
  -43.062,
  -43.0147,
  -42.957,
  -42.8876,
  -42.8044,
  -42.7065,
  -42.5933,
  -42.4647,
  -42.3228,
  -42.1713,
  -42.0153,
  -41.8616,
  -41.7155,
  -41.581,
  -41.4595,
  -41.3516,
  -41.2556,
  -41.1696,
  -41.0903,
  -41.0148,
  -40.9385,
  -40.9852,
  -41.0327,
  -41.0806,
  -41.1281,
  -41.1744,
  -41.221,
  -41.2676,
  -41.3141,
  -41.361,
  -41.408,
  -41.4549,
  -41.5013,
  -41.5466,
  -41.5904,
  -41.6329,
  -41.6741,
  -41.7148,
  -41.7554,
  -41.7961,
  -41.8355,
  -41.8755,
  -41.914,
  -41.951,
  -41.9862,
  -42.0196,
  -42.0512,
  -42.0808,
  -42.1085,
  -42.1336,
  -42.1559,
  -42.175,
  -42.1909,
  -42.2037,
  -42.2135,
  -42.2194,
  -42.224,
  -42.2265,
  -42.227,
  -42.226,
  -42.2243,
  -42.2227,
  -42.2219,
  -42.222,
  -42.2231,
  -42.2256,
  -42.2294,
  -42.2342,
  -42.2393,
  -42.2438,
  -42.2473,
  -42.2484,
  -42.2495,
  -42.2502,
  -42.2512,
  -42.2533,
  -42.2564,
  -42.2609,
  -42.2663,
  -42.2723,
  -42.2782,
  -42.2842,
  -42.2913,
  -42.2996,
  -42.3098,
  -42.3212,
  -42.3333,
  -42.3445,
  -42.3564,
  -42.3672,
  -42.3772,
  -42.3872,
  -42.397,
  -42.4076,
  -42.4194,
  -42.4325,
  -42.4465,
  -42.4615,
  -42.477,
  -42.493,
  -42.5092,
  -42.5253,
  -42.5406,
  -42.5552,
  -42.5689,
  -42.5815,
  -42.595,
  -42.6084,
  -42.6219,
  -42.6368,
  -42.6531,
  -42.6712,
  -42.6906,
  -42.7114,
  -42.7334,
  -42.7563,
  -42.7799,
  -42.8041,
  -42.8283,
  -42.8528,
  -42.878,
  -42.905,
  -42.9333,
  -42.9622,
  -42.9928,
  -43.0236,
  -43.0534,
  -43.0817,
  -43.1071,
  -43.1295,
  -43.1496,
  -43.1683,
  -43.1862,
  -43.2045,
  -43.2232,
  -43.2424,
  -43.2619,
  -43.2817,
  -43.3014,
  -43.3204,
  -43.3383,
  -43.3549,
  -43.3702,
  -43.3833,
  -43.3965,
  -43.4086,
  -43.4204,
  -43.4321,
  -43.4439,
  -43.456,
  -43.4685,
  -43.481,
  -43.4936,
  -43.5059,
  -43.5182,
  -43.5301,
  -43.5424,
  -43.5545,
  -43.567,
  -43.5793,
  -43.5919,
  -43.6048,
  -43.6181,
  -43.6316,
  -43.6438,
  -43.6566,
  -43.6688,
  -43.6806,
  -43.6918,
  -43.7026,
  -43.7132,
  -43.7236,
  -43.7336,
  -43.7431,
  -43.7523,
  -43.7607,
  -43.7681,
  -43.775,
  -43.7813,
  -43.7871,
  -43.7928,
  -43.7984,
  -43.804,
  -43.8092,
  -43.8141,
  -43.8186,
  -43.8228,
  -43.8256,
  -43.8287,
  -43.8318,
  -43.8353,
  -43.8393,
  -43.8437,
  -43.8482,
  -43.8528,
  -43.8568,
  -43.8597,
  -43.861,
  -43.8607,
  -43.8589,
  -43.8558,
  -43.8522,
  -43.8482,
  -43.8437,
  -43.8385,
  -43.8328,
  -43.8263,
  -43.8189,
  -43.8102,
  -43.8003,
  -43.7896,
  -43.7777,
  -43.7635,
  -43.7492,
  -43.7345,
  -43.7199,
  -43.7058,
  -43.6916,
  -43.6776,
  -43.6637,
  -43.6499,
  -43.6363,
  -43.623,
  -43.6101,
  -43.598,
  -43.5866,
  -43.5758,
  -43.5651,
  -43.5549,
  -43.5451,
  -43.5354,
  -43.5257,
  -43.5152,
  -43.5041,
  -43.4922,
  -43.4794,
  -43.466,
  -43.452,
  -43.4374,
  -43.423,
  -43.4091,
  -43.3944,
  -43.3809,
  -43.3669,
  -43.3526,
  -43.338,
  -43.3233,
  -43.3091,
  -43.2961,
  -43.2842,
  -43.274,
  -43.2655,
  -43.2588,
  -43.2536,
  -43.2496,
  -43.2461,
  -43.2426,
  -43.239,
  -43.2346,
  -43.2293,
  -43.2232,
  -43.2166,
  -43.2095,
  -43.2027,
  -43.1965,
  -43.1912,
  -43.187,
  -43.1838,
  -43.1815,
  -43.1798,
  -43.1782,
  -43.1767,
  -43.1754,
  -43.1742,
  -43.1733,
  -43.1725,
  -43.174,
  -43.1764,
  -43.1797,
  -43.1832,
  -43.1869,
  -43.1902,
  -43.1927,
  -43.1944,
  -43.1953,
  -43.1958,
  -43.1956,
  -43.1949,
  -43.1944,
  -43.1949,
  -43.1964,
  -43.1983,
  -43.1993,
  -43.1986,
  -43.195,
  -43.1879,
  -43.1767,
  -43.1613,
  -43.1412,
  -43.1159,
  -43.0841,
  -43.0444,
  -42.9965,
  -42.9384,
  -42.8687,
  -42.786,
  -42.6892,
  -42.5774,
  -42.4506,
  -42.3105,
  -42.1598,
  -42.0038,
  -41.8487,
  -41.7002,
  -41.5621,
  -41.437,
  -41.3255,
  -41.2267,
  -41.1382,
  -41.0566,
  -40.9808,
  -40.866,
  -40.9124,
  -40.9607,
  -41.009,
  -41.0569,
  -41.1041,
  -41.1509,
  -41.1974,
  -41.2438,
  -41.2905,
  -41.3375,
  -41.3844,
  -41.4308,
  -41.4761,
  -41.5203,
  -41.5621,
  -41.6039,
  -41.6453,
  -41.6863,
  -41.7272,
  -41.7675,
  -41.8065,
  -41.8439,
  -41.8796,
  -41.9137,
  -41.9462,
  -41.9773,
  -42.0066,
  -42.0342,
  -42.0596,
  -42.0812,
  -42.1006,
  -42.1167,
  -42.1295,
  -42.1393,
  -42.1465,
  -42.1514,
  -42.1545,
  -42.1561,
  -42.1563,
  -42.1559,
  -42.156,
  -42.1566,
  -42.158,
  -42.1604,
  -42.1636,
  -42.1667,
  -42.1716,
  -42.1766,
  -42.1813,
  -42.1853,
  -42.1885,
  -42.1909,
  -42.1933,
  -42.1961,
  -42.2002,
  -42.2056,
  -42.2121,
  -42.2192,
  -42.2263,
  -42.2334,
  -42.2402,
  -42.2466,
  -42.2554,
  -42.2659,
  -42.2771,
  -42.2892,
  -42.3007,
  -42.3117,
  -42.322,
  -42.3315,
  -42.3409,
  -42.3504,
  -42.3607,
  -42.3724,
  -42.3851,
  -42.3993,
  -42.4144,
  -42.4304,
  -42.446,
  -42.4627,
  -42.4791,
  -42.4947,
  -42.5094,
  -42.5232,
  -42.5365,
  -42.5497,
  -42.563,
  -42.5768,
  -42.5916,
  -42.6077,
  -42.6257,
  -42.6452,
  -42.6657,
  -42.6871,
  -42.7094,
  -42.7322,
  -42.7544,
  -42.7781,
  -42.8018,
  -42.8262,
  -42.8521,
  -42.879,
  -42.9072,
  -42.9364,
  -42.966,
  -42.9951,
  -43.0224,
  -43.0471,
  -43.0686,
  -43.0875,
  -43.105,
  -43.1219,
  -43.1393,
  -43.1573,
  -43.1758,
  -43.1938,
  -43.2128,
  -43.2317,
  -43.2501,
  -43.2672,
  -43.2831,
  -43.2978,
  -43.3116,
  -43.3244,
  -43.3363,
  -43.3476,
  -43.3589,
  -43.3702,
  -43.3817,
  -43.3932,
  -43.405,
  -43.4163,
  -43.4278,
  -43.4393,
  -43.4511,
  -43.4629,
  -43.4746,
  -43.4872,
  -43.5001,
  -43.5133,
  -43.5271,
  -43.5413,
  -43.5555,
  -43.5695,
  -43.5829,
  -43.5959,
  -43.6084,
  -43.6207,
  -43.6325,
  -43.6443,
  -43.6562,
  -43.6677,
  -43.6784,
  -43.6886,
  -43.6979,
  -43.7062,
  -43.7139,
  -43.721,
  -43.727,
  -43.7338,
  -43.7404,
  -43.7468,
  -43.7528,
  -43.7586,
  -43.7639,
  -43.7691,
  -43.7737,
  -43.7782,
  -43.7825,
  -43.7873,
  -43.7922,
  -43.7974,
  -43.8026,
  -43.8078,
  -43.8124,
  -43.8161,
  -43.8183,
  -43.8191,
  -43.8184,
  -43.8162,
  -43.8136,
  -43.8106,
  -43.8056,
  -43.8009,
  -43.7956,
  -43.7897,
  -43.783,
  -43.7753,
  -43.7662,
  -43.7563,
  -43.7452,
  -43.7326,
  -43.7191,
  -43.7054,
  -43.6915,
  -43.6779,
  -43.6644,
  -43.6508,
  -43.6374,
  -43.6242,
  -43.6112,
  -43.5988,
  -43.5871,
  -43.5764,
  -43.5662,
  -43.5564,
  -43.5467,
  -43.5371,
  -43.5276,
  -43.5177,
  -43.5067,
  -43.4961,
  -43.4848,
  -43.473,
  -43.4607,
  -43.4474,
  -43.4336,
  -43.4193,
  -43.4053,
  -43.3913,
  -43.3776,
  -43.3639,
  -43.3499,
  -43.336,
  -43.3216,
  -43.3077,
  -43.2948,
  -43.283,
  -43.2733,
  -43.2654,
  -43.259,
  -43.2548,
  -43.2517,
  -43.2494,
  -43.2477,
  -43.2462,
  -43.2442,
  -43.2416,
  -43.2379,
  -43.2334,
  -43.2281,
  -43.2223,
  -43.2153,
  -43.2094,
  -43.2039,
  -43.1992,
  -43.1957,
  -43.1931,
  -43.1907,
  -43.1884,
  -43.1863,
  -43.1842,
  -43.1824,
  -43.181,
  -43.1806,
  -43.1813,
  -43.1831,
  -43.1857,
  -43.1888,
  -43.1917,
  -43.1941,
  -43.1961,
  -43.1972,
  -43.1974,
  -43.1966,
  -43.1948,
  -43.1923,
  -43.19,
  -43.1884,
  -43.1875,
  -43.1872,
  -43.1864,
  -43.1841,
  -43.1794,
  -43.1718,
  -43.1605,
  -43.1449,
  -43.1243,
  -43.0983,
  -43.0656,
  -43.0253,
  -42.9763,
  -42.9165,
  -42.8467,
  -42.7645,
  -42.6686,
  -42.5581,
  -42.4329,
  -42.2945,
  -42.1453,
  -41.9899,
  -41.8342,
  -41.6841,
  -41.5434,
  -41.4151,
  -41.3003,
  -41.1984,
  -41.1073,
  -41.0249,
  -40.9476,
  -40.7822,
  -40.8305,
  -40.8793,
  -40.928,
  -40.9767,
  -41.0241,
  -41.0709,
  -41.1179,
  -41.1644,
  -41.2112,
  -41.257,
  -41.3039,
  -41.35,
  -41.3956,
  -41.44,
  -41.4835,
  -41.5261,
  -41.5682,
  -41.6099,
  -41.6507,
  -41.6905,
  -41.7286,
  -41.7651,
  -41.7997,
  -41.8325,
  -41.8632,
  -41.8935,
  -41.9226,
  -41.95,
  -41.9756,
  -41.9983,
  -42.0182,
  -42.0346,
  -42.048,
  -42.0581,
  -42.066,
  -42.0717,
  -42.0756,
  -42.0779,
  -42.0794,
  -42.0797,
  -42.0813,
  -42.0836,
  -42.0865,
  -42.0903,
  -42.0948,
  -42.0998,
  -42.105,
  -42.1104,
  -42.1153,
  -42.1197,
  -42.1238,
  -42.1279,
  -42.1318,
  -42.1366,
  -42.1423,
  -42.1484,
  -42.1567,
  -42.1652,
  -42.1736,
  -42.1812,
  -42.1887,
  -42.1967,
  -42.2056,
  -42.216,
  -42.2274,
  -42.2387,
  -42.2497,
  -42.2602,
  -42.2697,
  -42.2788,
  -42.2879,
  -42.2976,
  -42.3067,
  -42.3179,
  -42.3304,
  -42.3441,
  -42.3592,
  -42.3754,
  -42.3924,
  -42.4098,
  -42.4264,
  -42.4424,
  -42.4571,
  -42.4709,
  -42.484,
  -42.4968,
  -42.51,
  -42.524,
  -42.5392,
  -42.5555,
  -42.5724,
  -42.5919,
  -42.6121,
  -42.6327,
  -42.6541,
  -42.676,
  -42.6982,
  -42.721,
  -42.7442,
  -42.7681,
  -42.7929,
  -42.8185,
  -42.8452,
  -42.8729,
  -42.9012,
  -42.9292,
  -42.9555,
  -42.979,
  -42.9998,
  -43.0167,
  -43.0332,
  -43.0493,
  -43.066,
  -43.0837,
  -43.1019,
  -43.1204,
  -43.139,
  -43.1571,
  -43.1745,
  -43.1909,
  -43.206,
  -43.22,
  -43.233,
  -43.2455,
  -43.2571,
  -43.2682,
  -43.2789,
  -43.2897,
  -43.3006,
  -43.3105,
  -43.3212,
  -43.3316,
  -43.3423,
  -43.3533,
  -43.3649,
  -43.377,
  -43.3896,
  -43.4026,
  -43.4161,
  -43.4299,
  -43.4443,
  -43.4592,
  -43.4739,
  -43.4884,
  -43.5025,
  -43.5159,
  -43.5289,
  -43.5417,
  -43.5548,
  -43.5679,
  -43.5798,
  -43.5923,
  -43.6044,
  -43.6156,
  -43.6257,
  -43.6346,
  -43.6429,
  -43.6506,
  -43.6583,
  -43.6658,
  -43.6732,
  -43.6804,
  -43.6874,
  -43.6943,
  -43.7011,
  -43.7076,
  -43.7137,
  -43.7197,
  -43.7256,
  -43.7314,
  -43.7373,
  -43.7434,
  -43.7491,
  -43.7549,
  -43.7591,
  -43.7635,
  -43.7665,
  -43.7683,
  -43.7686,
  -43.7676,
  -43.7659,
  -43.7635,
  -43.7605,
  -43.7567,
  -43.7522,
  -43.7471,
  -43.7413,
  -43.7344,
  -43.7267,
  -43.7176,
  -43.7072,
  -43.6956,
  -43.6834,
  -43.6705,
  -43.6572,
  -43.6439,
  -43.6308,
  -43.6177,
  -43.6049,
  -43.5921,
  -43.5789,
  -43.5676,
  -43.5571,
  -43.5477,
  -43.5386,
  -43.5299,
  -43.5206,
  -43.5114,
  -43.5019,
  -43.4918,
  -43.4813,
  -43.4704,
  -43.459,
  -43.4473,
  -43.4349,
  -43.4222,
  -43.409,
  -43.3955,
  -43.3818,
  -43.3679,
  -43.3543,
  -43.3407,
  -43.3271,
  -43.3134,
  -43.3001,
  -43.2873,
  -43.2757,
  -43.266,
  -43.2581,
  -43.2526,
  -43.248,
  -43.2454,
  -43.2437,
  -43.243,
  -43.2426,
  -43.2424,
  -43.2417,
  -43.2404,
  -43.2382,
  -43.2352,
  -43.2314,
  -43.2269,
  -43.2216,
  -43.2158,
  -43.2101,
  -43.2053,
  -43.2014,
  -43.1982,
  -43.1954,
  -43.1929,
  -43.1904,
  -43.188,
  -43.1858,
  -43.184,
  -43.1827,
  -43.1827,
  -43.1838,
  -43.1857,
  -43.1881,
  -43.1901,
  -43.1919,
  -43.1932,
  -43.1939,
  -43.1935,
  -43.1917,
  -43.1888,
  -43.1851,
  -43.1802,
  -43.1766,
  -43.1736,
  -43.1711,
  -43.1686,
  -43.165,
  -43.1599,
  -43.1522,
  -43.1411,
  -43.1256,
  -43.1051,
  -43.0785,
  -43.0449,
  -43.0036,
  -42.9537,
  -42.8943,
  -42.8243,
  -42.7422,
  -42.6472,
  -42.5378,
  -42.4143,
  -42.2774,
  -42.1299,
  -41.9756,
  -41.8202,
  -41.6689,
  -41.5265,
  -41.3956,
  -41.278,
  -41.1731,
  -41.0795,
  -40.995,
  -40.9164,
  -40.6893,
  -40.7381,
  -40.7879,
  -40.8373,
  -40.8863,
  -40.9339,
  -40.9811,
  -41.028,
  -41.0748,
  -41.1217,
  -41.1686,
  -41.215,
  -41.2612,
  -41.3069,
  -41.3517,
  -41.3957,
  -41.4393,
  -41.4822,
  -41.5244,
  -41.5653,
  -41.6035,
  -41.6408,
  -41.6763,
  -41.7098,
  -41.7417,
  -41.7724,
  -41.8021,
  -41.8307,
  -41.8579,
  -41.8832,
  -41.9064,
  -41.9266,
  -41.9437,
  -41.9576,
  -41.9687,
  -41.9763,
  -41.9828,
  -41.9875,
  -41.9911,
  -41.9938,
  -41.9965,
  -41.9999,
  -42.0038,
  -42.0087,
  -42.0145,
  -42.0205,
  -42.0267,
  -42.0327,
  -42.0384,
  -42.0439,
  -42.049,
  -42.0531,
  -42.0585,
  -42.0641,
  -42.0703,
  -42.0774,
  -42.0858,
  -42.0953,
  -42.1053,
  -42.1144,
  -42.1228,
  -42.1305,
  -42.1387,
  -42.148,
  -42.1581,
  -42.169,
  -42.18,
  -42.1895,
  -42.1993,
  -42.2083,
  -42.217,
  -42.2259,
  -42.2355,
  -42.2458,
  -42.2568,
  -42.2691,
  -42.2826,
  -42.2976,
  -42.314,
  -42.3314,
  -42.349,
  -42.3661,
  -42.382,
  -42.3967,
  -42.4104,
  -42.4222,
  -42.435,
  -42.4481,
  -42.4625,
  -42.4782,
  -42.4948,
  -42.5128,
  -42.532,
  -42.5519,
  -42.572,
  -42.5926,
  -42.6132,
  -42.6348,
  -42.6568,
  -42.6797,
  -42.703,
  -42.7272,
  -42.7519,
  -42.7765,
  -42.803,
  -42.8297,
  -42.8566,
  -42.8822,
  -42.9044,
  -42.9242,
  -42.9414,
  -42.9568,
  -42.9724,
  -42.9886,
  -43.0058,
  -43.0237,
  -43.042,
  -43.06,
  -43.0773,
  -43.0937,
  -43.1092,
  -43.1234,
  -43.1365,
  -43.1476,
  -43.1593,
  -43.1705,
  -43.1814,
  -43.1919,
  -43.2022,
  -43.2125,
  -43.2227,
  -43.2326,
  -43.2425,
  -43.2526,
  -43.2632,
  -43.2747,
  -43.2869,
  -43.2999,
  -43.3133,
  -43.3272,
  -43.3416,
  -43.3565,
  -43.3718,
  -43.387,
  -43.4008,
  -43.4152,
  -43.429,
  -43.4425,
  -43.4558,
  -43.4694,
  -43.4833,
  -43.4972,
  -43.5108,
  -43.5239,
  -43.536,
  -43.5467,
  -43.5562,
  -43.5646,
  -43.5726,
  -43.5807,
  -43.5887,
  -43.5966,
  -43.6047,
  -43.613,
  -43.6211,
  -43.6294,
  -43.6377,
  -43.6447,
  -43.6527,
  -43.6603,
  -43.6677,
  -43.6747,
  -43.6815,
  -43.688,
  -43.6941,
  -43.6996,
  -43.7044,
  -43.7083,
  -43.7108,
  -43.7121,
  -43.7121,
  -43.7113,
  -43.71,
  -43.708,
  -43.7054,
  -43.7022,
  -43.6982,
  -43.6934,
  -43.6877,
  -43.6812,
  -43.6732,
  -43.6638,
  -43.6526,
  -43.6414,
  -43.6293,
  -43.6169,
  -43.6042,
  -43.5915,
  -43.5787,
  -43.5661,
  -43.5539,
  -43.5425,
  -43.5322,
  -43.5228,
  -43.5142,
  -43.5063,
  -43.4982,
  -43.4897,
  -43.4803,
  -43.4705,
  -43.4602,
  -43.4494,
  -43.4382,
  -43.4267,
  -43.4148,
  -43.4029,
  -43.3909,
  -43.3786,
  -43.3659,
  -43.3526,
  -43.3394,
  -43.3249,
  -43.3117,
  -43.2987,
  -43.2859,
  -43.2739,
  -43.2625,
  -43.2526,
  -43.245,
  -43.2394,
  -43.2358,
  -43.2339,
  -43.2328,
  -43.2324,
  -43.2327,
  -43.2332,
  -43.2336,
  -43.2339,
  -43.2336,
  -43.2328,
  -43.2312,
  -43.2289,
  -43.2253,
  -43.2207,
  -43.2152,
  -43.2097,
  -43.2048,
  -43.2006,
  -43.197,
  -43.1942,
  -43.1916,
  -43.1893,
  -43.1868,
  -43.1843,
  -43.1821,
  -43.179,
  -43.1781,
  -43.1783,
  -43.1793,
  -43.1804,
  -43.1817,
  -43.1828,
  -43.1838,
  -43.1839,
  -43.1828,
  -43.1804,
  -43.1772,
  -43.1727,
  -43.1677,
  -43.1626,
  -43.1576,
  -43.1532,
  -43.149,
  -43.1445,
  -43.1388,
  -43.1313,
  -43.1206,
  -43.1055,
  -43.0848,
  -43.0578,
  -43.0234,
  -42.9813,
  -42.9306,
  -42.8707,
  -42.8004,
  -42.7188,
  -42.6245,
  -42.5165,
  -42.3946,
  -42.2597,
  -42.114,
  -41.961,
  -41.8061,
  -41.6543,
  -41.5103,
  -41.3773,
  -41.2571,
  -41.1498,
  -41.0538,
  -40.9657,
  -40.8853,
  -40.5874,
  -40.6362,
  -40.6867,
  -40.7371,
  -40.787,
  -40.8357,
  -40.8833,
  -40.9303,
  -40.9772,
  -41.0239,
  -41.0705,
  -41.1169,
  -41.1631,
  -41.2089,
  -41.2542,
  -41.298,
  -41.3424,
  -41.386,
  -41.4285,
  -41.4693,
  -41.5079,
  -41.5447,
  -41.5791,
  -41.6118,
  -41.643,
  -41.6731,
  -41.702,
  -41.7301,
  -41.7571,
  -41.7824,
  -41.8045,
  -41.825,
  -41.8426,
  -41.8572,
  -41.8691,
  -41.8789,
  -41.8865,
  -41.8923,
  -41.8969,
  -41.9012,
  -41.9054,
  -41.9103,
  -41.9163,
  -41.9229,
  -41.9306,
  -41.9385,
  -41.9452,
  -41.9524,
  -41.9591,
  -41.965,
  -41.9711,
  -41.9772,
  -41.9837,
  -41.9906,
  -41.9983,
  -42.0065,
  -42.0159,
  -42.0261,
  -42.0366,
  -42.0466,
  -42.0553,
  -42.0634,
  -42.0708,
  -42.0801,
  -42.0902,
  -42.1009,
  -42.1114,
  -42.1212,
  -42.1303,
  -42.1389,
  -42.1472,
  -42.1562,
  -42.1661,
  -42.1767,
  -42.188,
  -42.2004,
  -42.2137,
  -42.2287,
  -42.2452,
  -42.2617,
  -42.2795,
  -42.2967,
  -42.3124,
  -42.3269,
  -42.3407,
  -42.3536,
  -42.3666,
  -42.3802,
  -42.3947,
  -42.4107,
  -42.428,
  -42.4461,
  -42.4652,
  -42.4847,
  -42.5045,
  -42.5244,
  -42.5449,
  -42.5648,
  -42.5862,
  -42.6085,
  -42.6315,
  -42.6554,
  -42.6797,
  -42.7041,
  -42.7294,
  -42.7552,
  -42.7809,
  -42.805,
  -42.8271,
  -42.8453,
  -42.8618,
  -42.8766,
  -42.8917,
  -42.9071,
  -42.9239,
  -42.9415,
  -42.9582,
  -42.9757,
  -42.9923,
  -43.0077,
  -43.0221,
  -43.0353,
  -43.0473,
  -43.0584,
  -43.069,
  -43.0794,
  -43.09,
  -43.1002,
  -43.1102,
  -43.1198,
  -43.1293,
  -43.1388,
  -43.1482,
  -43.1581,
  -43.1687,
  -43.1803,
  -43.1925,
  -43.2047,
  -43.2186,
  -43.2331,
  -43.248,
  -43.2634,
  -43.279,
  -43.2943,
  -43.3093,
  -43.324,
  -43.3382,
  -43.3518,
  -43.3656,
  -43.3795,
  -43.3939,
  -43.4085,
  -43.4232,
  -43.437,
  -43.4496,
  -43.4607,
  -43.4703,
  -43.479,
  -43.4874,
  -43.4945,
  -43.5028,
  -43.5112,
  -43.5203,
  -43.5295,
  -43.5393,
  -43.5496,
  -43.5596,
  -43.5698,
  -43.5796,
  -43.5891,
  -43.5983,
  -43.6068,
  -43.6145,
  -43.6215,
  -43.6279,
  -43.6335,
  -43.6386,
  -43.643,
  -43.6461,
  -43.6482,
  -43.6493,
  -43.6495,
  -43.6491,
  -43.6476,
  -43.6465,
  -43.6448,
  -43.6423,
  -43.6389,
  -43.6342,
  -43.6292,
  -43.6225,
  -43.6146,
  -43.6057,
  -43.5957,
  -43.5847,
  -43.5732,
  -43.5611,
  -43.5487,
  -43.5361,
  -43.5237,
  -43.512,
  -43.5013,
  -43.4915,
  -43.4829,
  -43.4754,
  -43.4682,
  -43.4605,
  -43.4522,
  -43.4429,
  -43.4329,
  -43.4227,
  -43.4109,
  -43.3996,
  -43.388,
  -43.3763,
  -43.3648,
  -43.3536,
  -43.3422,
  -43.3303,
  -43.3179,
  -43.3052,
  -43.2923,
  -43.2799,
  -43.2678,
  -43.2562,
  -43.2454,
  -43.2358,
  -43.2281,
  -43.2225,
  -43.2189,
  -43.2173,
  -43.2165,
  -43.2165,
  -43.2169,
  -43.2176,
  -43.2184,
  -43.2192,
  -43.22,
  -43.2205,
  -43.2209,
  -43.2206,
  -43.2196,
  -43.217,
  -43.2121,
  -43.2073,
  -43.2022,
  -43.1974,
  -43.1933,
  -43.1897,
  -43.1871,
  -43.1848,
  -43.1827,
  -43.1805,
  -43.178,
  -43.1751,
  -43.1726,
  -43.1705,
  -43.1694,
  -43.1688,
  -43.1688,
  -43.1691,
  -43.1696,
  -43.1698,
  -43.1691,
  -43.1675,
  -43.1652,
  -43.1617,
  -43.1571,
  -43.1517,
  -43.1455,
  -43.1391,
  -43.1332,
  -43.1277,
  -43.1222,
  -43.1161,
  -43.1086,
  -43.0981,
  -43.0832,
  -43.0623,
  -43.0346,
  -42.9997,
  -42.9565,
  -42.9053,
  -42.844,
  -42.7741,
  -42.6931,
  -42.5999,
  -42.4934,
  -42.3735,
  -42.2408,
  -42.0972,
  -41.9458,
  -41.7916,
  -41.6396,
  -41.4944,
  -41.3595,
  -41.2371,
  -41.1271,
  -41.0286,
  -40.9395,
  -40.8574,
  -40.4759,
  -40.5268,
  -40.5783,
  -40.6297,
  -40.6802,
  -40.7292,
  -40.7771,
  -40.8241,
  -40.8707,
  -40.9171,
  -40.9625,
  -41.0087,
  -41.055,
  -41.1012,
  -41.1472,
  -41.1928,
  -41.2377,
  -41.2815,
  -41.324,
  -41.3643,
  -41.4026,
  -41.4386,
  -41.4727,
  -41.5047,
  -41.5357,
  -41.5643,
  -41.5929,
  -41.6204,
  -41.647,
  -41.6722,
  -41.6953,
  -41.7159,
  -41.7341,
  -41.7495,
  -41.7625,
  -41.7731,
  -41.7817,
  -41.7888,
  -41.7948,
  -41.8005,
  -41.8054,
  -41.8121,
  -41.8198,
  -41.8284,
  -41.8378,
  -41.8473,
  -41.8567,
  -41.8653,
  -41.8729,
  -41.8801,
  -41.8869,
  -41.8941,
  -41.9017,
  -41.9099,
  -41.9186,
  -41.9278,
  -41.9367,
  -41.9473,
  -41.9579,
  -41.9679,
  -41.9768,
  -41.9851,
  -41.9938,
  -42.0034,
  -42.0137,
  -42.024,
  -42.0341,
  -42.0434,
  -42.0518,
  -42.0603,
  -42.0688,
  -42.078,
  -42.0882,
  -42.0986,
  -42.1107,
  -42.1233,
  -42.1369,
  -42.152,
  -42.1685,
  -42.1859,
  -42.2036,
  -42.2206,
  -42.2362,
  -42.2509,
  -42.2645,
  -42.2779,
  -42.2911,
  -42.3053,
  -42.3205,
  -42.3369,
  -42.3546,
  -42.3722,
  -42.3912,
  -42.4106,
  -42.4302,
  -42.4501,
  -42.4701,
  -42.4906,
  -42.5116,
  -42.5335,
  -42.5566,
  -42.5801,
  -42.6041,
  -42.6282,
  -42.6525,
  -42.6772,
  -42.7018,
  -42.725,
  -42.746,
  -42.7636,
  -42.7779,
  -42.792,
  -42.8064,
  -42.8217,
  -42.838,
  -42.8548,
  -42.8722,
  -42.8889,
  -42.9046,
  -42.9191,
  -42.9324,
  -42.9444,
  -42.9552,
  -42.9652,
  -42.9747,
  -42.984,
  -42.9935,
  -43.0032,
  -43.0128,
  -43.022,
  -43.0299,
  -43.0391,
  -43.0483,
  -43.058,
  -43.0688,
  -43.0803,
  -43.093,
  -43.1067,
  -43.1212,
  -43.1362,
  -43.1516,
  -43.1672,
  -43.1829,
  -43.1983,
  -43.2137,
  -43.2285,
  -43.2429,
  -43.2572,
  -43.2711,
  -43.2853,
  -43.2999,
  -43.314,
  -43.3288,
  -43.3432,
  -43.356,
  -43.3672,
  -43.3771,
  -43.3859,
  -43.3947,
  -43.4033,
  -43.412,
  -43.4207,
  -43.4304,
  -43.4408,
  -43.4524,
  -43.464,
  -43.4758,
  -43.4882,
  -43.5001,
  -43.5118,
  -43.5226,
  -43.5327,
  -43.5415,
  -43.5489,
  -43.5554,
  -43.5602,
  -43.5655,
  -43.5702,
  -43.574,
  -43.5767,
  -43.5785,
  -43.5798,
  -43.5808,
  -43.582,
  -43.5826,
  -43.5826,
  -43.5818,
  -43.5796,
  -43.577,
  -43.5733,
  -43.5682,
  -43.5617,
  -43.5541,
  -43.5455,
  -43.5357,
  -43.5252,
  -43.5137,
  -43.5017,
  -43.4893,
  -43.4771,
  -43.4656,
  -43.4542,
  -43.4449,
  -43.4368,
  -43.4299,
  -43.4231,
  -43.4158,
  -43.4076,
  -43.3985,
  -43.3888,
  -43.3787,
  -43.3681,
  -43.357,
  -43.3456,
  -43.3343,
  -43.3236,
  -43.313,
  -43.3023,
  -43.2914,
  -43.28,
  -43.2679,
  -43.256,
  -43.2445,
  -43.2333,
  -43.223,
  -43.2137,
  -43.2061,
  -43.2005,
  -43.197,
  -43.1953,
  -43.195,
  -43.1943,
  -43.195,
  -43.1959,
  -43.1968,
  -43.1975,
  -43.1984,
  -43.1994,
  -43.2007,
  -43.2018,
  -43.2028,
  -43.2028,
  -43.2014,
  -43.1985,
  -43.1946,
  -43.1903,
  -43.1858,
  -43.182,
  -43.1789,
  -43.1764,
  -43.1745,
  -43.1731,
  -43.1712,
  -43.1685,
  -43.1656,
  -43.1624,
  -43.1591,
  -43.1562,
  -43.154,
  -43.1527,
  -43.1519,
  -43.1512,
  -43.1503,
  -43.1489,
  -43.1472,
  -43.1449,
  -43.1417,
  -43.1375,
  -43.131,
  -43.1243,
  -43.1171,
  -43.1102,
  -43.1037,
  -43.0973,
  -43.0907,
  -43.0829,
  -43.0724,
  -43.0575,
  -43.0361,
  -43.0078,
  -42.9722,
  -42.9284,
  -42.8772,
  -42.8171,
  -42.7473,
  -42.6672,
  -42.5752,
  -42.4706,
  -42.3531,
  -42.223,
  -42.0818,
  -41.9324,
  -41.7792,
  -41.6273,
  -41.4812,
  -41.3447,
  -41.22,
  -41.1075,
  -41.0066,
  -40.9154,
  -40.8316,
  -40.3579,
  -40.4098,
  -40.4623,
  -40.5144,
  -40.5655,
  -40.614,
  -40.6617,
  -40.7085,
  -40.7548,
  -40.8008,
  -40.847,
  -40.8934,
  -40.94,
  -40.9866,
  -41.0331,
  -41.0793,
  -41.1245,
  -41.1683,
  -41.2103,
  -41.2498,
  -41.2864,
  -41.3219,
  -41.3555,
  -41.3877,
  -41.4184,
  -41.4482,
  -41.4767,
  -41.504,
  -41.5304,
  -41.5554,
  -41.5784,
  -41.5994,
  -41.6179,
  -41.6341,
  -41.6479,
  -41.6583,
  -41.6681,
  -41.6763,
  -41.6839,
  -41.6913,
  -41.699,
  -41.7074,
  -41.7167,
  -41.7271,
  -41.738,
  -41.7488,
  -41.7595,
  -41.7694,
  -41.7786,
  -41.7869,
  -41.7949,
  -41.802,
  -41.8109,
  -41.8203,
  -41.8301,
  -41.8403,
  -41.8507,
  -41.8607,
  -41.8707,
  -41.8806,
  -41.8896,
  -41.8982,
  -41.9073,
  -41.917,
  -41.9275,
  -41.9379,
  -41.9477,
  -41.9557,
  -41.9642,
  -41.9723,
  -41.9811,
  -41.991,
  -42.0018,
  -42.014,
  -42.0268,
  -42.0404,
  -42.0546,
  -42.0699,
  -42.0863,
  -42.1036,
  -42.121,
  -42.1378,
  -42.1536,
  -42.1682,
  -42.1821,
  -42.1949,
  -42.2092,
  -42.2241,
  -42.24,
  -42.257,
  -42.2749,
  -42.2937,
  -42.3131,
  -42.3326,
  -42.3522,
  -42.3722,
  -42.3924,
  -42.4127,
  -42.4336,
  -42.4553,
  -42.4778,
  -42.5011,
  -42.5251,
  -42.5479,
  -42.5717,
  -42.5955,
  -42.6191,
  -42.6412,
  -42.6609,
  -42.678,
  -42.6927,
  -42.7064,
  -42.72,
  -42.7346,
  -42.7503,
  -42.7667,
  -42.7833,
  -42.7993,
  -42.8143,
  -42.8277,
  -42.8398,
  -42.8505,
  -42.8601,
  -42.8677,
  -42.8761,
  -42.8841,
  -42.8924,
  -42.9009,
  -42.9097,
  -42.9185,
  -42.9269,
  -42.9357,
  -42.945,
  -42.9547,
  -42.9654,
  -42.9771,
  -42.9903,
  -43.0045,
  -43.0194,
  -43.035,
  -43.0507,
  -43.0667,
  -43.0826,
  -43.0983,
  -43.1129,
  -43.1281,
  -43.1429,
  -43.1574,
  -43.1716,
  -43.1861,
  -43.2007,
  -43.2157,
  -43.2307,
  -43.245,
  -43.2578,
  -43.2693,
  -43.2793,
  -43.2886,
  -43.2976,
  -43.3069,
  -43.316,
  -43.3253,
  -43.3355,
  -43.347,
  -43.3595,
  -43.3724,
  -43.3862,
  -43.3994,
  -43.4137,
  -43.4271,
  -43.4399,
  -43.4513,
  -43.4608,
  -43.4689,
  -43.4758,
  -43.4818,
  -43.4874,
  -43.4924,
  -43.4967,
  -43.5001,
  -43.5028,
  -43.5052,
  -43.5077,
  -43.5106,
  -43.5131,
  -43.5151,
  -43.516,
  -43.516,
  -43.5148,
  -43.5125,
  -43.5089,
  -43.5038,
  -43.4967,
  -43.4893,
  -43.4809,
  -43.4712,
  -43.4607,
  -43.4493,
  -43.4373,
  -43.4254,
  -43.414,
  -43.4035,
  -43.3944,
  -43.3867,
  -43.3801,
  -43.3736,
  -43.3665,
  -43.3587,
  -43.3498,
  -43.3406,
  -43.3309,
  -43.3208,
  -43.3102,
  -43.2994,
  -43.2888,
  -43.2785,
  -43.2684,
  -43.2585,
  -43.2483,
  -43.2376,
  -43.2266,
  -43.2148,
  -43.2042,
  -43.1942,
  -43.1853,
  -43.1775,
  -43.1719,
  -43.1683,
  -43.1666,
  -43.1665,
  -43.1674,
  -43.1687,
  -43.17,
  -43.1711,
  -43.172,
  -43.1727,
  -43.1737,
  -43.1749,
  -43.1764,
  -43.1782,
  -43.1799,
  -43.1809,
  -43.1808,
  -43.1793,
  -43.1766,
  -43.1731,
  -43.1694,
  -43.1662,
  -43.1636,
  -43.1616,
  -43.1601,
  -43.159,
  -43.1572,
  -43.155,
  -43.1518,
  -43.1468,
  -43.1423,
  -43.138,
  -43.1344,
  -43.1317,
  -43.1292,
  -43.127,
  -43.1248,
  -43.1229,
  -43.1211,
  -43.1189,
  -43.1163,
  -43.1125,
  -43.1074,
  -43.1008,
  -43.0935,
  -43.0857,
  -43.0783,
  -43.0715,
  -43.0643,
  -43.0561,
  -43.0452,
  -43.0296,
  -43.0079,
  -42.979,
  -42.9427,
  -42.8989,
  -42.8474,
  -42.7876,
  -42.7188,
  -42.6396,
  -42.5493,
  -42.447,
  -42.3323,
  -42.2052,
  -42.067,
  -41.9198,
  -41.7681,
  -41.6166,
  -41.4701,
  -41.3322,
  -41.2055,
  -41.0905,
  -40.9875,
  -40.8931,
  -40.808,
  -40.2325,
  -40.2848,
  -40.3383,
  -40.3911,
  -40.4428,
  -40.4924,
  -40.5403,
  -40.5868,
  -40.6326,
  -40.6783,
  -40.7243,
  -40.7708,
  -40.8177,
  -40.8648,
  -40.9119,
  -40.9574,
  -41.0025,
  -41.0458,
  -41.0869,
  -41.1259,
  -41.1625,
  -41.1972,
  -41.2308,
  -41.263,
  -41.2942,
  -41.3242,
  -41.353,
  -41.3805,
  -41.4068,
  -41.4316,
  -41.4537,
  -41.4749,
  -41.4936,
  -41.5103,
  -41.5249,
  -41.5373,
  -41.548,
  -41.5576,
  -41.5667,
  -41.5759,
  -41.5857,
  -41.5956,
  -41.6066,
  -41.6181,
  -41.6302,
  -41.6422,
  -41.6528,
  -41.664,
  -41.6745,
  -41.6842,
  -41.6934,
  -41.7027,
  -41.7127,
  -41.7235,
  -41.7346,
  -41.7458,
  -41.7561,
  -41.766,
  -41.7752,
  -41.7842,
  -41.7932,
  -41.8023,
  -41.811,
  -41.8211,
  -41.8318,
  -41.8422,
  -41.852,
  -41.8609,
  -41.8696,
  -41.8781,
  -41.8872,
  -41.8977,
  -41.9095,
  -41.9224,
  -41.9362,
  -41.9507,
  -41.9658,
  -41.9816,
  -41.9984,
  -42.0145,
  -42.0317,
  -42.0482,
  -42.064,
  -42.0791,
  -42.0938,
  -42.1085,
  -42.1237,
  -42.1394,
  -42.1561,
  -42.1735,
  -42.192,
  -42.2111,
  -42.2309,
  -42.2507,
  -42.2706,
  -42.2906,
  -42.3111,
  -42.3305,
  -42.3513,
  -42.3728,
  -42.3951,
  -42.418,
  -42.4417,
  -42.4654,
  -42.489,
  -42.5121,
  -42.5346,
  -42.5558,
  -42.5749,
  -42.5911,
  -42.6056,
  -42.6187,
  -42.6316,
  -42.6454,
  -42.6603,
  -42.6762,
  -42.6912,
  -42.7065,
  -42.7205,
  -42.7329,
  -42.7438,
  -42.7533,
  -42.7615,
  -42.7689,
  -42.7758,
  -42.7824,
  -42.7892,
  -42.7965,
  -42.804,
  -42.812,
  -42.8202,
  -42.829,
  -42.8379,
  -42.8475,
  -42.8586,
  -42.8705,
  -42.8841,
  -42.8977,
  -42.9133,
  -42.9293,
  -42.9455,
  -42.9616,
  -42.9775,
  -42.9935,
  -43.0094,
  -43.025,
  -43.0404,
  -43.0554,
  -43.0699,
  -43.0844,
  -43.0989,
  -43.1134,
  -43.1281,
  -43.142,
  -43.1547,
  -43.1665,
  -43.1771,
  -43.1871,
  -43.1966,
  -43.205,
  -43.2145,
  -43.2243,
  -43.2351,
  -43.2471,
  -43.2604,
  -43.2746,
  -43.2901,
  -43.306,
  -43.3222,
  -43.3376,
  -43.352,
  -43.3644,
  -43.3749,
  -43.3838,
  -43.3912,
  -43.3977,
  -43.4037,
  -43.4093,
  -43.4141,
  -43.4183,
  -43.4219,
  -43.4256,
  -43.4296,
  -43.4331,
  -43.4376,
  -43.4415,
  -43.4444,
  -43.446,
  -43.4467,
  -43.4459,
  -43.4436,
  -43.4399,
  -43.435,
  -43.4289,
  -43.4217,
  -43.4133,
  -43.4038,
  -43.3934,
  -43.3821,
  -43.3706,
  -43.3593,
  -43.3489,
  -43.3399,
  -43.3323,
  -43.3256,
  -43.3193,
  -43.3126,
  -43.3053,
  -43.2971,
  -43.2884,
  -43.2792,
  -43.2687,
  -43.2589,
  -43.2488,
  -43.2389,
  -43.229,
  -43.2194,
  -43.2099,
  -43.2002,
  -43.1904,
  -43.1805,
  -43.1706,
  -43.1609,
  -43.1519,
  -43.1443,
  -43.1384,
  -43.1346,
  -43.1327,
  -43.1327,
  -43.134,
  -43.1359,
  -43.1381,
  -43.14,
  -43.1414,
  -43.1425,
  -43.1433,
  -43.1444,
  -43.1457,
  -43.1475,
  -43.1498,
  -43.1519,
  -43.1539,
  -43.154,
  -43.1538,
  -43.1522,
  -43.1499,
  -43.1473,
  -43.145,
  -43.1429,
  -43.1414,
  -43.14,
  -43.1391,
  -43.1378,
  -43.1356,
  -43.1321,
  -43.1276,
  -43.1223,
  -43.117,
  -43.1122,
  -43.1077,
  -43.1033,
  -43.0992,
  -43.0961,
  -43.0935,
  -43.0916,
  -43.0897,
  -43.0875,
  -43.0844,
  -43.0798,
  -43.0738,
  -43.0666,
  -43.0587,
  -43.0509,
  -43.0433,
  -43.0353,
  -43.0263,
  -43.0146,
  -42.9986,
  -42.9763,
  -42.947,
  -42.9102,
  -42.8663,
  -42.8141,
  -42.755,
  -42.6871,
  -42.6094,
  -42.5211,
  -42.4215,
  -42.3102,
  -42.1868,
  -42.0519,
  -41.9076,
  -41.7578,
  -41.6073,
  -41.4607,
  -41.3217,
  -41.193,
  -41.0758,
  -40.9703,
  -40.8758,
  -40.7895,
  -40.1005,
  -40.1545,
  -40.2087,
  -40.2623,
  -40.3143,
  -40.3643,
  -40.4123,
  -40.4588,
  -40.5045,
  -40.55,
  -40.5949,
  -40.6414,
  -40.6885,
  -40.7359,
  -40.783,
  -40.8295,
  -40.8743,
  -40.9169,
  -40.9572,
  -40.9951,
  -41.031,
  -41.0654,
  -41.0987,
  -41.1313,
  -41.1629,
  -41.1923,
  -41.2214,
  -41.249,
  -41.2752,
  -41.3,
  -41.3231,
  -41.3443,
  -41.3636,
  -41.3807,
  -41.3957,
  -41.4091,
  -41.421,
  -41.4319,
  -41.443,
  -41.454,
  -41.4644,
  -41.4757,
  -41.4881,
  -41.5007,
  -41.5136,
  -41.5266,
  -41.5392,
  -41.5514,
  -41.5629,
  -41.574,
  -41.5845,
  -41.5951,
  -41.6062,
  -41.6182,
  -41.6306,
  -41.6424,
  -41.6526,
  -41.6623,
  -41.6712,
  -41.6798,
  -41.6885,
  -41.6981,
  -41.7083,
  -41.719,
  -41.7299,
  -41.7404,
  -41.7503,
  -41.7597,
  -41.7687,
  -41.778,
  -41.7877,
  -41.7987,
  -41.811,
  -41.8238,
  -41.8384,
  -41.8537,
  -41.8699,
  -41.8865,
  -41.9038,
  -41.9209,
  -41.9382,
  -41.9549,
  -41.9711,
  -41.9869,
  -42.0026,
  -42.0183,
  -42.0343,
  -42.0506,
  -42.0679,
  -42.0861,
  -42.1051,
  -42.1238,
  -42.1439,
  -42.1641,
  -42.1846,
  -42.2048,
  -42.2253,
  -42.2463,
  -42.2671,
  -42.2887,
  -42.3107,
  -42.3333,
  -42.3565,
  -42.3801,
  -42.4035,
  -42.4264,
  -42.4479,
  -42.468,
  -42.4867,
  -42.5026,
  -42.5155,
  -42.5282,
  -42.5405,
  -42.5535,
  -42.5678,
  -42.5827,
  -42.5981,
  -42.6126,
  -42.6255,
  -42.6369,
  -42.6465,
  -42.6547,
  -42.6618,
  -42.6679,
  -42.6735,
  -42.6785,
  -42.6839,
  -42.6896,
  -42.6959,
  -42.7029,
  -42.7097,
  -42.7182,
  -42.7271,
  -42.737,
  -42.7479,
  -42.7601,
  -42.7739,
  -42.789,
  -42.805,
  -42.8216,
  -42.838,
  -42.8542,
  -42.8702,
  -42.8863,
  -42.9023,
  -42.9183,
  -42.9339,
  -42.9491,
  -42.964,
  -42.9784,
  -42.9929,
  -43.0061,
  -43.0203,
  -43.0339,
  -43.0468,
  -43.0588,
  -43.0702,
  -43.0808,
  -43.0909,
  -43.1007,
  -43.1107,
  -43.1208,
  -43.1318,
  -43.1442,
  -43.1578,
  -43.173,
  -43.1895,
  -43.2069,
  -43.2245,
  -43.2416,
  -43.2572,
  -43.271,
  -43.2828,
  -43.2927,
  -43.3009,
  -43.3071,
  -43.3139,
  -43.32,
  -43.3257,
  -43.3308,
  -43.3357,
  -43.3406,
  -43.3463,
  -43.3525,
  -43.3584,
  -43.3639,
  -43.3685,
  -43.3722,
  -43.3744,
  -43.375,
  -43.3743,
  -43.3719,
  -43.3684,
  -43.3636,
  -43.3577,
  -43.3507,
  -43.3425,
  -43.3332,
  -43.3228,
  -43.3119,
  -43.3011,
  -43.2901,
  -43.2812,
  -43.2736,
  -43.267,
  -43.2608,
  -43.2546,
  -43.2478,
  -43.2403,
  -43.2321,
  -43.2235,
  -43.2146,
  -43.2055,
  -43.1962,
  -43.1869,
  -43.1775,
  -43.1682,
  -43.159,
  -43.1497,
  -43.1406,
  -43.1314,
  -43.1221,
  -43.1132,
  -43.1055,
  -43.0993,
  -43.095,
  -43.0929,
  -43.0927,
  -43.0941,
  -43.0965,
  -43.0998,
  -43.1019,
  -43.1042,
  -43.1061,
  -43.1075,
  -43.1087,
  -43.1099,
  -43.1115,
  -43.1136,
  -43.116,
  -43.1189,
  -43.1214,
  -43.1235,
  -43.1245,
  -43.124,
  -43.1227,
  -43.1214,
  -43.1197,
  -43.1182,
  -43.117,
  -43.1161,
  -43.1153,
  -43.1143,
  -43.1119,
  -43.1082,
  -43.1035,
  -43.0979,
  -43.0918,
  -43.0856,
  -43.0791,
  -43.073,
  -43.0676,
  -43.0632,
  -43.06,
  -43.0578,
  -43.0562,
  -43.0545,
  -43.0521,
  -43.0474,
  -43.042,
  -43.0352,
  -43.0276,
  -43.0196,
  -43.0113,
  -43.0026,
  -42.9925,
  -42.9799,
  -42.9629,
  -42.9401,
  -42.9104,
  -42.8737,
  -42.83,
  -42.7794,
  -42.7212,
  -42.6544,
  -42.5787,
  -42.493,
  -42.3965,
  -42.2888,
  -42.1694,
  -42.0383,
  -41.8974,
  -41.7501,
  -41.6011,
  -41.4549,
  -41.3154,
  -41.1852,
  -41.0666,
  -40.9594,
  -40.8632,
  -40.7765,
  -39.9646,
  -40.019,
  -40.0736,
  -40.1276,
  -40.1801,
  -40.2296,
  -40.278,
  -40.3245,
  -40.3703,
  -40.4157,
  -40.4615,
  -40.5078,
  -40.5548,
  -40.6021,
  -40.6492,
  -40.6953,
  -40.7395,
  -40.7812,
  -40.8206,
  -40.8578,
  -40.892,
  -40.9262,
  -40.9596,
  -40.9925,
  -41.0245,
  -41.0553,
  -41.0846,
  -41.1123,
  -41.1385,
  -41.1633,
  -41.1865,
  -41.2078,
  -41.2274,
  -41.2451,
  -41.2607,
  -41.2739,
  -41.2869,
  -41.2996,
  -41.3123,
  -41.3248,
  -41.3375,
  -41.3505,
  -41.3638,
  -41.3773,
  -41.3911,
  -41.4048,
  -41.4183,
  -41.4313,
  -41.4438,
  -41.456,
  -41.4677,
  -41.4785,
  -41.4908,
  -41.504,
  -41.5175,
  -41.5304,
  -41.5422,
  -41.5524,
  -41.5614,
  -41.57,
  -41.579,
  -41.5887,
  -41.5994,
  -41.6107,
  -41.6218,
  -41.6325,
  -41.6428,
  -41.6516,
  -41.6614,
  -41.6713,
  -41.6821,
  -41.6935,
  -41.7061,
  -41.7205,
  -41.7359,
  -41.7522,
  -41.7692,
  -41.787,
  -41.805,
  -41.8226,
  -41.8402,
  -41.8574,
  -41.8745,
  -41.8913,
  -41.9081,
  -41.9237,
  -41.9404,
  -41.9571,
  -41.9748,
  -41.9936,
  -42.0134,
  -42.0339,
  -42.0546,
  -42.0754,
  -42.0964,
  -42.1171,
  -42.1376,
  -42.1585,
  -42.1798,
  -42.2014,
  -42.2232,
  -42.2455,
  -42.2684,
  -42.2907,
  -42.3139,
  -42.3366,
  -42.3583,
  -42.378,
  -42.3957,
  -42.4114,
  -42.425,
  -42.4372,
  -42.449,
  -42.4615,
  -42.4746,
  -42.4888,
  -42.503,
  -42.5163,
  -42.5283,
  -42.5386,
  -42.5469,
  -42.5541,
  -42.5601,
  -42.5641,
  -42.5685,
  -42.5723,
  -42.576,
  -42.5804,
  -42.5856,
  -42.5916,
  -42.5987,
  -42.607,
  -42.6161,
  -42.626,
  -42.637,
  -42.6495,
  -42.6634,
  -42.6788,
  -42.6949,
  -42.7115,
  -42.728,
  -42.7444,
  -42.7604,
  -42.7763,
  -42.7915,
  -42.8074,
  -42.8231,
  -42.8386,
  -42.8539,
  -42.8686,
  -42.883,
  -42.8968,
  -42.9104,
  -42.9235,
  -42.9364,
  -42.949,
  -42.9611,
  -42.9726,
  -42.9835,
  -42.9936,
  -43.0039,
  -43.0142,
  -43.0253,
  -43.0376,
  -43.0512,
  -43.067,
  -43.0844,
  -43.1018,
  -43.1204,
  -43.1386,
  -43.1557,
  -43.1709,
  -43.1841,
  -43.1952,
  -43.2046,
  -43.2129,
  -43.2205,
  -43.2276,
  -43.2342,
  -43.2404,
  -43.2464,
  -43.2531,
  -43.2602,
  -43.2677,
  -43.2751,
  -43.2821,
  -43.2885,
  -43.2935,
  -43.2976,
  -43.3,
  -43.3008,
  -43.2999,
  -43.2969,
  -43.2933,
  -43.2888,
  -43.2832,
  -43.2762,
  -43.268,
  -43.2588,
  -43.2488,
  -43.239,
  -43.2293,
  -43.221,
  -43.2136,
  -43.207,
  -43.201,
  -43.1951,
  -43.1888,
  -43.1816,
  -43.1739,
  -43.1659,
  -43.1578,
  -43.1496,
  -43.141,
  -43.1323,
  -43.1234,
  -43.1143,
  -43.1052,
  -43.0963,
  -43.0874,
  -43.0774,
  -43.0687,
  -43.0609,
  -43.0543,
  -43.0496,
  -43.0469,
  -43.0462,
  -43.0473,
  -43.0499,
  -43.0538,
  -43.058,
  -43.0615,
  -43.0646,
  -43.0672,
  -43.0696,
  -43.0715,
  -43.0732,
  -43.0753,
  -43.0776,
  -43.0804,
  -43.0832,
  -43.0864,
  -43.089,
  -43.0907,
  -43.0912,
  -43.0911,
  -43.0905,
  -43.0897,
  -43.0888,
  -43.0879,
  -43.0873,
  -43.0868,
  -43.0854,
  -43.0828,
  -43.0783,
  -43.0736,
  -43.0679,
  -43.0611,
  -43.0537,
  -43.0461,
  -43.0387,
  -43.0321,
  -43.0267,
  -43.0226,
  -43.02,
  -43.0183,
  -43.017,
  -43.0153,
  -43.0122,
  -43.0077,
  -43.0018,
  -42.9945,
  -42.9865,
  -42.9778,
  -42.9682,
  -42.957,
  -42.9433,
  -42.9256,
  -42.902,
  -42.8721,
  -42.8356,
  -42.7925,
  -42.7424,
  -42.6851,
  -42.6199,
  -42.5463,
  -42.4634,
  -42.3705,
  -42.2669,
  -42.1517,
  -42.0248,
  -41.8877,
  -41.7435,
  -41.5966,
  -41.4515,
  -41.3121,
  -41.1814,
  -41.0615,
  -40.9535,
  -40.8556,
  -40.7681,
  -39.8252,
  -39.8783,
  -39.9328,
  -39.987,
  -40.0398,
  -40.0905,
  -40.1392,
  -40.1861,
  -40.232,
  -40.2777,
  -40.3232,
  -40.3694,
  -40.416,
  -40.463,
  -40.5097,
  -40.5541,
  -40.5976,
  -40.6386,
  -40.6772,
  -40.7139,
  -40.7488,
  -40.7829,
  -40.8165,
  -40.8496,
  -40.882,
  -40.9132,
  -40.9428,
  -40.9707,
  -40.9967,
  -41.0215,
  -41.044,
  -41.0654,
  -41.0852,
  -41.1034,
  -41.1197,
  -41.1349,
  -41.1489,
  -41.1628,
  -41.1768,
  -41.1909,
  -41.2051,
  -41.2194,
  -41.2335,
  -41.2477,
  -41.2621,
  -41.2766,
  -41.2899,
  -41.3038,
  -41.3171,
  -41.3302,
  -41.343,
  -41.3557,
  -41.3693,
  -41.3835,
  -41.3979,
  -41.4122,
  -41.425,
  -41.4361,
  -41.4459,
  -41.455,
  -41.4643,
  -41.4747,
  -41.4848,
  -41.4964,
  -41.5079,
  -41.5189,
  -41.5295,
  -41.54,
  -41.5505,
  -41.5612,
  -41.5724,
  -41.5844,
  -41.5978,
  -41.6125,
  -41.6285,
  -41.6459,
  -41.6641,
  -41.6826,
  -41.7013,
  -41.7187,
  -41.737,
  -41.7553,
  -41.7736,
  -41.7918,
  -41.8097,
  -41.8272,
  -41.8444,
  -41.8617,
  -41.8799,
  -41.8992,
  -41.9198,
  -41.9412,
  -41.9625,
  -41.9836,
  -42.005,
  -42.0259,
  -42.0468,
  -42.0667,
  -42.0881,
  -42.11,
  -42.1316,
  -42.1537,
  -42.1763,
  -42.1992,
  -42.2224,
  -42.2453,
  -42.2671,
  -42.2866,
  -42.3044,
  -42.3197,
  -42.333,
  -42.3451,
  -42.3564,
  -42.3679,
  -42.3801,
  -42.3929,
  -42.405,
  -42.4172,
  -42.4281,
  -42.4371,
  -42.4443,
  -42.4505,
  -42.4555,
  -42.4595,
  -42.4629,
  -42.4657,
  -42.4684,
  -42.4716,
  -42.4756,
  -42.4809,
  -42.4876,
  -42.4955,
  -42.5047,
  -42.5149,
  -42.5263,
  -42.539,
  -42.5529,
  -42.5671,
  -42.5832,
  -42.5995,
  -42.6159,
  -42.6318,
  -42.6477,
  -42.6635,
  -42.6795,
  -42.6954,
  -42.7112,
  -42.7268,
  -42.7423,
  -42.7573,
  -42.7717,
  -42.7852,
  -42.7983,
  -42.811,
  -42.8237,
  -42.8367,
  -42.8497,
  -42.8622,
  -42.8737,
  -42.8834,
  -42.8936,
  -42.9038,
  -42.915,
  -42.9271,
  -42.941,
  -42.9567,
  -42.9743,
  -42.9933,
  -43.0127,
  -43.0319,
  -43.0501,
  -43.0667,
  -43.0815,
  -43.0941,
  -43.1049,
  -43.1145,
  -43.1233,
  -43.1315,
  -43.1392,
  -43.1467,
  -43.1542,
  -43.1623,
  -43.1709,
  -43.1789,
  -43.1877,
  -43.1963,
  -43.2038,
  -43.2103,
  -43.2159,
  -43.2201,
  -43.2225,
  -43.2234,
  -43.2228,
  -43.2212,
  -43.218,
  -43.2136,
  -43.2077,
  -43.2007,
  -43.1925,
  -43.1839,
  -43.175,
  -43.1664,
  -43.1587,
  -43.1517,
  -43.1456,
  -43.1399,
  -43.1343,
  -43.128,
  -43.1212,
  -43.1139,
  -43.1054,
  -43.0981,
  -43.0905,
  -43.0827,
  -43.0742,
  -43.0658,
  -43.0567,
  -43.0477,
  -43.039,
  -43.0301,
  -43.0215,
  -43.0136,
  -43.0067,
  -43.0013,
  -42.9979,
  -42.9966,
  -42.997,
  -42.9992,
  -43.0031,
  -43.0079,
  -43.0129,
  -43.0174,
  -43.0218,
  -43.0254,
  -43.0285,
  -43.0312,
  -43.0338,
  -43.0364,
  -43.0389,
  -43.0417,
  -43.0449,
  -43.0481,
  -43.0499,
  -43.0522,
  -43.0538,
  -43.0546,
  -43.0548,
  -43.0547,
  -43.0547,
  -43.0537,
  -43.0531,
  -43.0526,
  -43.0509,
  -43.0484,
  -43.045,
  -43.0403,
  -43.0343,
  -43.0272,
  -43.0194,
  -43.0111,
  -43.0028,
  -42.9952,
  -42.9888,
  -42.9842,
  -42.981,
  -42.9791,
  -42.9779,
  -42.9765,
  -42.9743,
  -42.9707,
  -42.9653,
  -42.9586,
  -42.9506,
  -42.9418,
  -42.9315,
  -42.9196,
  -42.9049,
  -42.8861,
  -42.8621,
  -42.832,
  -42.7956,
  -42.7528,
  -42.7024,
  -42.646,
  -42.5823,
  -42.511,
  -42.4312,
  -42.3421,
  -42.2425,
  -42.1315,
  -42.0091,
  -41.8761,
  -41.7356,
  -41.5917,
  -41.4487,
  -41.3103,
  -41.1799,
  -41.0601,
  -40.9518,
  -40.8546,
  -40.7673,
  -39.6819,
  -39.7352,
  -39.7891,
  -39.8429,
  -39.8957,
  -39.9466,
  -39.9956,
  -40.043,
  -40.0893,
  -40.135,
  -40.1795,
  -40.2253,
  -40.2716,
  -40.318,
  -40.364,
  -40.4087,
  -40.4514,
  -40.4918,
  -40.5299,
  -40.5663,
  -40.6013,
  -40.6354,
  -40.6693,
  -40.7029,
  -40.7356,
  -40.7661,
  -40.796,
  -40.8241,
  -40.8503,
  -40.875,
  -40.8985,
  -40.9203,
  -40.9402,
  -40.9585,
  -40.9755,
  -40.9913,
  -41.0066,
  -41.0215,
  -41.0366,
  -41.0521,
  -41.0664,
  -41.0816,
  -41.0964,
  -41.1115,
  -41.1267,
  -41.142,
  -41.1571,
  -41.172,
  -41.1866,
  -41.2003,
  -41.2138,
  -41.2274,
  -41.2419,
  -41.2572,
  -41.2729,
  -41.2881,
  -41.3011,
  -41.3133,
  -41.3241,
  -41.3343,
  -41.3445,
  -41.3556,
  -41.3673,
  -41.3793,
  -41.391,
  -41.4025,
  -41.4137,
  -41.4246,
  -41.4357,
  -41.4473,
  -41.4593,
  -41.472,
  -41.4859,
  -41.5002,
  -41.517,
  -41.5353,
  -41.5544,
  -41.5737,
  -41.593,
  -41.6124,
  -41.6318,
  -41.6513,
  -41.6711,
  -41.6909,
  -41.7101,
  -41.7283,
  -41.746,
  -41.7638,
  -41.7825,
  -41.8021,
  -41.8233,
  -41.8445,
  -41.8666,
  -41.8883,
  -41.9097,
  -41.9309,
  -41.9521,
  -41.9731,
  -41.9945,
  -42.016,
  -42.0379,
  -42.0601,
  -42.0825,
  -42.1052,
  -42.1281,
  -42.151,
  -42.173,
  -42.1933,
  -42.2112,
  -42.2264,
  -42.2387,
  -42.2503,
  -42.2614,
  -42.2723,
  -42.2834,
  -42.2948,
  -42.3063,
  -42.3172,
  -42.3269,
  -42.3347,
  -42.3411,
  -42.3463,
  -42.3504,
  -42.3536,
  -42.3564,
  -42.3586,
  -42.3604,
  -42.3626,
  -42.3659,
  -42.3706,
  -42.3761,
  -42.3841,
  -42.3933,
  -42.4039,
  -42.4156,
  -42.4284,
  -42.4424,
  -42.4571,
  -42.4726,
  -42.4886,
  -42.5043,
  -42.5198,
  -42.5354,
  -42.5509,
  -42.5666,
  -42.5821,
  -42.5978,
  -42.6135,
  -42.6293,
  -42.6445,
  -42.6588,
  -42.6712,
  -42.6837,
  -42.6962,
  -42.7089,
  -42.7223,
  -42.7358,
  -42.7488,
  -42.7606,
  -42.7717,
  -42.7821,
  -42.7924,
  -42.8033,
  -42.8154,
  -42.8289,
  -42.8446,
  -42.8619,
  -42.881,
  -42.9012,
  -42.9212,
  -42.9405,
  -42.9586,
  -42.9748,
  -42.989,
  -43.0015,
  -43.0117,
  -43.0217,
  -43.0313,
  -43.0405,
  -43.0494,
  -43.0588,
  -43.0683,
  -43.0784,
  -43.0889,
  -43.099,
  -43.1088,
  -43.1176,
  -43.1254,
  -43.1324,
  -43.1383,
  -43.1426,
  -43.1454,
  -43.1465,
  -43.1463,
  -43.1447,
  -43.1414,
  -43.1367,
  -43.1307,
  -43.1238,
  -43.1163,
  -43.1088,
  -43.1005,
  -43.0936,
  -43.0874,
  -43.0821,
  -43.0766,
  -43.0712,
  -43.0651,
  -43.0585,
  -43.0515,
  -43.0446,
  -43.0376,
  -43.0304,
  -43.0231,
  -43.0151,
  -43.007,
  -42.998,
  -42.9891,
  -42.9801,
  -42.9716,
  -42.9637,
  -42.9566,
  -42.9506,
  -42.9465,
  -42.9442,
  -42.9438,
  -42.9453,
  -42.9488,
  -42.9535,
  -42.9591,
  -42.9651,
  -42.9698,
  -42.9752,
  -42.98,
  -42.9841,
  -42.9877,
  -42.9908,
  -42.9937,
  -42.9966,
  -42.9995,
  -43.0027,
  -43.0058,
  -43.0089,
  -43.0118,
  -43.0139,
  -43.0157,
  -43.0169,
  -43.0174,
  -43.0173,
  -43.0172,
  -43.0164,
  -43.0157,
  -43.0139,
  -43.0115,
  -43.0078,
  -43.0028,
  -42.9969,
  -42.9899,
  -42.982,
  -42.9735,
  -42.965,
  -42.9568,
  -42.9497,
  -42.9445,
  -42.9409,
  -42.9388,
  -42.9373,
  -42.936,
  -42.9333,
  -42.9303,
  -42.9258,
  -42.9197,
  -42.9119,
  -42.9027,
  -42.8921,
  -42.8794,
  -42.8639,
  -42.8446,
  -42.8202,
  -42.79,
  -42.7535,
  -42.7108,
  -42.6618,
  -42.6062,
  -42.5441,
  -42.4749,
  -42.3979,
  -42.3122,
  -42.2165,
  -42.1097,
  -41.9916,
  -41.8631,
  -41.7268,
  -41.5867,
  -41.4467,
  -41.3108,
  -41.1819,
  -41.0631,
  -40.9554,
  -40.8587,
  -40.7717,
  -39.5372,
  -39.5894,
  -39.6423,
  -39.6955,
  -39.7477,
  -39.7976,
  -39.8468,
  -39.8945,
  -39.9411,
  -39.9869,
  -40.0324,
  -40.078,
  -40.1238,
  -40.1695,
  -40.2147,
  -40.2587,
  -40.3007,
  -40.3407,
  -40.3787,
  -40.415,
  -40.4491,
  -40.4836,
  -40.5178,
  -40.5518,
  -40.585,
  -40.617,
  -40.6472,
  -40.6755,
  -40.7019,
  -40.7269,
  -40.7504,
  -40.772,
  -40.7921,
  -40.8105,
  -40.8277,
  -40.8431,
  -40.859,
  -40.875,
  -40.8912,
  -40.9076,
  -40.9239,
  -40.9398,
  -40.9558,
  -40.9715,
  -40.9879,
  -41.0042,
  -41.0203,
  -41.0364,
  -41.0516,
  -41.0661,
  -41.0806,
  -41.0941,
  -41.1096,
  -41.1259,
  -41.1426,
  -41.159,
  -41.174,
  -41.1874,
  -41.1993,
  -41.2106,
  -41.2223,
  -41.2341,
  -41.2463,
  -41.2588,
  -41.2712,
  -41.2832,
  -41.2951,
  -41.3058,
  -41.3175,
  -41.3294,
  -41.3423,
  -41.3558,
  -41.3706,
  -41.3868,
  -41.4046,
  -41.4237,
  -41.4434,
  -41.4634,
  -41.4836,
  -41.5038,
  -41.5243,
  -41.5454,
  -41.5667,
  -41.5877,
  -41.6079,
  -41.6261,
  -41.6445,
  -41.6627,
  -41.682,
  -41.7024,
  -41.7241,
  -41.7467,
  -41.7695,
  -41.7918,
  -41.8135,
  -41.8347,
  -41.8558,
  -41.877,
  -41.8984,
  -41.9197,
  -41.9416,
  -41.9637,
  -41.9861,
  -42.0079,
  -42.0307,
  -42.0534,
  -42.0756,
  -42.0962,
  -42.1148,
  -42.1303,
  -42.1435,
  -42.1551,
  -42.166,
  -42.1764,
  -42.1866,
  -42.1967,
  -42.2065,
  -42.2159,
  -42.2243,
  -42.2313,
  -42.2368,
  -42.2411,
  -42.2445,
  -42.2462,
  -42.2483,
  -42.2499,
  -42.2515,
  -42.2532,
  -42.2561,
  -42.2606,
  -42.2671,
  -42.2753,
  -42.2848,
  -42.2955,
  -42.3075,
  -42.3205,
  -42.3343,
  -42.3486,
  -42.3634,
  -42.3782,
  -42.3931,
  -42.408,
  -42.4231,
  -42.4384,
  -42.4528,
  -42.468,
  -42.4836,
  -42.4994,
  -42.5152,
  -42.5303,
  -42.5444,
  -42.5573,
  -42.5695,
  -42.5816,
  -42.5944,
  -42.6079,
  -42.6215,
  -42.6348,
  -42.647,
  -42.6582,
  -42.6686,
  -42.679,
  -42.6898,
  -42.7015,
  -42.7147,
  -42.7299,
  -42.7474,
  -42.7657,
  -42.7862,
  -42.8071,
  -42.8274,
  -42.8469,
  -42.8647,
  -42.8806,
  -42.8946,
  -42.9073,
  -42.919,
  -42.93,
  -42.9406,
  -42.9514,
  -42.9622,
  -42.9737,
  -42.9856,
  -42.9975,
  -43.0091,
  -43.0199,
  -43.0299,
  -43.039,
  -43.0473,
  -43.0547,
  -43.0606,
  -43.0651,
  -43.0672,
  -43.0687,
  -43.0684,
  -43.0665,
  -43.063,
  -43.0579,
  -43.0521,
  -43.0458,
  -43.0396,
  -43.0336,
  -43.028,
  -43.0231,
  -43.0182,
  -43.0134,
  -43.0079,
  -43.0022,
  -42.996,
  -42.9896,
  -42.9829,
  -42.9761,
  -42.9691,
  -42.9618,
  -42.9543,
  -42.9462,
  -42.9375,
  -42.9284,
  -42.9196,
  -42.9117,
  -42.9036,
  -42.8975,
  -42.8929,
  -42.8897,
  -42.8881,
  -42.8887,
  -42.8912,
  -42.8953,
  -42.9009,
  -42.9074,
  -42.9144,
  -42.9212,
  -42.9278,
  -42.9337,
  -42.9387,
  -42.9429,
  -42.9462,
  -42.9492,
  -42.9524,
  -42.9554,
  -42.9585,
  -42.9618,
  -42.9654,
  -42.9687,
  -42.9718,
  -42.9743,
  -42.9762,
  -42.9771,
  -42.9779,
  -42.9776,
  -42.9775,
  -42.9763,
  -42.9742,
  -42.9713,
  -42.9664,
  -42.9614,
  -42.9556,
  -42.9488,
  -42.9411,
  -42.9326,
  -42.9241,
  -42.916,
  -42.9088,
  -42.9032,
  -42.8993,
  -42.8965,
  -42.8948,
  -42.8934,
  -42.8918,
  -42.8895,
  -42.8856,
  -42.8799,
  -42.8724,
  -42.8631,
  -42.8523,
  -42.839,
  -42.823,
  -42.8032,
  -42.7785,
  -42.7482,
  -42.7119,
  -42.6691,
  -42.6202,
  -42.5653,
  -42.5043,
  -42.4368,
  -42.3622,
  -42.2794,
  -42.187,
  -42.0842,
  -41.9704,
  -41.8464,
  -41.7147,
  -41.5789,
  -41.4428,
  -41.3104,
  -41.1847,
  -41.068,
  -40.9619,
  -40.8651,
  -40.7786,
  -39.3911,
  -39.4411,
  -39.4927,
  -39.5447,
  -39.596,
  -39.6463,
  -39.6953,
  -39.7431,
  -39.7898,
  -39.8358,
  -39.8813,
  -39.9266,
  -39.972,
  -40.0172,
  -40.0617,
  -40.1039,
  -40.1455,
  -40.1852,
  -40.2232,
  -40.2596,
  -40.2952,
  -40.3302,
  -40.365,
  -40.3995,
  -40.4332,
  -40.4656,
  -40.4962,
  -40.5249,
  -40.5517,
  -40.5766,
  -40.5988,
  -40.6202,
  -40.6401,
  -40.6585,
  -40.6757,
  -40.6923,
  -40.7089,
  -40.7257,
  -40.7427,
  -40.76,
  -40.7773,
  -40.7946,
  -40.8115,
  -40.8286,
  -40.8459,
  -40.8633,
  -40.8796,
  -40.8965,
  -40.9129,
  -40.9287,
  -40.9443,
  -40.96,
  -40.9763,
  -40.9932,
  -41.0107,
  -41.0279,
  -41.0439,
  -41.0584,
  -41.0716,
  -41.0843,
  -41.0968,
  -41.1096,
  -41.1216,
  -41.1346,
  -41.1478,
  -41.1608,
  -41.1735,
  -41.1859,
  -41.1983,
  -41.2111,
  -41.2245,
  -41.2392,
  -41.2552,
  -41.2728,
  -41.2917,
  -41.3114,
  -41.3315,
  -41.352,
  -41.3729,
  -41.393,
  -41.4149,
  -41.4373,
  -41.4597,
  -41.4817,
  -41.5027,
  -41.5228,
  -41.5421,
  -41.5611,
  -41.5807,
  -41.6017,
  -41.6241,
  -41.6473,
  -41.6709,
  -41.6935,
  -41.7155,
  -41.7367,
  -41.7577,
  -41.7778,
  -41.7992,
  -41.8208,
  -41.8426,
  -41.8646,
  -41.8872,
  -41.9098,
  -41.9323,
  -41.9549,
  -41.9769,
  -41.998,
  -42.0172,
  -42.0335,
  -42.047,
  -42.0584,
  -42.0691,
  -42.079,
  -42.0885,
  -42.0975,
  -42.105,
  -42.1131,
  -42.1202,
  -42.1263,
  -42.131,
  -42.1346,
  -42.1373,
  -42.1393,
  -42.1409,
  -42.1423,
  -42.1438,
  -42.1459,
  -42.1488,
  -42.1534,
  -42.1599,
  -42.1681,
  -42.1778,
  -42.1888,
  -42.2009,
  -42.2139,
  -42.2275,
  -42.2404,
  -42.2544,
  -42.2682,
  -42.282,
  -42.2963,
  -42.3109,
  -42.3258,
  -42.3408,
  -42.3562,
  -42.3716,
  -42.3873,
  -42.4027,
  -42.4175,
  -42.431,
  -42.4433,
  -42.455,
  -42.4668,
  -42.4795,
  -42.4928,
  -42.5064,
  -42.5197,
  -42.5321,
  -42.5423,
  -42.5528,
  -42.5632,
  -42.5738,
  -42.5853,
  -42.5984,
  -42.6134,
  -42.6308,
  -42.6502,
  -42.6713,
  -42.693,
  -42.7146,
  -42.7352,
  -42.7543,
  -42.7717,
  -42.7873,
  -42.8015,
  -42.8146,
  -42.8271,
  -42.8394,
  -42.8518,
  -42.8645,
  -42.878,
  -42.8915,
  -42.9041,
  -42.9171,
  -42.9293,
  -42.9405,
  -42.9507,
  -42.9601,
  -42.9686,
  -42.9761,
  -42.9823,
  -42.9872,
  -42.9902,
  -42.9915,
  -42.9907,
  -42.9881,
  -42.9843,
  -42.9795,
  -42.9746,
  -42.9697,
  -42.9652,
  -42.961,
  -42.9571,
  -42.9533,
  -42.9488,
  -42.944,
  -42.9387,
  -42.933,
  -42.9268,
  -42.9191,
  -42.9125,
  -42.9056,
  -42.8986,
  -42.891,
  -42.883,
  -42.8743,
  -42.8655,
  -42.8575,
  -42.8501,
  -42.8439,
  -42.8389,
  -42.8353,
  -42.833,
  -42.8323,
  -42.8339,
  -42.8371,
  -42.8419,
  -42.8481,
  -42.8554,
  -42.8631,
  -42.871,
  -42.8785,
  -42.8852,
  -42.8908,
  -42.8952,
  -42.8986,
  -42.9017,
  -42.905,
  -42.9082,
  -42.9118,
  -42.9155,
  -42.9184,
  -42.9225,
  -42.9263,
  -42.9295,
  -42.9319,
  -42.9336,
  -42.9347,
  -42.9354,
  -42.9353,
  -42.9342,
  -42.9314,
  -42.9282,
  -42.9241,
  -42.9191,
  -42.9134,
  -42.9069,
  -42.8995,
  -42.8913,
  -42.8829,
  -42.8748,
  -42.868,
  -42.8621,
  -42.8578,
  -42.8547,
  -42.8524,
  -42.851,
  -42.8495,
  -42.8475,
  -42.8441,
  -42.8389,
  -42.8319,
  -42.8228,
  -42.8115,
  -42.7979,
  -42.7813,
  -42.7609,
  -42.7361,
  -42.7057,
  -42.6694,
  -42.6269,
  -42.5773,
  -42.523,
  -42.4626,
  -42.3964,
  -42.3235,
  -42.2427,
  -42.153,
  -42.0534,
  -41.9436,
  -41.8239,
  -41.6969,
  -41.5659,
  -41.4347,
  -41.3068,
  -41.1853,
  -41.0719,
  -40.9683,
  -40.8741,
  -40.7885,
  -39.2422,
  -39.2923,
  -39.3429,
  -39.3936,
  -39.444,
  -39.4934,
  -39.5417,
  -39.5889,
  -39.6353,
  -39.6812,
  -39.7256,
  -39.7708,
  -39.8159,
  -39.8608,
  -39.9049,
  -39.9477,
  -39.9888,
  -40.0283,
  -40.0663,
  -40.103,
  -40.139,
  -40.1746,
  -40.2099,
  -40.245,
  -40.2793,
  -40.3113,
  -40.3424,
  -40.3714,
  -40.3981,
  -40.4228,
  -40.4455,
  -40.4665,
  -40.4859,
  -40.5043,
  -40.5217,
  -40.5386,
  -40.5558,
  -40.5734,
  -40.5913,
  -40.6097,
  -40.6273,
  -40.6456,
  -40.664,
  -40.6823,
  -40.7008,
  -40.7194,
  -40.7377,
  -40.7559,
  -40.7736,
  -40.7908,
  -40.8076,
  -40.8246,
  -40.8419,
  -40.8595,
  -40.8774,
  -40.8951,
  -40.9109,
  -40.9262,
  -40.9406,
  -40.9542,
  -40.9678,
  -40.9816,
  -40.9955,
  -41.0094,
  -41.0234,
  -41.0375,
  -41.0514,
  -41.0649,
  -41.0784,
  -41.0921,
  -41.1067,
  -41.1225,
  -41.1399,
  -41.1575,
  -41.1772,
  -41.1978,
  -41.2184,
  -41.2393,
  -41.2606,
  -41.2827,
  -41.3056,
  -41.329,
  -41.3526,
  -41.3755,
  -41.3972,
  -41.4179,
  -41.4379,
  -41.4581,
  -41.4787,
  -41.5001,
  -41.5231,
  -41.5459,
  -41.5699,
  -41.593,
  -41.6152,
  -41.6366,
  -41.6576,
  -41.6785,
  -41.6998,
  -41.7214,
  -41.7433,
  -41.7655,
  -41.7879,
  -41.8106,
  -41.8329,
  -41.855,
  -41.8768,
  -41.8978,
  -41.9173,
  -41.9342,
  -41.9476,
  -41.9594,
  -41.9698,
  -41.9792,
  -41.9881,
  -41.9964,
  -42.0038,
  -42.0106,
  -42.0167,
  -42.022,
  -42.0261,
  -42.0289,
  -42.0309,
  -42.0325,
  -42.0338,
  -42.0352,
  -42.0367,
  -42.0392,
  -42.0425,
  -42.0474,
  -42.0532,
  -42.0614,
  -42.0713,
  -42.0824,
  -42.0947,
  -42.1075,
  -42.1208,
  -42.134,
  -42.1471,
  -42.16,
  -42.1731,
  -42.1867,
  -42.2008,
  -42.2155,
  -42.2305,
  -42.2456,
  -42.2608,
  -42.2762,
  -42.2911,
  -42.3051,
  -42.3179,
  -42.3285,
  -42.3398,
  -42.3512,
  -42.3634,
  -42.3765,
  -42.3898,
  -42.4029,
  -42.4154,
  -42.4268,
  -42.4373,
  -42.4476,
  -42.4582,
  -42.4699,
  -42.4829,
  -42.498,
  -42.5154,
  -42.5354,
  -42.557,
  -42.5795,
  -42.6021,
  -42.6241,
  -42.6445,
  -42.6632,
  -42.6799,
  -42.6943,
  -42.7087,
  -42.7227,
  -42.7364,
  -42.7503,
  -42.7647,
  -42.78,
  -42.7954,
  -42.8106,
  -42.8252,
  -42.8387,
  -42.8511,
  -42.8625,
  -42.8727,
  -42.8823,
  -42.8912,
  -42.899,
  -42.9055,
  -42.9101,
  -42.9126,
  -42.913,
  -42.9115,
  -42.9087,
  -42.9053,
  -42.9017,
  -42.8981,
  -42.8942,
  -42.8914,
  -42.8887,
  -42.8856,
  -42.8822,
  -42.878,
  -42.8735,
  -42.8683,
  -42.8622,
  -42.8558,
  -42.8492,
  -42.8422,
  -42.835,
  -42.8273,
  -42.8191,
  -42.8109,
  -42.8028,
  -42.7952,
  -42.7888,
  -42.7835,
  -42.7796,
  -42.7769,
  -42.7753,
  -42.7758,
  -42.7778,
  -42.7818,
  -42.7874,
  -42.7944,
  -42.8021,
  -42.8106,
  -42.818,
  -42.8259,
  -42.8331,
  -42.8388,
  -42.8432,
  -42.8467,
  -42.85,
  -42.8534,
  -42.8573,
  -42.8617,
  -42.8666,
  -42.8713,
  -42.8759,
  -42.88,
  -42.8834,
  -42.8863,
  -42.8888,
  -42.8905,
  -42.8914,
  -42.8915,
  -42.8902,
  -42.8879,
  -42.8847,
  -42.8806,
  -42.8757,
  -42.8701,
  -42.8638,
  -42.8569,
  -42.8491,
  -42.841,
  -42.8334,
  -42.8263,
  -42.8203,
  -42.8154,
  -42.8117,
  -42.8091,
  -42.8073,
  -42.8048,
  -42.8031,
  -42.8003,
  -42.7958,
  -42.7892,
  -42.7804,
  -42.7691,
  -42.7552,
  -42.7381,
  -42.7172,
  -42.6918,
  -42.6613,
  -42.6252,
  -42.5831,
  -42.5353,
  -42.4815,
  -42.4219,
  -42.3565,
  -42.2846,
  -42.2053,
  -42.1176,
  -42.0206,
  -41.914,
  -41.7983,
  -41.6758,
  -41.5498,
  -41.4237,
  -41.3008,
  -41.1838,
  -41.0748,
  -40.9744,
  -40.8825,
  -40.7979,
  -39.0935,
  -39.1429,
  -39.1927,
  -39.2423,
  -39.2914,
  -39.3386,
  -39.3858,
  -39.4321,
  -39.4779,
  -39.5231,
  -39.5683,
  -39.6133,
  -39.6582,
  -39.7029,
  -39.7468,
  -39.7894,
  -39.8304,
  -39.8698,
  -39.9077,
  -39.9447,
  -39.98,
  -40.016,
  -40.0519,
  -40.0875,
  -40.1223,
  -40.1557,
  -40.1872,
  -40.2162,
  -40.2429,
  -40.2671,
  -40.2891,
  -40.3097,
  -40.3288,
  -40.3471,
  -40.3647,
  -40.3813,
  -40.3992,
  -40.4177,
  -40.437,
  -40.4567,
  -40.4766,
  -40.4963,
  -40.5159,
  -40.5354,
  -40.5549,
  -40.5746,
  -40.5942,
  -40.6136,
  -40.6329,
  -40.6516,
  -40.6701,
  -40.6873,
  -40.7054,
  -40.7237,
  -40.7421,
  -40.7601,
  -40.7775,
  -40.7937,
  -40.8089,
  -40.8237,
  -40.8385,
  -40.8532,
  -40.8679,
  -40.8827,
  -40.8977,
  -40.9129,
  -40.928,
  -40.9419,
  -40.9566,
  -40.9718,
  -40.9875,
  -41.0047,
  -41.0229,
  -41.0426,
  -41.0631,
  -41.0843,
  -41.1057,
  -41.1273,
  -41.1492,
  -41.1722,
  -41.196,
  -41.2204,
  -41.2447,
  -41.2684,
  -41.2909,
  -41.3112,
  -41.332,
  -41.3529,
  -41.3746,
  -41.3969,
  -41.4203,
  -41.4445,
  -41.469,
  -41.4924,
  -41.5148,
  -41.5365,
  -41.5577,
  -41.5788,
  -41.6001,
  -41.6217,
  -41.6438,
  -41.6663,
  -41.6886,
  -41.71,
  -41.7322,
  -41.7537,
  -41.7751,
  -41.7958,
  -41.8153,
  -41.8326,
  -41.8475,
  -41.8601,
  -41.8707,
  -41.8798,
  -41.8878,
  -41.895,
  -41.9015,
  -41.9074,
  -41.9128,
  -41.9174,
  -41.9207,
  -41.923,
  -41.9244,
  -41.9246,
  -41.9257,
  -41.9271,
  -41.929,
  -41.9317,
  -41.9356,
  -41.9411,
  -41.9481,
  -41.9566,
  -41.9666,
  -41.9775,
  -41.9897,
  -42.0023,
  -42.0152,
  -42.0278,
  -42.0402,
  -42.0524,
  -42.0649,
  -42.0779,
  -42.0916,
  -42.106,
  -42.1199,
  -42.135,
  -42.1501,
  -42.1649,
  -42.1792,
  -42.1925,
  -42.2044,
  -42.2154,
  -42.2261,
  -42.2371,
  -42.2489,
  -42.2614,
  -42.2745,
  -42.2875,
  -42.2998,
  -42.3112,
  -42.322,
  -42.3325,
  -42.3433,
  -42.355,
  -42.3684,
  -42.3838,
  -42.4017,
  -42.4211,
  -42.4433,
  -42.4668,
  -42.4904,
  -42.5135,
  -42.535,
  -42.5546,
  -42.5723,
  -42.5888,
  -42.6041,
  -42.619,
  -42.6339,
  -42.6493,
  -42.6652,
  -42.6819,
  -42.699,
  -42.716,
  -42.7321,
  -42.7471,
  -42.7606,
  -42.7729,
  -42.7842,
  -42.7948,
  -42.8049,
  -42.8143,
  -42.821,
  -42.827,
  -42.8307,
  -42.8321,
  -42.8321,
  -42.8306,
  -42.8284,
  -42.8261,
  -42.8242,
  -42.8226,
  -42.821,
  -42.8194,
  -42.8177,
  -42.815,
  -42.812,
  -42.808,
  -42.8035,
  -42.7979,
  -42.7917,
  -42.7851,
  -42.7779,
  -42.7703,
  -42.7626,
  -42.7545,
  -42.7466,
  -42.7391,
  -42.7324,
  -42.7267,
  -42.7212,
  -42.7178,
  -42.7159,
  -42.7153,
  -42.7167,
  -42.7196,
  -42.7246,
  -42.7308,
  -42.7384,
  -42.7465,
  -42.7554,
  -42.7641,
  -42.7721,
  -42.7791,
  -42.7847,
  -42.7891,
  -42.7929,
  -42.7967,
  -42.8006,
  -42.8055,
  -42.8108,
  -42.8165,
  -42.8219,
  -42.8268,
  -42.8313,
  -42.8353,
  -42.8388,
  -42.8415,
  -42.8436,
  -42.8449,
  -42.8452,
  -42.8445,
  -42.8425,
  -42.8397,
  -42.8349,
  -42.8303,
  -42.8251,
  -42.8191,
  -42.8124,
  -42.8051,
  -42.7975,
  -42.7898,
  -42.7829,
  -42.7765,
  -42.771,
  -42.7665,
  -42.7633,
  -42.761,
  -42.7595,
  -42.7579,
  -42.7556,
  -42.7516,
  -42.7456,
  -42.7373,
  -42.7262,
  -42.7123,
  -42.695,
  -42.6736,
  -42.6479,
  -42.6175,
  -42.5816,
  -42.5403,
  -42.4932,
  -42.4404,
  -42.3817,
  -42.317,
  -42.2456,
  -42.1672,
  -42.0808,
  -41.9859,
  -41.882,
  -41.7699,
  -41.6517,
  -41.5305,
  -41.4096,
  -41.2915,
  -41.1792,
  -41.0741,
  -40.9772,
  -40.887,
  -40.8047,
  -38.9442,
  -38.9924,
  -39.0413,
  -39.0898,
  -39.1376,
  -39.1844,
  -39.2301,
  -39.2751,
  -39.3198,
  -39.3646,
  -39.4093,
  -39.4542,
  -39.499,
  -39.5436,
  -39.5874,
  -39.6289,
  -39.6699,
  -39.7093,
  -39.7472,
  -39.7841,
  -39.8206,
  -39.8569,
  -39.8932,
  -39.9291,
  -39.9643,
  -39.998,
  -40.0296,
  -40.0587,
  -40.0848,
  -40.1083,
  -40.1286,
  -40.1488,
  -40.1678,
  -40.1862,
  -40.2043,
  -40.2225,
  -40.2414,
  -40.2614,
  -40.282,
  -40.3032,
  -40.3246,
  -40.3459,
  -40.3668,
  -40.3874,
  -40.408,
  -40.4287,
  -40.4485,
  -40.4692,
  -40.4901,
  -40.5108,
  -40.5307,
  -40.5502,
  -40.5692,
  -40.5882,
  -40.6069,
  -40.6253,
  -40.6432,
  -40.6601,
  -40.6762,
  -40.6921,
  -40.7079,
  -40.7236,
  -40.7382,
  -40.7539,
  -40.77,
  -40.7861,
  -40.8025,
  -40.8188,
  -40.8354,
  -40.8521,
  -40.8695,
  -40.8875,
  -40.9067,
  -40.9272,
  -40.9484,
  -40.9699,
  -40.9919,
  -41.0144,
  -41.0376,
  -41.0605,
  -41.0852,
  -41.1106,
  -41.1356,
  -41.1596,
  -41.1826,
  -41.2045,
  -41.226,
  -41.2475,
  -41.27,
  -41.2933,
  -41.3173,
  -41.3421,
  -41.3666,
  -41.3903,
  -41.4134,
  -41.4356,
  -41.4571,
  -41.4776,
  -41.4993,
  -41.5211,
  -41.5435,
  -41.5662,
  -41.5889,
  -41.6112,
  -41.6331,
  -41.6543,
  -41.6748,
  -41.6951,
  -41.7141,
  -41.7314,
  -41.7469,
  -41.7601,
  -41.7711,
  -41.7798,
  -41.7872,
  -41.7936,
  -41.7982,
  -41.8032,
  -41.8078,
  -41.8115,
  -41.8142,
  -41.8159,
  -41.8169,
  -41.8178,
  -41.8187,
  -41.82,
  -41.8222,
  -41.8254,
  -41.8297,
  -41.8356,
  -41.843,
  -41.8516,
  -41.8616,
  -41.8726,
  -41.8843,
  -41.8966,
  -41.9093,
  -41.9204,
  -41.9323,
  -41.9442,
  -41.9562,
  -41.9689,
  -41.9823,
  -41.9965,
  -42.0113,
  -42.0263,
  -42.0411,
  -42.0556,
  -42.0692,
  -42.0815,
  -42.0929,
  -42.1035,
  -42.1139,
  -42.1248,
  -42.1362,
  -42.1482,
  -42.1608,
  -42.1733,
  -42.1855,
  -42.1961,
  -42.2071,
  -42.2182,
  -42.2295,
  -42.2418,
  -42.2554,
  -42.2713,
  -42.2895,
  -42.3104,
  -42.3333,
  -42.3576,
  -42.382,
  -42.4059,
  -42.4282,
  -42.4485,
  -42.4668,
  -42.4839,
  -42.5001,
  -42.5158,
  -42.5315,
  -42.5479,
  -42.565,
  -42.5832,
  -42.6018,
  -42.6192,
  -42.6367,
  -42.6529,
  -42.6673,
  -42.6807,
  -42.693,
  -42.7047,
  -42.7161,
  -42.7267,
  -42.7355,
  -42.7428,
  -42.7473,
  -42.75,
  -42.7511,
  -42.751,
  -42.7503,
  -42.7497,
  -42.7493,
  -42.7492,
  -42.7491,
  -42.7487,
  -42.748,
  -42.7465,
  -42.7441,
  -42.7411,
  -42.7371,
  -42.7322,
  -42.7253,
  -42.7186,
  -42.7111,
  -42.7033,
  -42.6958,
  -42.6882,
  -42.681,
  -42.6741,
  -42.668,
  -42.6628,
  -42.6585,
  -42.6555,
  -42.6541,
  -42.6544,
  -42.6568,
  -42.661,
  -42.667,
  -42.6741,
  -42.6821,
  -42.6906,
  -42.6996,
  -42.7083,
  -42.7161,
  -42.7227,
  -42.7284,
  -42.7331,
  -42.737,
  -42.741,
  -42.7458,
  -42.7515,
  -42.7576,
  -42.7637,
  -42.7686,
  -42.774,
  -42.779,
  -42.7838,
  -42.7872,
  -42.7905,
  -42.7927,
  -42.7943,
  -42.7954,
  -42.7954,
  -42.7944,
  -42.7923,
  -42.789,
  -42.785,
  -42.7803,
  -42.7748,
  -42.7685,
  -42.7617,
  -42.7543,
  -42.7468,
  -42.7395,
  -42.7326,
  -42.7263,
  -42.7208,
  -42.717,
  -42.7144,
  -42.7127,
  -42.7112,
  -42.709,
  -42.7056,
  -42.7001,
  -42.6925,
  -42.6818,
  -42.6681,
  -42.6507,
  -42.6292,
  -42.6034,
  -42.573,
  -42.5377,
  -42.4972,
  -42.4503,
  -42.3985,
  -42.3409,
  -42.2769,
  -42.206,
  -42.1284,
  -42.043,
  -41.9499,
  -41.8486,
  -41.7399,
  -41.6258,
  -41.5088,
  -41.3922,
  -41.2784,
  -41.17,
  -41.0691,
  -40.9757,
  -40.8892,
  -40.8094,
  -38.7934,
  -38.8422,
  -38.8905,
  -38.9378,
  -38.9842,
  -39.0295,
  -39.0739,
  -39.1176,
  -39.1614,
  -39.2052,
  -39.2485,
  -39.2931,
  -39.3378,
  -39.3823,
  -39.4262,
  -39.4687,
  -39.5097,
  -39.549,
  -39.587,
  -39.6239,
  -39.6603,
  -39.6966,
  -39.7329,
  -39.7689,
  -39.804,
  -39.8367,
  -39.8683,
  -39.8969,
  -39.9225,
  -39.9455,
  -39.9667,
  -39.9867,
  -40.0057,
  -40.0245,
  -40.0432,
  -40.0625,
  -40.0826,
  -40.1039,
  -40.1263,
  -40.1491,
  -40.1711,
  -40.1937,
  -40.2157,
  -40.2375,
  -40.2589,
  -40.2804,
  -40.3023,
  -40.3247,
  -40.3472,
  -40.3696,
  -40.3912,
  -40.412,
  -40.4322,
  -40.4519,
  -40.4711,
  -40.49,
  -40.5073,
  -40.5247,
  -40.5418,
  -40.5588,
  -40.5758,
  -40.5924,
  -40.6089,
  -40.6255,
  -40.6426,
  -40.66,
  -40.6776,
  -40.6955,
  -40.7134,
  -40.7315,
  -40.75,
  -40.7693,
  -40.7893,
  -40.8093,
  -40.8311,
  -40.8533,
  -40.8762,
  -40.8997,
  -40.9241,
  -40.9493,
  -40.9749,
  -41.0009,
  -41.0265,
  -41.051,
  -41.0745,
  -41.0969,
  -41.1192,
  -41.1415,
  -41.1644,
  -41.1882,
  -41.2126,
  -41.2368,
  -41.262,
  -41.2865,
  -41.3103,
  -41.3331,
  -41.3553,
  -41.3773,
  -41.3993,
  -41.4215,
  -41.4444,
  -41.4674,
  -41.4904,
  -41.5129,
  -41.5348,
  -41.5557,
  -41.576,
  -41.5956,
  -41.614,
  -41.6311,
  -41.6454,
  -41.6588,
  -41.67,
  -41.679,
  -41.6858,
  -41.6915,
  -41.6962,
  -41.7002,
  -41.704,
  -41.7069,
  -41.7089,
  -41.71,
  -41.7106,
  -41.7113,
  -41.7121,
  -41.7136,
  -41.716,
  -41.7194,
  -41.7243,
  -41.7304,
  -41.737,
  -41.7456,
  -41.7554,
  -41.7663,
  -41.7779,
  -41.7898,
  -41.802,
  -41.8142,
  -41.826,
  -41.8376,
  -41.8493,
  -41.8618,
  -41.8748,
  -41.8889,
  -41.9036,
  -41.9183,
  -41.9329,
  -41.9468,
  -41.9598,
  -41.9719,
  -41.9828,
  -41.9921,
  -42.0025,
  -42.0132,
  -42.0243,
  -42.036,
  -42.0482,
  -42.0604,
  -42.0727,
  -42.0848,
  -42.0964,
  -42.1078,
  -42.1199,
  -42.1326,
  -42.1468,
  -42.1631,
  -42.1818,
  -42.2031,
  -42.2266,
  -42.2513,
  -42.2763,
  -42.3004,
  -42.3229,
  -42.3436,
  -42.3624,
  -42.3789,
  -42.3954,
  -42.412,
  -42.4283,
  -42.4457,
  -42.4639,
  -42.4829,
  -42.5026,
  -42.522,
  -42.5404,
  -42.5575,
  -42.5731,
  -42.5876,
  -42.6015,
  -42.6146,
  -42.6269,
  -42.6386,
  -42.6487,
  -42.6568,
  -42.6625,
  -42.6665,
  -42.6687,
  -42.6699,
  -42.6707,
  -42.6715,
  -42.6726,
  -42.673,
  -42.6743,
  -42.6752,
  -42.6756,
  -42.675,
  -42.6735,
  -42.6712,
  -42.6676,
  -42.6632,
  -42.6576,
  -42.651,
  -42.6437,
  -42.6363,
  -42.6291,
  -42.622,
  -42.6157,
  -42.6096,
  -42.6037,
  -42.5986,
  -42.5942,
  -42.5915,
  -42.5908,
  -42.5921,
  -42.5957,
  -42.601,
  -42.6081,
  -42.6161,
  -42.6245,
  -42.6334,
  -42.6424,
  -42.6496,
  -42.6571,
  -42.6638,
  -42.6695,
  -42.6744,
  -42.6788,
  -42.6834,
  -42.6887,
  -42.6948,
  -42.701,
  -42.7074,
  -42.7136,
  -42.7197,
  -42.7254,
  -42.7301,
  -42.7343,
  -42.738,
  -42.7409,
  -42.7429,
  -42.7443,
  -42.7454,
  -42.7453,
  -42.7439,
  -42.7418,
  -42.7387,
  -42.7346,
  -42.7297,
  -42.7237,
  -42.7172,
  -42.7103,
  -42.7027,
  -42.6949,
  -42.6873,
  -42.6802,
  -42.6741,
  -42.6695,
  -42.6665,
  -42.6634,
  -42.6619,
  -42.6599,
  -42.6567,
  -42.6517,
  -42.6444,
  -42.6343,
  -42.6208,
  -42.6038,
  -42.5827,
  -42.5571,
  -42.5274,
  -42.4929,
  -42.4533,
  -42.4081,
  -42.3573,
  -42.3005,
  -42.2376,
  -42.168,
  -42.0914,
  -42.0074,
  -41.9161,
  -41.8173,
  -41.7117,
  -41.6011,
  -41.4878,
  -41.3749,
  -41.2649,
  -41.1597,
  -41.0621,
  -40.9714,
  -40.8874,
  -40.8102,
  -38.6428,
  -38.6912,
  -38.7387,
  -38.7849,
  -38.83,
  -38.873,
  -38.9163,
  -38.9591,
  -39.002,
  -39.0453,
  -39.0893,
  -39.1335,
  -39.178,
  -39.2221,
  -39.2656,
  -39.308,
  -39.349,
  -39.3885,
  -39.4265,
  -39.4634,
  -39.4986,
  -39.5346,
  -39.5705,
  -39.606,
  -39.6409,
  -39.6742,
  -39.7055,
  -39.734,
  -39.7596,
  -39.7825,
  -39.8034,
  -39.8235,
  -39.8428,
  -39.8621,
  -39.8815,
  -39.9008,
  -39.9224,
  -39.9453,
  -39.9693,
  -39.9939,
  -40.0183,
  -40.0424,
  -40.0656,
  -40.0879,
  -40.1102,
  -40.1328,
  -40.156,
  -40.1797,
  -40.2038,
  -40.2277,
  -40.2509,
  -40.2721,
  -40.2934,
  -40.3139,
  -40.3336,
  -40.3528,
  -40.3717,
  -40.3899,
  -40.4079,
  -40.4258,
  -40.4436,
  -40.4617,
  -40.4792,
  -40.4968,
  -40.5147,
  -40.5332,
  -40.5522,
  -40.5712,
  -40.5895,
  -40.6089,
  -40.6284,
  -40.6487,
  -40.6696,
  -40.6915,
  -40.7139,
  -40.7369,
  -40.7608,
  -40.7854,
  -40.8109,
  -40.8373,
  -40.864,
  -40.8904,
  -40.916,
  -40.9411,
  -40.9649,
  -40.9871,
  -41.01,
  -41.0333,
  -41.0569,
  -41.081,
  -41.1059,
  -41.1315,
  -41.1573,
  -41.1827,
  -41.2075,
  -41.2312,
  -41.2541,
  -41.2766,
  -41.299,
  -41.3218,
  -41.3451,
  -41.3684,
  -41.392,
  -41.414,
  -41.4363,
  -41.4576,
  -41.4775,
  -41.4966,
  -41.5146,
  -41.5309,
  -41.5457,
  -41.5588,
  -41.5698,
  -41.5787,
  -41.5856,
  -41.5908,
  -41.5947,
  -41.5976,
  -41.6005,
  -41.6026,
  -41.6042,
  -41.6049,
  -41.6053,
  -41.6048,
  -41.6054,
  -41.6072,
  -41.6095,
  -41.6135,
  -41.6186,
  -41.6248,
  -41.6322,
  -41.6407,
  -41.6503,
  -41.6609,
  -41.6721,
  -41.684,
  -41.6961,
  -41.7083,
  -41.72,
  -41.7317,
  -41.7435,
  -41.7556,
  -41.7685,
  -41.7822,
  -41.7956,
  -41.8103,
  -41.8245,
  -41.8382,
  -41.8509,
  -41.8625,
  -41.8734,
  -41.8838,
  -41.8941,
  -41.9047,
  -41.9159,
  -41.9277,
  -41.9399,
  -41.9523,
  -41.9647,
  -41.9773,
  -41.9898,
  -42.002,
  -42.0144,
  -42.0278,
  -42.0424,
  -42.0591,
  -42.0783,
  -42.0989,
  -42.1225,
  -42.1471,
  -42.1721,
  -42.1963,
  -42.2188,
  -42.2394,
  -42.2583,
  -42.2759,
  -42.293,
  -42.3098,
  -42.327,
  -42.3453,
  -42.3643,
  -42.3842,
  -42.4042,
  -42.4239,
  -42.4427,
  -42.4604,
  -42.4771,
  -42.493,
  -42.5084,
  -42.523,
  -42.5369,
  -42.5496,
  -42.5596,
  -42.5688,
  -42.5758,
  -42.5807,
  -42.5841,
  -42.5867,
  -42.5889,
  -42.5912,
  -42.5937,
  -42.5964,
  -42.5989,
  -42.6011,
  -42.6027,
  -42.603,
  -42.6021,
  -42.6,
  -42.5968,
  -42.5925,
  -42.5872,
  -42.5809,
  -42.5744,
  -42.5677,
  -42.5613,
  -42.5554,
  -42.5496,
  -42.544,
  -42.5382,
  -42.5328,
  -42.5286,
  -42.5249,
  -42.5249,
  -42.5271,
  -42.5318,
  -42.5384,
  -42.5466,
  -42.5555,
  -42.5646,
  -42.5738,
  -42.5826,
  -42.5907,
  -42.5981,
  -42.6048,
  -42.6105,
  -42.6158,
  -42.6208,
  -42.626,
  -42.6317,
  -42.6377,
  -42.6439,
  -42.6499,
  -42.6566,
  -42.6629,
  -42.6686,
  -42.6738,
  -42.6784,
  -42.6827,
  -42.6865,
  -42.6894,
  -42.6924,
  -42.6941,
  -42.6948,
  -42.6947,
  -42.6932,
  -42.6901,
  -42.6867,
  -42.6823,
  -42.6772,
  -42.6708,
  -42.664,
  -42.6562,
  -42.648,
  -42.6397,
  -42.632,
  -42.6253,
  -42.6204,
  -42.617,
  -42.6146,
  -42.6127,
  -42.6105,
  -42.6073,
  -42.6026,
  -42.5957,
  -42.5859,
  -42.5729,
  -42.5562,
  -42.5356,
  -42.5108,
  -42.4818,
  -42.4483,
  -42.4095,
  -42.3652,
  -42.3156,
  -42.2599,
  -42.1983,
  -42.1303,
  -42.0552,
  -41.9732,
  -41.8841,
  -41.7879,
  -41.6852,
  -41.5778,
  -41.4678,
  -41.3579,
  -41.2505,
  -41.1475,
  -41.0518,
  -40.9638,
  -40.8812,
  -40.8059,
  -38.4907,
  -38.5374,
  -38.5838,
  -38.629,
  -38.6732,
  -38.7166,
  -38.7592,
  -38.8017,
  -38.8444,
  -38.8875,
  -38.9311,
  -38.9752,
  -39.019,
  -39.0625,
  -39.1054,
  -39.1464,
  -39.1872,
  -39.2266,
  -39.2646,
  -39.3015,
  -39.3376,
  -39.3733,
  -39.4085,
  -39.4434,
  -39.4776,
  -39.5103,
  -39.5413,
  -39.5699,
  -39.5957,
  -39.6188,
  -39.6391,
  -39.6594,
  -39.6791,
  -39.6988,
  -39.7192,
  -39.7406,
  -39.7635,
  -39.7879,
  -39.8136,
  -39.8398,
  -39.8657,
  -39.8909,
  -39.9149,
  -39.9382,
  -39.9615,
  -39.9853,
  -40.0087,
  -40.0338,
  -40.0593,
  -40.0846,
  -40.1091,
  -40.1326,
  -40.155,
  -40.1763,
  -40.1967,
  -40.2163,
  -40.2356,
  -40.2544,
  -40.2733,
  -40.2924,
  -40.3113,
  -40.3302,
  -40.3479,
  -40.367,
  -40.3859,
  -40.4053,
  -40.4252,
  -40.4452,
  -40.4654,
  -40.4858,
  -40.5067,
  -40.5281,
  -40.5503,
  -40.5732,
  -40.5967,
  -40.6207,
  -40.6452,
  -40.6708,
  -40.6972,
  -40.7233,
  -40.7507,
  -40.7778,
  -40.8038,
  -40.8289,
  -40.8532,
  -40.8771,
  -40.901,
  -40.9251,
  -40.9496,
  -40.9745,
  -40.9998,
  -41.0256,
  -41.0517,
  -41.0779,
  -41.1036,
  -41.1285,
  -41.1523,
  -41.1745,
  -41.1973,
  -41.2206,
  -41.2445,
  -41.2684,
  -41.2926,
  -41.3163,
  -41.3393,
  -41.361,
  -41.3809,
  -41.3999,
  -41.4173,
  -41.4328,
  -41.447,
  -41.4594,
  -41.4697,
  -41.4786,
  -41.4851,
  -41.4904,
  -41.4927,
  -41.4948,
  -41.4967,
  -41.4981,
  -41.4991,
  -41.4998,
  -41.5,
  -41.5004,
  -41.5013,
  -41.5028,
  -41.5057,
  -41.5097,
  -41.5147,
  -41.521,
  -41.5282,
  -41.5365,
  -41.5457,
  -41.5559,
  -41.5668,
  -41.5783,
  -41.5905,
  -41.6019,
  -41.6141,
  -41.6262,
  -41.6379,
  -41.6497,
  -41.6623,
  -41.6757,
  -41.6897,
  -41.704,
  -41.7182,
  -41.7317,
  -41.7442,
  -41.7557,
  -41.7666,
  -41.7771,
  -41.7878,
  -41.7988,
  -41.8105,
  -41.8224,
  -41.8348,
  -41.8477,
  -41.861,
  -41.8734,
  -41.8864,
  -41.8995,
  -41.9125,
  -41.9264,
  -41.9415,
  -41.9585,
  -41.9778,
  -41.9993,
  -42.0228,
  -42.0471,
  -42.0717,
  -42.0953,
  -42.1176,
  -42.1381,
  -42.157,
  -42.1748,
  -42.192,
  -42.2093,
  -42.2271,
  -42.246,
  -42.2655,
  -42.2857,
  -42.3057,
  -42.3244,
  -42.343,
  -42.3611,
  -42.379,
  -42.3963,
  -42.4136,
  -42.43,
  -42.4455,
  -42.4595,
  -42.4718,
  -42.4817,
  -42.4895,
  -42.4955,
  -42.5001,
  -42.5041,
  -42.5077,
  -42.5114,
  -42.515,
  -42.519,
  -42.5228,
  -42.5261,
  -42.5284,
  -42.5292,
  -42.5285,
  -42.5265,
  -42.5236,
  -42.5196,
  -42.5147,
  -42.5081,
  -42.5025,
  -42.4966,
  -42.4912,
  -42.4862,
  -42.4812,
  -42.4761,
  -42.4704,
  -42.4651,
  -42.4609,
  -42.4587,
  -42.4588,
  -42.4618,
  -42.4676,
  -42.4755,
  -42.4847,
  -42.4944,
  -42.5043,
  -42.5139,
  -42.5227,
  -42.5309,
  -42.5384,
  -42.5449,
  -42.5509,
  -42.5565,
  -42.5619,
  -42.5673,
  -42.573,
  -42.5788,
  -42.5848,
  -42.591,
  -42.5965,
  -42.6029,
  -42.6087,
  -42.6143,
  -42.6195,
  -42.6243,
  -42.6291,
  -42.6333,
  -42.637,
  -42.6395,
  -42.6414,
  -42.6426,
  -42.6424,
  -42.6411,
  -42.6386,
  -42.635,
  -42.6304,
  -42.6244,
  -42.6174,
  -42.6096,
  -42.6008,
  -42.5922,
  -42.5842,
  -42.5774,
  -42.5724,
  -42.5687,
  -42.5658,
  -42.5634,
  -42.5608,
  -42.5574,
  -42.5526,
  -42.5457,
  -42.5363,
  -42.5237,
  -42.5076,
  -42.4877,
  -42.4639,
  -42.4358,
  -42.4032,
  -42.3652,
  -42.321,
  -42.2719,
  -42.2175,
  -42.1575,
  -42.0914,
  -42.0189,
  -41.9396,
  -41.8533,
  -41.7603,
  -41.6608,
  -41.5564,
  -41.4492,
  -41.3413,
  -41.2357,
  -41.1348,
  -41.0403,
  -40.9524,
  -40.8724,
  -40.7985,
  -38.336,
  -38.3827,
  -38.4282,
  -38.4726,
  -38.5161,
  -38.5593,
  -38.6019,
  -38.6446,
  -38.6876,
  -38.7307,
  -38.7734,
  -38.8167,
  -38.8599,
  -38.9027,
  -38.9448,
  -38.9861,
  -39.0264,
  -39.0657,
  -39.1038,
  -39.1407,
  -39.1768,
  -39.2122,
  -39.247,
  -39.2811,
  -39.3143,
  -39.3457,
  -39.3763,
  -39.4047,
  -39.4308,
  -39.4543,
  -39.4761,
  -39.4967,
  -39.5169,
  -39.5375,
  -39.559,
  -39.5818,
  -39.6059,
  -39.6318,
  -39.6589,
  -39.6865,
  -39.7125,
  -39.7385,
  -39.7635,
  -39.7876,
  -39.8119,
  -39.8367,
  -39.8623,
  -39.8887,
  -39.9155,
  -39.9422,
  -39.9682,
  -39.9929,
  -40.0163,
  -40.0385,
  -40.0595,
  -40.0796,
  -40.0982,
  -40.1177,
  -40.1375,
  -40.1574,
  -40.1773,
  -40.1971,
  -40.2172,
  -40.2372,
  -40.2575,
  -40.278,
  -40.2986,
  -40.3194,
  -40.3405,
  -40.362,
  -40.3842,
  -40.4071,
  -40.4307,
  -40.4539,
  -40.4786,
  -40.5034,
  -40.5288,
  -40.5549,
  -40.582,
  -40.6097,
  -40.6375,
  -40.6649,
  -40.6917,
  -40.7175,
  -40.7422,
  -40.7667,
  -40.7915,
  -40.8165,
  -40.8417,
  -40.8673,
  -40.8936,
  -40.9187,
  -40.9447,
  -40.9713,
  -40.9976,
  -41.0235,
  -41.0485,
  -41.0728,
  -41.0966,
  -41.1204,
  -41.1446,
  -41.169,
  -41.1939,
  -41.2183,
  -41.2417,
  -41.2637,
  -41.2841,
  -41.3027,
  -41.3198,
  -41.3349,
  -41.3475,
  -41.3593,
  -41.3694,
  -41.3775,
  -41.3838,
  -41.3891,
  -41.3924,
  -41.3941,
  -41.3951,
  -41.3959,
  -41.3963,
  -41.3966,
  -41.397,
  -41.3972,
  -41.398,
  -41.3998,
  -41.4026,
  -41.4067,
  -41.412,
  -41.4179,
  -41.424,
  -41.4318,
  -41.4408,
  -41.4508,
  -41.4616,
  -41.473,
  -41.4851,
  -41.4976,
  -41.5101,
  -41.5225,
  -41.5343,
  -41.5462,
  -41.5584,
  -41.5715,
  -41.5852,
  -41.5992,
  -41.6133,
  -41.6265,
  -41.639,
  -41.6505,
  -41.6616,
  -41.6714,
  -41.6826,
  -41.6943,
  -41.7065,
  -41.7189,
  -41.732,
  -41.7458,
  -41.76,
  -41.7743,
  -41.7884,
  -41.8021,
  -41.8158,
  -41.8299,
  -41.8454,
  -41.8627,
  -41.8819,
  -41.9034,
  -41.9263,
  -41.9501,
  -41.9735,
  -41.9962,
  -42.018,
  -42.0382,
  -42.0572,
  -42.0743,
  -42.0921,
  -42.1098,
  -42.1279,
  -42.1469,
  -42.1669,
  -42.1869,
  -42.2065,
  -42.2257,
  -42.2445,
  -42.2631,
  -42.2817,
  -42.3009,
  -42.3199,
  -42.3383,
  -42.3556,
  -42.3711,
  -42.3839,
  -42.3946,
  -42.4034,
  -42.4105,
  -42.4161,
  -42.4213,
  -42.4264,
  -42.4317,
  -42.4366,
  -42.4407,
  -42.4453,
  -42.4495,
  -42.4521,
  -42.453,
  -42.4522,
  -42.4504,
  -42.4476,
  -42.4441,
  -42.4401,
  -42.4357,
  -42.4309,
  -42.426,
  -42.4214,
  -42.417,
  -42.4125,
  -42.4075,
  -42.4023,
  -42.3974,
  -42.3936,
  -42.3915,
  -42.3921,
  -42.3956,
  -42.4022,
  -42.411,
  -42.4212,
  -42.4322,
  -42.4427,
  -42.4527,
  -42.4622,
  -42.4695,
  -42.4767,
  -42.4832,
  -42.4894,
  -42.4955,
  -42.5012,
  -42.5068,
  -42.5123,
  -42.5177,
  -42.5236,
  -42.5296,
  -42.5359,
  -42.542,
  -42.5481,
  -42.5541,
  -42.56,
  -42.5656,
  -42.5713,
  -42.5765,
  -42.5814,
  -42.5853,
  -42.5885,
  -42.5906,
  -42.5915,
  -42.5913,
  -42.5898,
  -42.587,
  -42.5828,
  -42.5771,
  -42.5703,
  -42.5622,
  -42.5535,
  -42.5447,
  -42.5369,
  -42.5302,
  -42.5251,
  -42.5212,
  -42.5169,
  -42.514,
  -42.5108,
  -42.5069,
  -42.502,
  -42.4952,
  -42.4858,
  -42.4732,
  -42.4575,
  -42.4383,
  -42.4153,
  -42.3884,
  -42.3567,
  -42.3197,
  -42.2772,
  -42.2291,
  -42.1763,
  -42.1182,
  -42.0546,
  -41.9848,
  -41.9088,
  -41.8259,
  -41.7361,
  -41.64,
  -41.5385,
  -41.4337,
  -41.328,
  -41.2238,
  -41.1233,
  -41.0286,
  -40.9407,
  -40.8605,
  -40.7868,
  -38.1803,
  -38.226,
  -38.2706,
  -38.3142,
  -38.3576,
  -38.4008,
  -38.4433,
  -38.4869,
  -38.5307,
  -38.5742,
  -38.6176,
  -38.6608,
  -38.7034,
  -38.7452,
  -38.7861,
  -38.8265,
  -38.8663,
  -38.9053,
  -38.9434,
  -38.9805,
  -39.0158,
  -39.0511,
  -39.0855,
  -39.1189,
  -39.1514,
  -39.1828,
  -39.2129,
  -39.2411,
  -39.2675,
  -39.2915,
  -39.3139,
  -39.3353,
  -39.3564,
  -39.3779,
  -39.4005,
  -39.4235,
  -39.4491,
  -39.4763,
  -39.5048,
  -39.5334,
  -39.5615,
  -39.5884,
  -39.6141,
  -39.6392,
  -39.6644,
  -39.6901,
  -39.7166,
  -39.744,
  -39.7719,
  -39.7997,
  -39.8268,
  -39.8516,
  -39.8761,
  -39.8992,
  -39.9209,
  -39.9416,
  -39.9619,
  -39.9821,
  -40.0025,
  -40.0233,
  -40.0441,
  -40.0649,
  -40.086,
  -40.1072,
  -40.1288,
  -40.1503,
  -40.1719,
  -40.1933,
  -40.2142,
  -40.2369,
  -40.2607,
  -40.2852,
  -40.3105,
  -40.336,
  -40.3617,
  -40.3875,
  -40.4134,
  -40.44,
  -40.4674,
  -40.4952,
  -40.5237,
  -40.5515,
  -40.5788,
  -40.6056,
  -40.6317,
  -40.6564,
  -40.6817,
  -40.7076,
  -40.7334,
  -40.7596,
  -40.7858,
  -40.8123,
  -40.8387,
  -40.8652,
  -40.8918,
  -40.9184,
  -40.9443,
  -40.9698,
  -40.9947,
  -41.0193,
  -41.0439,
  -41.0687,
  -41.0939,
  -41.1177,
  -41.1418,
  -41.1642,
  -41.1849,
  -41.2035,
  -41.2204,
  -41.2353,
  -41.2487,
  -41.2601,
  -41.2697,
  -41.2778,
  -41.2842,
  -41.289,
  -41.292,
  -41.2936,
  -41.2944,
  -41.2946,
  -41.2949,
  -41.2951,
  -41.2953,
  -41.295,
  -41.2959,
  -41.2977,
  -41.3006,
  -41.3043,
  -41.309,
  -41.3146,
  -41.3213,
  -41.3291,
  -41.338,
  -41.3481,
  -41.3586,
  -41.37,
  -41.382,
  -41.3945,
  -41.4072,
  -41.4199,
  -41.432,
  -41.4439,
  -41.4561,
  -41.4688,
  -41.4812,
  -41.495,
  -41.5087,
  -41.5221,
  -41.5346,
  -41.5464,
  -41.558,
  -41.5694,
  -41.5811,
  -41.5934,
  -41.6062,
  -41.6192,
  -41.6332,
  -41.6481,
  -41.6636,
  -41.6791,
  -41.6939,
  -41.7081,
  -41.7223,
  -41.7369,
  -41.7528,
  -41.7702,
  -41.7895,
  -41.8095,
  -41.8318,
  -41.8544,
  -41.8767,
  -41.8984,
  -41.9195,
  -41.9398,
  -41.9588,
  -41.9773,
  -41.9953,
  -42.0133,
  -42.032,
  -42.0513,
  -42.0712,
  -42.0909,
  -42.11,
  -42.1287,
  -42.1471,
  -42.1659,
  -42.1859,
  -42.2065,
  -42.2276,
  -42.2479,
  -42.2666,
  -42.2832,
  -42.2962,
  -42.3079,
  -42.3176,
  -42.3255,
  -42.3323,
  -42.3384,
  -42.3448,
  -42.3512,
  -42.3575,
  -42.3636,
  -42.369,
  -42.3733,
  -42.3761,
  -42.3768,
  -42.376,
  -42.3738,
  -42.3712,
  -42.3685,
  -42.3654,
  -42.362,
  -42.3584,
  -42.3548,
  -42.3511,
  -42.3472,
  -42.3428,
  -42.3382,
  -42.3334,
  -42.3288,
  -42.3254,
  -42.3229,
  -42.324,
  -42.328,
  -42.3352,
  -42.3448,
  -42.356,
  -42.3678,
  -42.3793,
  -42.3901,
  -42.3998,
  -42.4079,
  -42.4152,
  -42.4217,
  -42.4282,
  -42.4346,
  -42.4406,
  -42.4463,
  -42.4518,
  -42.4574,
  -42.4629,
  -42.4685,
  -42.4744,
  -42.4805,
  -42.4865,
  -42.4928,
  -42.4991,
  -42.5054,
  -42.512,
  -42.5185,
  -42.5245,
  -42.5299,
  -42.5345,
  -42.5379,
  -42.5401,
  -42.5399,
  -42.5395,
  -42.5375,
  -42.5339,
  -42.5287,
  -42.5218,
  -42.5137,
  -42.505,
  -42.4966,
  -42.4891,
  -42.4828,
  -42.4779,
  -42.4736,
  -42.47,
  -42.4664,
  -42.4626,
  -42.4582,
  -42.453,
  -42.4461,
  -42.4369,
  -42.4245,
  -42.4091,
  -42.3904,
  -42.3681,
  -42.3418,
  -42.3109,
  -42.2748,
  -42.2331,
  -42.1862,
  -42.1347,
  -42.0789,
  -42.018,
  -41.9517,
  -41.8791,
  -41.7998,
  -41.7136,
  -41.6208,
  -41.5222,
  -41.4199,
  -41.3161,
  -41.2127,
  -41.1122,
  -41.0166,
  -40.9273,
  -40.8445,
  -40.7698,
  -38.0232,
  -38.0668,
  -38.1106,
  -38.154,
  -38.1975,
  -38.2414,
  -38.286,
  -38.3304,
  -38.3746,
  -38.4187,
  -38.4623,
  -38.5051,
  -38.5471,
  -38.588,
  -38.6281,
  -38.6667,
  -38.706,
  -38.7448,
  -38.7829,
  -38.8203,
  -38.8567,
  -38.892,
  -38.9262,
  -38.9592,
  -38.991,
  -39.0216,
  -39.051,
  -39.0791,
  -39.1056,
  -39.1299,
  -39.152,
  -39.1741,
  -39.1961,
  -39.2189,
  -39.2429,
  -39.2683,
  -39.2953,
  -39.3238,
  -39.3534,
  -39.383,
  -39.4119,
  -39.4398,
  -39.4663,
  -39.4924,
  -39.5184,
  -39.545,
  -39.5715,
  -39.5996,
  -39.6282,
  -39.6572,
  -39.6851,
  -39.7118,
  -39.7371,
  -39.761,
  -39.7836,
  -39.805,
  -39.8259,
  -39.8468,
  -39.8679,
  -39.8893,
  -39.9108,
  -39.9325,
  -39.9534,
  -39.9757,
  -39.9983,
  -40.0208,
  -40.0434,
  -40.066,
  -40.0892,
  -40.1133,
  -40.1384,
  -40.1645,
  -40.1914,
  -40.2182,
  -40.2448,
  -40.2714,
  -40.2978,
  -40.325,
  -40.3531,
  -40.3805,
  -40.4091,
  -40.4376,
  -40.4658,
  -40.4935,
  -40.5205,
  -40.5473,
  -40.5739,
  -40.6001,
  -40.6264,
  -40.6525,
  -40.6787,
  -40.7051,
  -40.7321,
  -40.7593,
  -40.7862,
  -40.8132,
  -40.8398,
  -40.8648,
  -40.8904,
  -40.9156,
  -40.9407,
  -40.9658,
  -40.991,
  -41.016,
  -41.0401,
  -41.0628,
  -41.084,
  -41.1032,
  -41.1203,
  -41.1354,
  -41.1488,
  -41.1603,
  -41.1699,
  -41.1779,
  -41.1843,
  -41.1889,
  -41.1908,
  -41.1924,
  -41.193,
  -41.1931,
  -41.1932,
  -41.1935,
  -41.1941,
  -41.1949,
  -41.1961,
  -41.1979,
  -41.2004,
  -41.2035,
  -41.2076,
  -41.2126,
  -41.2189,
  -41.2266,
  -41.2357,
  -41.2459,
  -41.2566,
  -41.2679,
  -41.2799,
  -41.2915,
  -41.3043,
  -41.3172,
  -41.3296,
  -41.3417,
  -41.3539,
  -41.3666,
  -41.38,
  -41.3939,
  -41.4077,
  -41.4209,
  -41.4336,
  -41.4459,
  -41.4581,
  -41.4702,
  -41.4824,
  -41.4952,
  -41.5084,
  -41.5226,
  -41.5376,
  -41.5536,
  -41.5704,
  -41.5858,
  -41.6013,
  -41.6163,
  -41.6308,
  -41.6458,
  -41.6618,
  -41.6796,
  -41.6987,
  -41.719,
  -41.7401,
  -41.7615,
  -41.7826,
  -41.8034,
  -41.824,
  -41.8441,
  -41.8636,
  -41.8824,
  -41.9009,
  -41.9196,
  -41.9388,
  -41.9584,
  -41.9781,
  -41.9975,
  -42.0162,
  -42.033,
  -42.0513,
  -42.0707,
  -42.0915,
  -42.1136,
  -42.1361,
  -42.1579,
  -42.1779,
  -42.1954,
  -42.2106,
  -42.2231,
  -42.2334,
  -42.2422,
  -42.2499,
  -42.2571,
  -42.2645,
  -42.2723,
  -42.2799,
  -42.2866,
  -42.2926,
  -42.2972,
  -42.2999,
  -42.3003,
  -42.2993,
  -42.2974,
  -42.2949,
  -42.2924,
  -42.29,
  -42.2866,
  -42.2842,
  -42.2818,
  -42.2789,
  -42.2755,
  -42.2716,
  -42.267,
  -42.2626,
  -42.2586,
  -42.2557,
  -42.255,
  -42.2566,
  -42.2612,
  -42.2688,
  -42.2791,
  -42.2909,
  -42.3039,
  -42.3163,
  -42.3274,
  -42.3368,
  -42.3451,
  -42.3523,
  -42.3594,
  -42.3661,
  -42.3727,
  -42.379,
  -42.3852,
  -42.391,
  -42.3966,
  -42.4019,
  -42.4072,
  -42.4124,
  -42.4171,
  -42.4231,
  -42.4294,
  -42.4361,
  -42.4435,
  -42.4509,
  -42.4585,
  -42.4659,
  -42.473,
  -42.4792,
  -42.4839,
  -42.4873,
  -42.4893,
  -42.4897,
  -42.4886,
  -42.4857,
  -42.4809,
  -42.4743,
  -42.4664,
  -42.4581,
  -42.4503,
  -42.4433,
  -42.4375,
  -42.4328,
  -42.4284,
  -42.4241,
  -42.42,
  -42.4157,
  -42.4109,
  -42.4054,
  -42.3986,
  -42.3894,
  -42.3772,
  -42.3619,
  -42.3434,
  -42.3213,
  -42.2953,
  -42.265,
  -42.2296,
  -42.188,
  -42.1426,
  -42.0928,
  -42.0388,
  -41.9806,
  -41.9175,
  -41.8485,
  -41.7727,
  -41.6902,
  -41.6009,
  -41.5054,
  -41.4055,
  -41.3035,
  -41.201,
  -41.0999,
  -41.0026,
  -40.9114,
  -40.827,
  -40.7505,
  -37.8647,
  -37.9082,
  -37.9513,
  -37.9946,
  -38.0385,
  -38.0829,
  -38.128,
  -38.1733,
  -38.2183,
  -38.2627,
  -38.3053,
  -38.3479,
  -38.3893,
  -38.4298,
  -38.4694,
  -38.5086,
  -38.5476,
  -38.5863,
  -38.6245,
  -38.662,
  -38.6986,
  -38.7342,
  -38.7682,
  -38.801,
  -38.8324,
  -38.8616,
  -38.8907,
  -38.9185,
  -38.9445,
  -38.9691,
  -38.9928,
  -39.0157,
  -39.0389,
  -39.0628,
  -39.088,
  -39.1146,
  -39.143,
  -39.1727,
  -39.2033,
  -39.234,
  -39.2638,
  -39.2916,
  -39.3192,
  -39.3463,
  -39.3735,
  -39.4008,
  -39.4289,
  -39.4576,
  -39.4871,
  -39.5164,
  -39.5452,
  -39.5727,
  -39.5988,
  -39.6234,
  -39.6467,
  -39.6689,
  -39.6906,
  -39.7111,
  -39.7328,
  -39.7548,
  -39.7769,
  -39.7993,
  -39.8219,
  -39.8451,
  -39.8685,
  -39.892,
  -39.9155,
  -39.9396,
  -39.9642,
  -39.9899,
  -40.0166,
  -40.0441,
  -40.0722,
  -40.0992,
  -40.1268,
  -40.1541,
  -40.1812,
  -40.2089,
  -40.2375,
  -40.2667,
  -40.2962,
  -40.3257,
  -40.3546,
  -40.3831,
  -40.4111,
  -40.4387,
  -40.4657,
  -40.4926,
  -40.5188,
  -40.5449,
  -40.5711,
  -40.5968,
  -40.6243,
  -40.6519,
  -40.6797,
  -40.7072,
  -40.7342,
  -40.7606,
  -40.7864,
  -40.8116,
  -40.8366,
  -40.8617,
  -40.8869,
  -40.9119,
  -40.9358,
  -40.959,
  -40.9804,
  -41,
  -41.0179,
  -41.0338,
  -41.0468,
  -41.0587,
  -41.0686,
  -41.0764,
  -41.0827,
  -41.0871,
  -41.0899,
  -41.0914,
  -41.092,
  -41.0924,
  -41.0927,
  -41.0931,
  -41.0941,
  -41.0955,
  -41.0971,
  -41.0991,
  -41.1014,
  -41.1041,
  -41.1073,
  -41.1117,
  -41.1167,
  -41.1241,
  -41.1331,
  -41.1431,
  -41.1539,
  -41.1655,
  -41.1774,
  -41.1901,
  -41.2033,
  -41.2165,
  -41.2292,
  -41.2416,
  -41.254,
  -41.2668,
  -41.2803,
  -41.2944,
  -41.3086,
  -41.3223,
  -41.3354,
  -41.3481,
  -41.3608,
  -41.3722,
  -41.3852,
  -41.3986,
  -41.4127,
  -41.4277,
  -41.4439,
  -41.461,
  -41.4785,
  -41.4954,
  -41.5118,
  -41.5274,
  -41.5423,
  -41.5579,
  -41.5741,
  -41.5915,
  -41.6102,
  -41.6295,
  -41.6495,
  -41.6699,
  -41.6899,
  -41.7099,
  -41.7299,
  -41.7499,
  -41.7699,
  -41.7884,
  -41.8077,
  -41.8271,
  -41.8467,
  -41.8667,
  -41.8863,
  -41.9055,
  -41.9236,
  -41.9412,
  -41.9593,
  -41.9792,
  -42.0009,
  -42.0241,
  -42.0477,
  -42.0705,
  -42.0917,
  -42.1103,
  -42.1264,
  -42.1398,
  -42.1506,
  -42.1598,
  -42.1681,
  -42.1764,
  -42.1849,
  -42.1937,
  -42.2023,
  -42.2088,
  -42.2151,
  -42.2198,
  -42.2225,
  -42.2229,
  -42.2218,
  -42.2198,
  -42.2172,
  -42.215,
  -42.2131,
  -42.2115,
  -42.2101,
  -42.2087,
  -42.2067,
  -42.204,
  -42.2004,
  -42.1963,
  -42.1925,
  -42.1892,
  -42.1874,
  -42.1873,
  -42.1895,
  -42.1948,
  -42.2028,
  -42.2136,
  -42.2262,
  -42.2395,
  -42.2521,
  -42.2632,
  -42.2727,
  -42.2801,
  -42.2876,
  -42.2947,
  -42.3017,
  -42.309,
  -42.3161,
  -42.3229,
  -42.3291,
  -42.3346,
  -42.3399,
  -42.3446,
  -42.3495,
  -42.3546,
  -42.3604,
  -42.3666,
  -42.3736,
  -42.3814,
  -42.3899,
  -42.3989,
  -42.4079,
  -42.4165,
  -42.4243,
  -42.4305,
  -42.4351,
  -42.4381,
  -42.4396,
  -42.4392,
  -42.4371,
  -42.433,
  -42.4271,
  -42.4199,
  -42.4125,
  -42.4053,
  -42.3988,
  -42.3933,
  -42.3884,
  -42.3837,
  -42.378,
  -42.3733,
  -42.3687,
  -42.3638,
  -42.3583,
  -42.3517,
  -42.3427,
  -42.3309,
  -42.3156,
  -42.297,
  -42.2747,
  -42.2487,
  -42.2184,
  -42.1835,
  -42.1438,
  -42.0995,
  -42.0515,
  -41.9993,
  -41.9438,
  -41.8834,
  -41.8177,
  -41.7454,
  -41.6665,
  -41.5808,
  -41.4885,
  -41.3914,
  -41.2911,
  -41.1892,
  -41.0877,
  -40.9886,
  -40.8947,
  -40.8078,
  -40.7285,
  -37.7069,
  -37.7495,
  -37.7922,
  -37.8355,
  -37.8799,
  -37.9248,
  -37.9692,
  -38.0148,
  -38.06,
  -38.1044,
  -38.1477,
  -38.1903,
  -38.2316,
  -38.2719,
  -38.3116,
  -38.3508,
  -38.3896,
  -38.4284,
  -38.4668,
  -38.5045,
  -38.5403,
  -38.5759,
  -38.6102,
  -38.643,
  -38.6742,
  -38.7042,
  -38.7329,
  -38.7604,
  -38.7867,
  -38.8114,
  -38.8354,
  -38.8591,
  -38.8832,
  -38.9081,
  -38.9344,
  -38.9612,
  -38.9906,
  -39.0214,
  -39.053,
  -39.0846,
  -39.1154,
  -39.1453,
  -39.174,
  -39.2024,
  -39.2307,
  -39.259,
  -39.2877,
  -39.3172,
  -39.3472,
  -39.377,
  -39.4064,
  -39.4335,
  -39.4602,
  -39.4856,
  -39.5096,
  -39.5326,
  -39.5552,
  -39.5774,
  -39.5997,
  -39.6222,
  -39.6448,
  -39.6677,
  -39.691,
  -39.7148,
  -39.739,
  -39.7633,
  -39.788,
  -39.8132,
  -39.8384,
  -39.8658,
  -39.8943,
  -39.9233,
  -39.9522,
  -39.981,
  -40.0093,
  -40.0373,
  -40.0652,
  -40.0938,
  -40.1231,
  -40.153,
  -40.1834,
  -40.2139,
  -40.244,
  -40.2734,
  -40.3021,
  -40.3291,
  -40.3563,
  -40.3828,
  -40.4089,
  -40.4352,
  -40.4618,
  -40.4888,
  -40.5169,
  -40.5452,
  -40.5737,
  -40.602,
  -40.6296,
  -40.6562,
  -40.6819,
  -40.7067,
  -40.7311,
  -40.7556,
  -40.7803,
  -40.8042,
  -40.8287,
  -40.852,
  -40.8743,
  -40.8946,
  -40.9133,
  -40.9303,
  -40.9451,
  -40.9579,
  -40.9682,
  -40.9763,
  -40.9822,
  -40.986,
  -40.9882,
  -40.9894,
  -40.9901,
  -40.9908,
  -40.9917,
  -40.9929,
  -40.9943,
  -40.9951,
  -40.9971,
  -40.9993,
  -41.0017,
  -41.0044,
  -41.0076,
  -41.0116,
  -41.017,
  -41.024,
  -41.0328,
  -41.0427,
  -41.0534,
  -41.065,
  -41.077,
  -41.0897,
  -41.1031,
  -41.1165,
  -41.1296,
  -41.1424,
  -41.1554,
  -41.1687,
  -41.1816,
  -41.1961,
  -41.2105,
  -41.2247,
  -41.2384,
  -41.2519,
  -41.2651,
  -41.2784,
  -41.2918,
  -41.3056,
  -41.3202,
  -41.3362,
  -41.3532,
  -41.3707,
  -41.3891,
  -41.4068,
  -41.4238,
  -41.4397,
  -41.4552,
  -41.471,
  -41.4874,
  -41.5045,
  -41.5224,
  -41.54,
  -41.5591,
  -41.5784,
  -41.5974,
  -41.6165,
  -41.636,
  -41.6561,
  -41.6761,
  -41.696,
  -41.7163,
  -41.7365,
  -41.7572,
  -41.7778,
  -41.7974,
  -41.816,
  -41.8338,
  -41.8513,
  -41.8698,
  -41.8901,
  -41.9123,
  -41.9365,
  -41.9612,
  -41.9852,
  -42.0073,
  -42.0266,
  -42.0423,
  -42.0562,
  -42.0676,
  -42.0772,
  -42.0863,
  -42.0953,
  -42.1048,
  -42.1143,
  -42.1235,
  -42.1315,
  -42.1381,
  -42.1429,
  -42.1455,
  -42.146,
  -42.1447,
  -42.1427,
  -42.1404,
  -42.1382,
  -42.1368,
  -42.1363,
  -42.1362,
  -42.1355,
  -42.1346,
  -42.1324,
  -42.1291,
  -42.1256,
  -42.1224,
  -42.1199,
  -42.1191,
  -42.1189,
  -42.122,
  -42.1279,
  -42.1369,
  -42.1484,
  -42.1612,
  -42.1746,
  -42.1867,
  -42.1974,
  -42.2069,
  -42.2152,
  -42.2229,
  -42.2301,
  -42.2378,
  -42.246,
  -42.2537,
  -42.2611,
  -42.2679,
  -42.2736,
  -42.2787,
  -42.2834,
  -42.288,
  -42.2928,
  -42.2982,
  -42.3043,
  -42.3117,
  -42.3202,
  -42.3296,
  -42.3396,
  -42.3498,
  -42.36,
  -42.3693,
  -42.3769,
  -42.3829,
  -42.386,
  -42.3883,
  -42.389,
  -42.3877,
  -42.3845,
  -42.3795,
  -42.3732,
  -42.3664,
  -42.36,
  -42.3541,
  -42.3486,
  -42.3435,
  -42.3386,
  -42.3337,
  -42.3288,
  -42.3241,
  -42.3192,
  -42.314,
  -42.3078,
  -42.299,
  -42.2872,
  -42.2717,
  -42.2525,
  -42.2297,
  -42.2031,
  -42.1726,
  -42.138,
  -42.099,
  -42.0559,
  -42.0089,
  -41.959,
  -41.9054,
  -41.8478,
  -41.7849,
  -41.7158,
  -41.6406,
  -41.5584,
  -41.4697,
  -41.3756,
  -41.2774,
  -41.1765,
  -41.0743,
  -40.9736,
  -40.8769,
  -40.7858,
  -40.7037,
  -37.5495,
  -37.5904,
  -37.6328,
  -37.6762,
  -37.7205,
  -37.7657,
  -37.8111,
  -37.8563,
  -37.9011,
  -37.9452,
  -37.9888,
  -38.0316,
  -38.0732,
  -38.1135,
  -38.1533,
  -38.1918,
  -38.231,
  -38.2701,
  -38.3087,
  -38.3466,
  -38.3835,
  -38.4193,
  -38.4537,
  -38.4866,
  -38.5179,
  -38.548,
  -38.5766,
  -38.6041,
  -38.6303,
  -38.6555,
  -38.679,
  -38.7033,
  -38.7281,
  -38.754,
  -38.781,
  -38.8096,
  -38.8398,
  -38.8714,
  -38.9038,
  -38.9361,
  -38.9678,
  -38.9989,
  -39.0291,
  -39.0589,
  -39.0883,
  -39.1178,
  -39.1465,
  -39.1768,
  -39.2074,
  -39.2379,
  -39.2676,
  -39.2964,
  -39.3238,
  -39.3497,
  -39.3748,
  -39.3987,
  -39.4219,
  -39.4449,
  -39.4676,
  -39.4905,
  -39.5136,
  -39.5371,
  -39.5601,
  -39.5845,
  -39.6092,
  -39.6344,
  -39.6599,
  -39.6863,
  -39.7138,
  -39.7428,
  -39.7727,
  -39.8029,
  -39.8331,
  -39.8625,
  -39.8915,
  -39.92,
  -39.9491,
  -39.9786,
  -40.0089,
  -40.0387,
  -40.0699,
  -40.1013,
  -40.1323,
  -40.1625,
  -40.1916,
  -40.2195,
  -40.2465,
  -40.2727,
  -40.2987,
  -40.325,
  -40.3519,
  -40.3798,
  -40.4085,
  -40.4379,
  -40.4676,
  -40.4965,
  -40.5248,
  -40.5508,
  -40.5764,
  -40.6007,
  -40.6244,
  -40.6479,
  -40.6718,
  -40.6962,
  -40.7208,
  -40.7446,
  -40.7679,
  -40.7895,
  -40.8094,
  -40.8274,
  -40.8433,
  -40.8572,
  -40.8683,
  -40.8764,
  -40.8823,
  -40.8859,
  -40.8864,
  -40.8867,
  -40.8871,
  -40.8877,
  -40.889,
  -40.8907,
  -40.893,
  -40.8955,
  -40.8978,
  -40.9005,
  -40.9035,
  -40.9065,
  -40.9097,
  -40.9139,
  -40.9193,
  -40.926,
  -40.9343,
  -40.9439,
  -40.9543,
  -40.9658,
  -40.9781,
  -40.9898,
  -41.0032,
  -41.017,
  -41.0304,
  -41.0438,
  -41.0575,
  -41.0715,
  -41.086,
  -41.1008,
  -41.1155,
  -41.1301,
  -41.1445,
  -41.1586,
  -41.1726,
  -41.1866,
  -41.2007,
  -41.2152,
  -41.2305,
  -41.2468,
  -41.2642,
  -41.2826,
  -41.3011,
  -41.3184,
  -41.3357,
  -41.3519,
  -41.3678,
  -41.3838,
  -41.4001,
  -41.4168,
  -41.4342,
  -41.4522,
  -41.4702,
  -41.4884,
  -41.5066,
  -41.525,
  -41.5439,
  -41.5634,
  -41.5836,
  -41.604,
  -41.6253,
  -41.6466,
  -41.668,
  -41.6887,
  -41.7086,
  -41.7272,
  -41.7446,
  -41.7612,
  -41.78,
  -41.8009,
  -41.8241,
  -41.8493,
  -41.875,
  -41.8999,
  -41.9228,
  -41.9429,
  -41.9601,
  -41.9744,
  -41.9861,
  -41.9963,
  -42.0058,
  -42.0155,
  -42.0253,
  -42.0355,
  -42.0448,
  -42.0531,
  -42.0599,
  -42.0648,
  -42.0675,
  -42.0682,
  -42.067,
  -42.0651,
  -42.0628,
  -42.0612,
  -42.0603,
  -42.0596,
  -42.0605,
  -42.061,
  -42.0609,
  -42.0593,
  -42.057,
  -42.0542,
  -42.0517,
  -42.0503,
  -42.0503,
  -42.052,
  -42.056,
  -42.0628,
  -42.0726,
  -42.0844,
  -42.0971,
  -42.1099,
  -42.1216,
  -42.1321,
  -42.141,
  -42.1493,
  -42.1571,
  -42.165,
  -42.1734,
  -42.1821,
  -42.1906,
  -42.1987,
  -42.2059,
  -42.2124,
  -42.218,
  -42.2229,
  -42.2275,
  -42.2311,
  -42.2363,
  -42.2424,
  -42.2499,
  -42.2588,
  -42.2688,
  -42.2799,
  -42.2914,
  -42.303,
  -42.3134,
  -42.3223,
  -42.3293,
  -42.3345,
  -42.3379,
  -42.3394,
  -42.339,
  -42.337,
  -42.3331,
  -42.3281,
  -42.3224,
  -42.3165,
  -42.3108,
  -42.3054,
  -42.3001,
  -42.2952,
  -42.2902,
  -42.2853,
  -42.2806,
  -42.2757,
  -42.2709,
  -42.2645,
  -42.2557,
  -42.2437,
  -42.2279,
  -42.208,
  -42.1843,
  -42.1569,
  -42.1259,
  -42.0912,
  -42.0531,
  -42.0103,
  -41.9648,
  -41.9162,
  -41.8647,
  -41.8091,
  -41.7487,
  -41.6826,
  -41.6107,
  -41.5324,
  -41.4475,
  -41.3566,
  -41.2605,
  -41.1604,
  -41.0581,
  -40.9561,
  -40.8573,
  -40.7641,
  -40.6787,
  -37.3918,
  -37.4334,
  -37.4756,
  -37.5188,
  -37.5628,
  -37.6077,
  -37.6525,
  -37.6971,
  -37.7414,
  -37.7855,
  -37.8288,
  -37.8708,
  -37.9132,
  -37.9544,
  -37.9946,
  -38.0345,
  -38.0743,
  -38.1137,
  -38.1524,
  -38.1902,
  -38.2269,
  -38.2627,
  -38.2972,
  -38.3303,
  -38.3621,
  -38.3914,
  -38.4203,
  -38.4478,
  -38.4744,
  -38.5,
  -38.5251,
  -38.5501,
  -38.5756,
  -38.6019,
  -38.6294,
  -38.6584,
  -38.6891,
  -38.7211,
  -38.754,
  -38.7871,
  -38.8199,
  -38.8511,
  -38.8828,
  -38.914,
  -38.945,
  -38.9759,
  -39.0069,
  -39.0382,
  -39.0696,
  -39.1005,
  -39.1307,
  -39.1601,
  -39.1882,
  -39.2152,
  -39.241,
  -39.2659,
  -39.2899,
  -39.3126,
  -39.3358,
  -39.359,
  -39.3825,
  -39.4066,
  -39.4312,
  -39.4561,
  -39.4813,
  -39.507,
  -39.5334,
  -39.5609,
  -39.5898,
  -39.62,
  -39.6513,
  -39.6826,
  -39.7137,
  -39.743,
  -39.7726,
  -39.8021,
  -39.832,
  -39.8624,
  -39.8934,
  -39.9253,
  -39.9575,
  -39.9895,
  -40.0209,
  -40.0517,
  -40.0809,
  -40.1086,
  -40.135,
  -40.1613,
  -40.1874,
  -40.2138,
  -40.2414,
  -40.2692,
  -40.299,
  -40.3294,
  -40.3597,
  -40.3896,
  -40.4186,
  -40.4461,
  -40.4719,
  -40.4962,
  -40.5194,
  -40.5422,
  -40.5654,
  -40.5892,
  -40.6135,
  -40.6378,
  -40.6616,
  -40.684,
  -40.7051,
  -40.7242,
  -40.7404,
  -40.7551,
  -40.7673,
  -40.7761,
  -40.7823,
  -40.7854,
  -40.7865,
  -40.7862,
  -40.786,
  -40.7862,
  -40.7872,
  -40.7894,
  -40.7923,
  -40.7954,
  -40.799,
  -40.8023,
  -40.8062,
  -40.8098,
  -40.8137,
  -40.818,
  -40.8221,
  -40.8285,
  -40.8363,
  -40.8454,
  -40.8556,
  -40.8671,
  -40.8798,
  -40.8928,
  -40.9065,
  -40.9201,
  -40.9341,
  -40.9481,
  -40.9624,
  -40.9773,
  -40.9924,
  -41.0078,
  -41.0231,
  -41.0381,
  -41.0529,
  -41.0677,
  -41.0824,
  -41.097,
  -41.1108,
  -41.1261,
  -41.1422,
  -41.1591,
  -41.1769,
  -41.1953,
  -41.2137,
  -41.232,
  -41.2494,
  -41.2661,
  -41.2823,
  -41.2986,
  -41.3146,
  -41.3311,
  -41.3478,
  -41.3646,
  -41.3818,
  -41.399,
  -41.4165,
  -41.4342,
  -41.4527,
  -41.4721,
  -41.4923,
  -41.5122,
  -41.5342,
  -41.5566,
  -41.5783,
  -41.5994,
  -41.6189,
  -41.6372,
  -41.6543,
  -41.672,
  -41.6915,
  -41.7134,
  -41.7378,
  -41.7637,
  -41.7903,
  -41.8161,
  -41.84,
  -41.8611,
  -41.8787,
  -41.8935,
  -41.9057,
  -41.9161,
  -41.926,
  -41.9359,
  -41.946,
  -41.9561,
  -41.9656,
  -41.9732,
  -41.9803,
  -41.9853,
  -41.9881,
  -41.989,
  -41.9879,
  -41.9861,
  -41.984,
  -41.9825,
  -41.9823,
  -41.9833,
  -41.9849,
  -41.9866,
  -41.9876,
  -41.9874,
  -41.986,
  -41.9844,
  -41.983,
  -41.9822,
  -41.9829,
  -41.9856,
  -41.9908,
  -41.9985,
  -42.0086,
  -42.0205,
  -42.033,
  -42.045,
  -42.0561,
  -42.0656,
  -42.074,
  -42.0822,
  -42.0892,
  -42.0976,
  -42.1065,
  -42.1158,
  -42.1249,
  -42.1338,
  -42.142,
  -42.1493,
  -42.1557,
  -42.1612,
  -42.1661,
  -42.1708,
  -42.1759,
  -42.1821,
  -42.1899,
  -42.1992,
  -42.2099,
  -42.2217,
  -42.2344,
  -42.247,
  -42.2585,
  -42.2682,
  -42.2764,
  -42.2825,
  -42.2869,
  -42.2896,
  -42.2906,
  -42.2898,
  -42.2873,
  -42.2837,
  -42.2788,
  -42.2734,
  -42.2678,
  -42.2624,
  -42.2568,
  -42.2515,
  -42.2455,
  -42.2406,
  -42.2359,
  -42.2311,
  -42.226,
  -42.2195,
  -42.2105,
  -42.1982,
  -42.1821,
  -42.1615,
  -42.1369,
  -42.1088,
  -42.0771,
  -42.0426,
  -42.0051,
  -41.9644,
  -41.9205,
  -41.8738,
  -41.8235,
  -41.7695,
  -41.7114,
  -41.648,
  -41.5792,
  -41.5044,
  -41.4231,
  -41.3353,
  -41.2415,
  -41.1427,
  -41.0409,
  -40.9379,
  -40.8373,
  -40.7416,
  -40.6531,
  -37.2361,
  -37.2772,
  -37.3193,
  -37.3621,
  -37.4059,
  -37.4499,
  -37.4932,
  -37.5371,
  -37.5807,
  -37.6245,
  -37.6679,
  -37.7114,
  -37.754,
  -37.7962,
  -37.8374,
  -37.8781,
  -37.9183,
  -37.9579,
  -37.9967,
  -38.0343,
  -38.0697,
  -38.1053,
  -38.1397,
  -38.1731,
  -38.2053,
  -38.2359,
  -38.2651,
  -38.2932,
  -38.3202,
  -38.3467,
  -38.3723,
  -38.398,
  -38.424,
  -38.4508,
  -38.4787,
  -38.5079,
  -38.5377,
  -38.57,
  -38.6032,
  -38.6369,
  -38.6706,
  -38.704,
  -38.7371,
  -38.7699,
  -38.8025,
  -38.8349,
  -38.8673,
  -38.8998,
  -38.932,
  -38.9635,
  -38.9942,
  -39.023,
  -39.0518,
  -39.08,
  -39.1069,
  -39.1329,
  -39.1578,
  -39.182,
  -39.2057,
  -39.2294,
  -39.2533,
  -39.2779,
  -39.303,
  -39.3285,
  -39.3543,
  -39.3806,
  -39.4076,
  -39.4361,
  -39.4652,
  -39.4967,
  -39.5291,
  -39.5615,
  -39.5933,
  -39.6243,
  -39.6549,
  -39.6853,
  -39.7162,
  -39.7476,
  -39.7793,
  -39.8117,
  -39.8443,
  -39.8771,
  -39.9094,
  -39.9401,
  -39.9691,
  -39.9956,
  -40.022,
  -40.048,
  -40.0744,
  -40.1016,
  -40.1302,
  -40.1599,
  -40.1906,
  -40.2217,
  -40.2527,
  -40.2831,
  -40.3126,
  -40.3408,
  -40.3669,
  -40.3915,
  -40.415,
  -40.438,
  -40.4611,
  -40.4846,
  -40.5076,
  -40.532,
  -40.5559,
  -40.5789,
  -40.6003,
  -40.62,
  -40.6379,
  -40.6536,
  -40.6666,
  -40.6765,
  -40.683,
  -40.6866,
  -40.6876,
  -40.687,
  -40.6866,
  -40.6863,
  -40.6869,
  -40.6888,
  -40.6914,
  -40.6942,
  -40.6986,
  -40.7032,
  -40.7079,
  -40.7127,
  -40.7173,
  -40.722,
  -40.7274,
  -40.7335,
  -40.7406,
  -40.7492,
  -40.7591,
  -40.7705,
  -40.7831,
  -40.7966,
  -40.8106,
  -40.8247,
  -40.8391,
  -40.8538,
  -40.869,
  -40.8845,
  -40.8994,
  -40.9155,
  -40.9313,
  -40.9468,
  -40.9622,
  -40.9777,
  -40.9931,
  -41.0085,
  -41.024,
  -41.0402,
  -41.0569,
  -41.0745,
  -41.0923,
  -41.1106,
  -41.1287,
  -41.1468,
  -41.1642,
  -41.1811,
  -41.1976,
  -41.214,
  -41.2301,
  -41.2461,
  -41.2622,
  -41.2772,
  -41.2934,
  -41.3095,
  -41.326,
  -41.3433,
  -41.3612,
  -41.3802,
  -41.4007,
  -41.4224,
  -41.445,
  -41.4676,
  -41.4898,
  -41.5105,
  -41.5298,
  -41.5476,
  -41.5648,
  -41.5829,
  -41.6034,
  -41.6261,
  -41.6511,
  -41.678,
  -41.7055,
  -41.7325,
  -41.7573,
  -41.7793,
  -41.797,
  -41.8123,
  -41.825,
  -41.8358,
  -41.8456,
  -41.8554,
  -41.8654,
  -41.8757,
  -41.8854,
  -41.8941,
  -41.9012,
  -41.9063,
  -41.9092,
  -41.9099,
  -41.9091,
  -41.9073,
  -41.9056,
  -41.9047,
  -41.9049,
  -41.9064,
  -41.909,
  -41.9117,
  -41.914,
  -41.9151,
  -41.915,
  -41.9142,
  -41.9138,
  -41.9141,
  -41.9159,
  -41.9186,
  -41.9247,
  -41.9331,
  -41.9439,
  -41.9557,
  -41.9678,
  -41.979,
  -41.989,
  -41.9975,
  -42.0055,
  -42.0133,
  -42.0211,
  -42.0297,
  -42.039,
  -42.0487,
  -42.0586,
  -42.0683,
  -42.0774,
  -42.0858,
  -42.0934,
  -42.0999,
  -42.1055,
  -42.1106,
  -42.1159,
  -42.1225,
  -42.1305,
  -42.1403,
  -42.1517,
  -42.1645,
  -42.1777,
  -42.1909,
  -42.203,
  -42.2134,
  -42.2223,
  -42.2286,
  -42.2343,
  -42.2383,
  -42.2407,
  -42.2412,
  -42.2402,
  -42.2377,
  -42.2338,
  -42.2289,
  -42.2234,
  -42.2177,
  -42.2121,
  -42.2064,
  -42.2012,
  -42.196,
  -42.1909,
  -42.1859,
  -42.1804,
  -42.1737,
  -42.1645,
  -42.1521,
  -42.1356,
  -42.1147,
  -42.0893,
  -42.0607,
  -42.0287,
  -41.9941,
  -41.9572,
  -41.9176,
  -41.8756,
  -41.83,
  -41.7815,
  -41.729,
  -41.6724,
  -41.6111,
  -41.5451,
  -41.4734,
  -41.3954,
  -41.3105,
  -41.219,
  -41.1221,
  -41.0211,
  -40.9184,
  -40.8165,
  -40.7178,
  -40.6265,
  -37.0816,
  -37.1213,
  -37.1629,
  -37.2054,
  -37.2485,
  -37.292,
  -37.3354,
  -37.3786,
  -37.4218,
  -37.4651,
  -37.5086,
  -37.5524,
  -37.5957,
  -37.6386,
  -37.6807,
  -37.7223,
  -37.7621,
  -37.8019,
  -37.8404,
  -37.8777,
  -37.9139,
  -37.9489,
  -37.9833,
  -38.0168,
  -38.0494,
  -38.0806,
  -38.1104,
  -38.139,
  -38.1667,
  -38.1935,
  -38.219,
  -38.2455,
  -38.2722,
  -38.2995,
  -38.3278,
  -38.3572,
  -38.3882,
  -38.4205,
  -38.454,
  -38.4883,
  -38.5228,
  -38.5573,
  -38.5917,
  -38.626,
  -38.6601,
  -38.6941,
  -38.7269,
  -38.7603,
  -38.7933,
  -38.8254,
  -38.8566,
  -38.8871,
  -38.917,
  -38.9462,
  -38.9743,
  -39.0012,
  -39.027,
  -39.0519,
  -39.0761,
  -39.1004,
  -39.1248,
  -39.1498,
  -39.1745,
  -39.2006,
  -39.2271,
  -39.2539,
  -39.2817,
  -39.311,
  -39.3422,
  -39.375,
  -39.4084,
  -39.4416,
  -39.4741,
  -39.5058,
  -39.5373,
  -39.5689,
  -39.6008,
  -39.6329,
  -39.6651,
  -39.6968,
  -39.7301,
  -39.7631,
  -39.7956,
  -39.8267,
  -39.8559,
  -39.8833,
  -39.9097,
  -39.9358,
  -39.9627,
  -39.9909,
  -40.0203,
  -40.051,
  -40.0823,
  -40.1138,
  -40.1454,
  -40.1764,
  -40.2061,
  -40.2337,
  -40.2608,
  -40.2861,
  -40.3098,
  -40.3333,
  -40.3568,
  -40.3806,
  -40.405,
  -40.4295,
  -40.4536,
  -40.4765,
  -40.4979,
  -40.5177,
  -40.5359,
  -40.5517,
  -40.5652,
  -40.5757,
  -40.583,
  -40.5869,
  -40.5886,
  -40.5876,
  -40.5868,
  -40.5865,
  -40.5869,
  -40.5886,
  -40.5912,
  -40.5951,
  -40.6,
  -40.6054,
  -40.6113,
  -40.6171,
  -40.6227,
  -40.6279,
  -40.6334,
  -40.6395,
  -40.6463,
  -40.6543,
  -40.6637,
  -40.6749,
  -40.6873,
  -40.6997,
  -40.714,
  -40.7286,
  -40.7441,
  -40.7598,
  -40.776,
  -40.7923,
  -40.8088,
  -40.8254,
  -40.8416,
  -40.8577,
  -40.8737,
  -40.8898,
  -40.9062,
  -40.9226,
  -40.9395,
  -40.9567,
  -40.974,
  -40.9915,
  -41.0093,
  -41.0271,
  -41.0448,
  -41.0613,
  -41.0785,
  -41.0956,
  -41.1125,
  -41.1289,
  -41.1449,
  -41.1609,
  -41.1766,
  -41.1919,
  -41.207,
  -41.2221,
  -41.238,
  -41.2548,
  -41.2726,
  -41.2915,
  -41.3119,
  -41.3336,
  -41.3561,
  -41.3785,
  -41.4004,
  -41.421,
  -41.4397,
  -41.4574,
  -41.4752,
  -41.4937,
  -41.5137,
  -41.537,
  -41.5628,
  -41.5907,
  -41.619,
  -41.647,
  -41.673,
  -41.6963,
  -41.7161,
  -41.7322,
  -41.7452,
  -41.7561,
  -41.7663,
  -41.7762,
  -41.7861,
  -41.796,
  -41.806,
  -41.8146,
  -41.822,
  -41.8271,
  -41.8298,
  -41.8308,
  -41.83,
  -41.8286,
  -41.8274,
  -41.8269,
  -41.8277,
  -41.8288,
  -41.8321,
  -41.8356,
  -41.8388,
  -41.841,
  -41.8418,
  -41.8421,
  -41.8426,
  -41.844,
  -41.8468,
  -41.8516,
  -41.8586,
  -41.868,
  -41.8792,
  -41.8911,
  -41.9027,
  -41.9131,
  -41.9221,
  -41.9299,
  -41.9371,
  -41.9444,
  -41.9521,
  -41.9605,
  -41.97,
  -41.9802,
  -41.9908,
  -42.0014,
  -42.0116,
  -42.0213,
  -42.0302,
  -42.0378,
  -42.0444,
  -42.0492,
  -42.0551,
  -42.0622,
  -42.0708,
  -42.0813,
  -42.0935,
  -42.1068,
  -42.1205,
  -42.1336,
  -42.1459,
  -42.1567,
  -42.1663,
  -42.1746,
  -42.1816,
  -42.1869,
  -42.1905,
  -42.1924,
  -42.1928,
  -42.1916,
  -42.1887,
  -42.1844,
  -42.1791,
  -42.1734,
  -42.1677,
  -42.162,
  -42.1562,
  -42.1506,
  -42.1451,
  -42.1397,
  -42.1336,
  -42.1265,
  -42.1169,
  -42.1042,
  -42.0875,
  -42.0663,
  -42.0408,
  -42.0116,
  -41.9795,
  -41.9453,
  -41.9089,
  -41.8697,
  -41.8289,
  -41.7848,
  -41.7374,
  -41.6862,
  -41.631,
  -41.5716,
  -41.5078,
  -41.4385,
  -41.3633,
  -41.2813,
  -41.1924,
  -41.0977,
  -40.9983,
  -40.8961,
  -40.7939,
  -40.6945,
  -40.6007,
  -36.9273,
  -36.9678,
  -37.0088,
  -37.0507,
  -37.0932,
  -37.136,
  -37.1787,
  -37.2213,
  -37.2641,
  -37.3071,
  -37.3506,
  -37.3934,
  -37.4373,
  -37.4809,
  -37.5238,
  -37.5659,
  -37.607,
  -37.647,
  -37.6856,
  -37.7226,
  -37.7584,
  -37.7933,
  -37.8275,
  -37.8611,
  -37.8938,
  -37.9244,
  -37.9547,
  -37.9839,
  -38.0123,
  -38.0401,
  -38.0675,
  -38.0949,
  -38.1225,
  -38.1505,
  -38.1792,
  -38.2091,
  -38.2403,
  -38.2728,
  -38.3065,
  -38.3412,
  -38.3763,
  -38.4108,
  -38.4463,
  -38.4819,
  -38.5173,
  -38.5527,
  -38.5876,
  -38.622,
  -38.6557,
  -38.6885,
  -38.7203,
  -38.7516,
  -38.7824,
  -38.8125,
  -38.8418,
  -38.8698,
  -38.8965,
  -38.9211,
  -38.9461,
  -38.9708,
  -38.9959,
  -39.0216,
  -39.0476,
  -39.0745,
  -39.1015,
  -39.129,
  -39.1576,
  -39.1878,
  -39.2199,
  -39.2536,
  -39.2881,
  -39.3221,
  -39.3556,
  -39.3884,
  -39.4197,
  -39.452,
  -39.4845,
  -39.517,
  -39.5497,
  -39.5826,
  -39.6159,
  -39.6494,
  -39.682,
  -39.7133,
  -39.7431,
  -39.7711,
  -39.7979,
  -39.8247,
  -39.8521,
  -39.8811,
  -39.9112,
  -39.9415,
  -39.9735,
  -40.0051,
  -40.0369,
  -40.0683,
  -40.0987,
  -40.1279,
  -40.1557,
  -40.1818,
  -40.2065,
  -40.2305,
  -40.2543,
  -40.2786,
  -40.3034,
  -40.3282,
  -40.3526,
  -40.3756,
  -40.397,
  -40.4166,
  -40.4335,
  -40.4495,
  -40.4628,
  -40.4734,
  -40.4809,
  -40.4856,
  -40.4878,
  -40.4886,
  -40.4885,
  -40.4886,
  -40.4891,
  -40.4907,
  -40.4934,
  -40.4974,
  -40.5027,
  -40.5086,
  -40.5153,
  -40.5221,
  -40.5284,
  -40.5343,
  -40.5392,
  -40.5453,
  -40.552,
  -40.5597,
  -40.5688,
  -40.5795,
  -40.5917,
  -40.6052,
  -40.6197,
  -40.635,
  -40.6511,
  -40.6678,
  -40.6851,
  -40.7024,
  -40.7197,
  -40.7368,
  -40.7535,
  -40.77,
  -40.7864,
  -40.803,
  -40.82,
  -40.8377,
  -40.8545,
  -40.8726,
  -40.8909,
  -40.9089,
  -40.9267,
  -40.944,
  -40.9609,
  -40.9779,
  -40.9948,
  -41.0118,
  -41.0289,
  -41.0454,
  -41.0612,
  -41.077,
  -41.0924,
  -41.1072,
  -41.1218,
  -41.1364,
  -41.1519,
  -41.168,
  -41.1853,
  -41.2041,
  -41.2243,
  -41.2449,
  -41.267,
  -41.2891,
  -41.3105,
  -41.3306,
  -41.349,
  -41.3666,
  -41.3846,
  -41.4035,
  -41.4246,
  -41.4486,
  -41.4749,
  -41.5033,
  -41.5327,
  -41.5616,
  -41.5887,
  -41.613,
  -41.6336,
  -41.6503,
  -41.664,
  -41.6757,
  -41.6863,
  -41.6964,
  -41.7066,
  -41.7169,
  -41.7269,
  -41.7359,
  -41.7422,
  -41.7472,
  -41.7498,
  -41.7508,
  -41.7507,
  -41.7495,
  -41.7487,
  -41.7488,
  -41.7501,
  -41.7526,
  -41.7563,
  -41.7605,
  -41.7641,
  -41.7669,
  -41.7685,
  -41.7698,
  -41.7711,
  -41.7732,
  -41.7773,
  -41.7834,
  -41.7915,
  -41.8016,
  -41.8133,
  -41.825,
  -41.8359,
  -41.8455,
  -41.8541,
  -41.8614,
  -41.8681,
  -41.8749,
  -41.8813,
  -41.8899,
  -41.8995,
  -41.9102,
  -41.9213,
  -41.9327,
  -41.944,
  -41.9549,
  -41.9651,
  -41.9742,
  -41.9819,
  -41.9888,
  -41.9956,
  -42.0035,
  -42.0129,
  -42.024,
  -42.0367,
  -42.0503,
  -42.064,
  -42.0772,
  -42.0895,
  -42.1006,
  -42.1109,
  -42.1202,
  -42.1281,
  -42.1345,
  -42.1393,
  -42.1425,
  -42.1441,
  -42.1441,
  -42.1423,
  -42.1387,
  -42.1339,
  -42.1284,
  -42.1227,
  -42.117,
  -42.1101,
  -42.1043,
  -42.0983,
  -42.0922,
  -42.0855,
  -42.0776,
  -42.0678,
  -42.0547,
  -42.0376,
  -42.0161,
  -41.9903,
  -41.9611,
  -41.9291,
  -41.8951,
  -41.8595,
  -41.8224,
  -41.7829,
  -41.7403,
  -41.6941,
  -41.6442,
  -41.5902,
  -41.5321,
  -41.4699,
  -41.4027,
  -41.3298,
  -41.2504,
  -41.1638,
  -41.0714,
  -40.9738,
  -40.8729,
  -40.7708,
  -40.6703,
  -40.5744,
  -36.7753,
  -36.8153,
  -36.8559,
  -36.8973,
  -36.9391,
  -36.9812,
  -37.0223,
  -37.0644,
  -37.1069,
  -37.1498,
  -37.1933,
  -37.2372,
  -37.2814,
  -37.3253,
  -37.3686,
  -37.411,
  -37.4524,
  -37.4925,
  -37.5311,
  -37.5681,
  -37.6036,
  -37.6374,
  -37.6716,
  -37.7053,
  -37.7382,
  -37.7701,
  -37.8009,
  -37.8306,
  -37.8598,
  -37.8886,
  -37.9171,
  -37.9455,
  -37.9741,
  -38.003,
  -38.0326,
  -38.0631,
  -38.0937,
  -38.1265,
  -38.1605,
  -38.1955,
  -38.2311,
  -38.2673,
  -38.3039,
  -38.3406,
  -38.3772,
  -38.4135,
  -38.4493,
  -38.4844,
  -38.5186,
  -38.5519,
  -38.5846,
  -38.6157,
  -38.6473,
  -38.6783,
  -38.7086,
  -38.7376,
  -38.7652,
  -38.7917,
  -38.8174,
  -38.8429,
  -38.8685,
  -38.8947,
  -38.9212,
  -38.9485,
  -38.9765,
  -39.0048,
  -39.0342,
  -39.0654,
  -39.0973,
  -39.1318,
  -39.1671,
  -39.2024,
  -39.2369,
  -39.2706,
  -39.3038,
  -39.3368,
  -39.3695,
  -39.4022,
  -39.435,
  -39.468,
  -39.5015,
  -39.5352,
  -39.5683,
  -39.6003,
  -39.6306,
  -39.6583,
  -39.6859,
  -39.7137,
  -39.7416,
  -39.7708,
  -39.8016,
  -39.8332,
  -39.8654,
  -39.8975,
  -39.9296,
  -39.9614,
  -39.9924,
  -40.0226,
  -40.0511,
  -40.078,
  -40.1037,
  -40.1287,
  -40.1532,
  -40.1781,
  -40.2022,
  -40.2272,
  -40.2515,
  -40.2745,
  -40.2959,
  -40.3154,
  -40.3332,
  -40.3488,
  -40.3617,
  -40.3722,
  -40.3799,
  -40.385,
  -40.3879,
  -40.3896,
  -40.3905,
  -40.3911,
  -40.3923,
  -40.394,
  -40.3971,
  -40.4005,
  -40.4061,
  -40.4126,
  -40.4198,
  -40.4272,
  -40.434,
  -40.4402,
  -40.4466,
  -40.453,
  -40.4599,
  -40.4675,
  -40.4765,
  -40.4868,
  -40.4985,
  -40.5118,
  -40.5263,
  -40.5422,
  -40.559,
  -40.5767,
  -40.5949,
  -40.6132,
  -40.6304,
  -40.6481,
  -40.6655,
  -40.6825,
  -40.6994,
  -40.7165,
  -40.7339,
  -40.7521,
  -40.7707,
  -40.7899,
  -40.8091,
  -40.8275,
  -40.8451,
  -40.8621,
  -40.8788,
  -40.8954,
  -40.9121,
  -40.929,
  -40.9458,
  -40.9622,
  -40.9778,
  -40.9931,
  -41.0082,
  -41.0217,
  -41.0361,
  -41.0502,
  -41.0652,
  -41.0812,
  -41.0983,
  -41.1166,
  -41.1365,
  -41.1577,
  -41.1793,
  -41.2012,
  -41.2223,
  -41.2422,
  -41.2604,
  -41.278,
  -41.2958,
  -41.315,
  -41.3364,
  -41.3607,
  -41.3876,
  -41.4162,
  -41.4461,
  -41.4757,
  -41.5035,
  -41.5287,
  -41.5505,
  -41.5672,
  -41.5819,
  -41.5944,
  -41.6057,
  -41.6167,
  -41.6277,
  -41.6384,
  -41.6486,
  -41.6576,
  -41.6645,
  -41.6694,
  -41.6719,
  -41.6725,
  -41.6725,
  -41.6718,
  -41.6714,
  -41.6721,
  -41.6739,
  -41.677,
  -41.6808,
  -41.685,
  -41.6888,
  -41.6921,
  -41.6945,
  -41.6963,
  -41.6983,
  -41.7014,
  -41.7061,
  -41.7121,
  -41.7214,
  -41.7321,
  -41.7437,
  -41.7551,
  -41.7659,
  -41.7758,
  -41.7841,
  -41.7911,
  -41.7976,
  -41.8042,
  -41.8117,
  -41.8203,
  -41.8303,
  -41.8414,
  -41.8532,
  -41.8653,
  -41.8773,
  -41.8893,
  -41.9006,
  -41.9109,
  -41.9198,
  -41.9281,
  -41.9362,
  -41.945,
  -41.9552,
  -41.9669,
  -41.9799,
  -41.9935,
  -42.0071,
  -42.0203,
  -42.0325,
  -42.0441,
  -42.055,
  -42.0641,
  -42.0729,
  -42.0803,
  -42.0861,
  -42.0903,
  -42.093,
  -42.0941,
  -42.0932,
  -42.0906,
  -42.0864,
  -42.0814,
  -42.0761,
  -42.0707,
  -42.0651,
  -42.0592,
  -42.0528,
  -42.046,
  -42.0387,
  -42.0302,
  -42.0197,
  -42.0058,
  -41.9882,
  -41.9665,
  -41.9406,
  -41.9113,
  -41.8796,
  -41.8461,
  -41.8114,
  -41.7754,
  -41.7373,
  -41.6962,
  -41.6511,
  -41.6021,
  -41.5491,
  -41.4923,
  -41.4312,
  -41.3655,
  -41.2943,
  -41.2169,
  -41.1325,
  -41.0421,
  -40.9465,
  -40.8468,
  -40.7452,
  -40.6441,
  -40.5452,
  -36.6245,
  -36.663,
  -36.7031,
  -36.7438,
  -36.7851,
  -36.8266,
  -36.8683,
  -36.9104,
  -36.9528,
  -36.9958,
  -37.0393,
  -37.0834,
  -37.1276,
  -37.1716,
  -37.2148,
  -37.2572,
  -37.2975,
  -37.3375,
  -37.3761,
  -37.4131,
  -37.4487,
  -37.4835,
  -37.5178,
  -37.5516,
  -37.5848,
  -37.617,
  -37.6483,
  -37.6787,
  -37.7089,
  -37.7386,
  -37.7684,
  -37.797,
  -37.8267,
  -37.8568,
  -37.8874,
  -37.9188,
  -37.9511,
  -37.9843,
  -38.0185,
  -38.0538,
  -38.0898,
  -38.1266,
  -38.1639,
  -38.2015,
  -38.239,
  -38.2761,
  -38.3113,
  -38.3468,
  -38.3814,
  -38.4153,
  -38.4485,
  -38.4815,
  -38.5139,
  -38.5457,
  -38.5766,
  -38.6064,
  -38.6349,
  -38.6624,
  -38.689,
  -38.7153,
  -38.7417,
  -38.7683,
  -38.7946,
  -38.8225,
  -38.8511,
  -38.8804,
  -38.9109,
  -38.9428,
  -38.9765,
  -39.0118,
  -39.0479,
  -39.0841,
  -39.1198,
  -39.1547,
  -39.1889,
  -39.2224,
  -39.2554,
  -39.288,
  -39.3206,
  -39.3534,
  -39.386,
  -39.4198,
  -39.4535,
  -39.4866,
  -39.5181,
  -39.548,
  -39.5763,
  -39.6047,
  -39.6333,
  -39.6627,
  -39.6938,
  -39.7253,
  -39.7573,
  -39.7897,
  -39.8221,
  -39.8544,
  -39.8863,
  -39.9172,
  -39.9457,
  -39.9736,
  -40.0003,
  -40.0262,
  -40.0518,
  -40.0774,
  -40.1031,
  -40.1282,
  -40.1526,
  -40.1753,
  -40.1965,
  -40.2158,
  -40.2334,
  -40.2484,
  -40.2612,
  -40.2713,
  -40.2792,
  -40.285,
  -40.2891,
  -40.291,
  -40.2926,
  -40.2938,
  -40.2955,
  -40.298,
  -40.3017,
  -40.3066,
  -40.3126,
  -40.3197,
  -40.3273,
  -40.3349,
  -40.3418,
  -40.3482,
  -40.3549,
  -40.3614,
  -40.3685,
  -40.3764,
  -40.3856,
  -40.3961,
  -40.4076,
  -40.4196,
  -40.4339,
  -40.4499,
  -40.467,
  -40.4854,
  -40.5044,
  -40.5235,
  -40.5425,
  -40.5611,
  -40.5791,
  -40.5967,
  -40.6141,
  -40.6316,
  -40.6496,
  -40.6682,
  -40.6875,
  -40.7073,
  -40.727,
  -40.7458,
  -40.7637,
  -40.7807,
  -40.7972,
  -40.8126,
  -40.829,
  -40.8454,
  -40.8616,
  -40.8775,
  -40.8929,
  -40.9082,
  -40.923,
  -40.9374,
  -40.9515,
  -40.9656,
  -40.9803,
  -40.996,
  -41.0129,
  -41.0311,
  -41.0504,
  -41.0709,
  -41.0919,
  -41.1131,
  -41.1337,
  -41.1528,
  -41.171,
  -41.189,
  -41.2071,
  -41.2266,
  -41.2476,
  -41.2721,
  -41.2992,
  -41.3283,
  -41.3584,
  -41.3882,
  -41.4169,
  -41.443,
  -41.4657,
  -41.4847,
  -41.5006,
  -41.5143,
  -41.5269,
  -41.5391,
  -41.5508,
  -41.562,
  -41.572,
  -41.581,
  -41.5879,
  -41.5924,
  -41.5947,
  -41.5952,
  -41.5947,
  -41.5945,
  -41.5948,
  -41.5961,
  -41.5984,
  -41.6004,
  -41.6044,
  -41.6085,
  -41.6128,
  -41.6164,
  -41.6191,
  -41.6214,
  -41.624,
  -41.6276,
  -41.6332,
  -41.6408,
  -41.6504,
  -41.6614,
  -41.6731,
  -41.6849,
  -41.6959,
  -41.7056,
  -41.7139,
  -41.7212,
  -41.728,
  -41.7349,
  -41.7428,
  -41.752,
  -41.7623,
  -41.774,
  -41.7861,
  -41.7988,
  -41.8118,
  -41.8242,
  -41.8363,
  -41.8474,
  -41.8576,
  -41.8661,
  -41.8757,
  -41.8855,
  -41.8963,
  -41.9084,
  -41.9214,
  -41.935,
  -41.9485,
  -41.9617,
  -41.9742,
  -41.9863,
  -41.9979,
  -42.0087,
  -42.0181,
  -42.0265,
  -42.033,
  -42.0378,
  -42.0412,
  -42.0431,
  -42.0433,
  -42.0419,
  -42.0389,
  -42.0348,
  -42.0302,
  -42.0252,
  -42.0201,
  -42.0144,
  -42.0079,
  -42.0009,
  -41.9927,
  -41.9834,
  -41.9719,
  -41.9575,
  -41.9392,
  -41.9169,
  -41.891,
  -41.8617,
  -41.8304,
  -41.7976,
  -41.7639,
  -41.7281,
  -41.6916,
  -41.6518,
  -41.6079,
  -41.5596,
  -41.5074,
  -41.4514,
  -41.3914,
  -41.3267,
  -41.2567,
  -41.1805,
  -41.0978,
  -41.0091,
  -40.9148,
  -40.8163,
  -40.7149,
  -40.613,
  -40.5136,
  -36.4744,
  -36.5134,
  -36.5529,
  -36.5932,
  -36.6341,
  -36.6753,
  -36.7168,
  -36.7587,
  -36.8011,
  -36.8442,
  -36.888,
  -36.9312,
  -36.9753,
  -37.019,
  -37.0619,
  -37.1039,
  -37.1449,
  -37.1849,
  -37.2234,
  -37.2604,
  -37.296,
  -37.3308,
  -37.3652,
  -37.3994,
  -37.4329,
  -37.4655,
  -37.4964,
  -37.5278,
  -37.559,
  -37.59,
  -37.6208,
  -37.6515,
  -37.6824,
  -37.7138,
  -37.7456,
  -37.778,
  -37.811,
  -37.8448,
  -37.8793,
  -37.9146,
  -37.9509,
  -37.9871,
  -38.0251,
  -38.0634,
  -38.1015,
  -38.139,
  -38.1757,
  -38.2116,
  -38.2466,
  -38.2809,
  -38.3147,
  -38.3481,
  -38.381,
  -38.4133,
  -38.4448,
  -38.4753,
  -38.5047,
  -38.5321,
  -38.5598,
  -38.5872,
  -38.6145,
  -38.6419,
  -38.67,
  -38.6987,
  -38.728,
  -38.7583,
  -38.7896,
  -38.8224,
  -38.857,
  -38.8931,
  -38.93,
  -38.967,
  -39.0038,
  -39.0398,
  -39.0738,
  -39.108,
  -39.1412,
  -39.1739,
  -39.2063,
  -39.2392,
  -39.2725,
  -39.3066,
  -39.3405,
  -39.3742,
  -39.4067,
  -39.4379,
  -39.4674,
  -39.4961,
  -39.5249,
  -39.5544,
  -39.5852,
  -39.6169,
  -39.6481,
  -39.6806,
  -39.7133,
  -39.7462,
  -39.7788,
  -39.8106,
  -39.8407,
  -39.8698,
  -39.8976,
  -39.9244,
  -39.9511,
  -39.9778,
  -40.0039,
  -40.0294,
  -40.0534,
  -40.0761,
  -40.0969,
  -40.1157,
  -40.1319,
  -40.1467,
  -40.1592,
  -40.1695,
  -40.178,
  -40.1847,
  -40.1901,
  -40.1941,
  -40.1971,
  -40.1994,
  -40.2019,
  -40.2047,
  -40.2089,
  -40.2144,
  -40.2209,
  -40.2282,
  -40.236,
  -40.2438,
  -40.251,
  -40.2578,
  -40.2633,
  -40.2703,
  -40.2778,
  -40.286,
  -40.2955,
  -40.306,
  -40.3179,
  -40.3309,
  -40.3454,
  -40.3615,
  -40.3787,
  -40.3971,
  -40.4164,
  -40.4361,
  -40.4556,
  -40.4748,
  -40.4935,
  -40.5118,
  -40.5298,
  -40.5478,
  -40.5661,
  -40.5851,
  -40.6037,
  -40.6238,
  -40.6438,
  -40.6629,
  -40.6809,
  -40.6979,
  -40.7143,
  -40.7304,
  -40.7466,
  -40.7625,
  -40.7782,
  -40.7937,
  -40.8088,
  -40.824,
  -40.8388,
  -40.8533,
  -40.8675,
  -40.882,
  -40.897,
  -40.9125,
  -40.929,
  -40.9464,
  -40.965,
  -40.9834,
  -41.0034,
  -41.0236,
  -41.0437,
  -41.0628,
  -41.0812,
  -41.0994,
  -41.118,
  -41.1378,
  -41.16,
  -41.1848,
  -41.2122,
  -41.2416,
  -41.272,
  -41.3023,
  -41.3314,
  -41.3581,
  -41.3817,
  -41.4017,
  -41.4189,
  -41.4343,
  -41.4484,
  -41.4618,
  -41.4746,
  -41.4863,
  -41.4967,
  -41.5054,
  -41.5111,
  -41.5153,
  -41.5172,
  -41.5174,
  -41.5171,
  -41.5171,
  -41.5179,
  -41.5197,
  -41.5222,
  -41.5255,
  -41.5296,
  -41.5338,
  -41.538,
  -41.5417,
  -41.5446,
  -41.5473,
  -41.5505,
  -41.5548,
  -41.5608,
  -41.5686,
  -41.5785,
  -41.5899,
  -41.6018,
  -41.6135,
  -41.6246,
  -41.6344,
  -41.6431,
  -41.651,
  -41.6584,
  -41.6662,
  -41.6739,
  -41.6837,
  -41.6948,
  -41.7068,
  -41.7195,
  -41.7326,
  -41.7459,
  -41.7588,
  -41.7714,
  -41.7832,
  -41.7945,
  -41.8053,
  -41.816,
  -41.8269,
  -41.8384,
  -41.8506,
  -41.8638,
  -41.8772,
  -41.8906,
  -41.9037,
  -41.9164,
  -41.9291,
  -41.9415,
  -41.9529,
  -41.9631,
  -41.9719,
  -41.9789,
  -41.984,
  -41.9878,
  -41.9901,
  -41.9915,
  -41.9914,
  -41.9899,
  -41.9871,
  -41.9835,
  -41.9794,
  -41.9747,
  -41.9683,
  -41.9619,
  -41.9544,
  -41.9457,
  -41.9354,
  -41.9232,
  -41.9081,
  -41.8895,
  -41.867,
  -41.8408,
  -41.8118,
  -41.781,
  -41.7491,
  -41.7165,
  -41.6831,
  -41.6477,
  -41.6093,
  -41.5667,
  -41.5191,
  -41.4672,
  -41.4118,
  -41.3525,
  -41.2886,
  -41.2194,
  -41.1442,
  -41.0626,
  -40.9748,
  -40.8812,
  -40.7829,
  -40.6814,
  -40.5784,
  -40.477,
  -36.3268,
  -36.3652,
  -36.4043,
  -36.4442,
  -36.4848,
  -36.5259,
  -36.5665,
  -36.6087,
  -36.6514,
  -36.6947,
  -36.7386,
  -36.7829,
  -36.8268,
  -36.8699,
  -36.9122,
  -36.9538,
  -36.9942,
  -37.0338,
  -37.0722,
  -37.1092,
  -37.1449,
  -37.1787,
  -37.2134,
  -37.2478,
  -37.2819,
  -37.3153,
  -37.3482,
  -37.3805,
  -37.4128,
  -37.4447,
  -37.4765,
  -37.5083,
  -37.5404,
  -37.5728,
  -37.6058,
  -37.6392,
  -37.672,
  -37.7062,
  -37.7409,
  -37.7765,
  -37.8131,
  -37.8507,
  -37.8891,
  -37.9279,
  -37.9664,
  -38.0042,
  -38.0412,
  -38.0774,
  -38.1128,
  -38.1475,
  -38.1817,
  -38.2154,
  -38.2476,
  -38.2802,
  -38.3122,
  -38.3433,
  -38.3734,
  -38.4029,
  -38.4318,
  -38.4604,
  -38.4889,
  -38.5175,
  -38.5465,
  -38.576,
  -38.6061,
  -38.6372,
  -38.6696,
  -38.7034,
  -38.7379,
  -38.7749,
  -38.8126,
  -38.8506,
  -38.8882,
  -38.925,
  -38.9609,
  -38.9955,
  -39.0291,
  -39.0621,
  -39.0946,
  -39.1274,
  -39.1608,
  -39.1948,
  -39.2291,
  -39.2632,
  -39.2963,
  -39.3279,
  -39.3571,
  -39.3864,
  -39.4156,
  -39.4452,
  -39.4759,
  -39.5074,
  -39.5396,
  -39.5723,
  -39.6055,
  -39.6389,
  -39.6717,
  -39.7042,
  -39.7352,
  -39.7653,
  -39.7939,
  -39.8225,
  -39.8503,
  -39.8777,
  -39.9034,
  -39.9289,
  -39.953,
  -39.9753,
  -39.9956,
  -40.0141,
  -40.0306,
  -40.045,
  -40.0574,
  -40.0682,
  -40.0774,
  -40.0853,
  -40.0924,
  -40.0984,
  -40.1029,
  -40.1065,
  -40.1098,
  -40.1136,
  -40.1184,
  -40.124,
  -40.1296,
  -40.1371,
  -40.1451,
  -40.153,
  -40.1604,
  -40.1675,
  -40.1747,
  -40.1821,
  -40.1901,
  -40.1989,
  -40.2085,
  -40.2191,
  -40.2311,
  -40.2442,
  -40.2589,
  -40.2749,
  -40.2923,
  -40.311,
  -40.3305,
  -40.3505,
  -40.3706,
  -40.3893,
  -40.4084,
  -40.4273,
  -40.4457,
  -40.4637,
  -40.4821,
  -40.5014,
  -40.521,
  -40.5412,
  -40.5611,
  -40.5804,
  -40.5986,
  -40.6157,
  -40.6321,
  -40.6482,
  -40.6638,
  -40.6793,
  -40.6946,
  -40.7097,
  -40.7246,
  -40.7397,
  -40.7546,
  -40.7687,
  -40.7836,
  -40.7986,
  -40.8137,
  -40.8294,
  -40.8454,
  -40.8617,
  -40.879,
  -40.8973,
  -40.9164,
  -40.9357,
  -40.9552,
  -40.9744,
  -40.993,
  -41.0115,
  -41.0306,
  -41.0512,
  -41.0738,
  -41.0992,
  -41.127,
  -41.1568,
  -41.1874,
  -41.2178,
  -41.2471,
  -41.2743,
  -41.2985,
  -41.3186,
  -41.3372,
  -41.354,
  -41.3696,
  -41.3846,
  -41.3985,
  -41.411,
  -41.4217,
  -41.4305,
  -41.4369,
  -41.4408,
  -41.4423,
  -41.4422,
  -41.4419,
  -41.4419,
  -41.4428,
  -41.445,
  -41.4478,
  -41.4513,
  -41.4551,
  -41.4594,
  -41.4634,
  -41.467,
  -41.4703,
  -41.4733,
  -41.4769,
  -41.4816,
  -41.4879,
  -41.4964,
  -41.5057,
  -41.5173,
  -41.5293,
  -41.5409,
  -41.5518,
  -41.5619,
  -41.571,
  -41.5796,
  -41.5882,
  -41.5972,
  -41.607,
  -41.6178,
  -41.6295,
  -41.642,
  -41.655,
  -41.6683,
  -41.6818,
  -41.6952,
  -41.7082,
  -41.7209,
  -41.7331,
  -41.745,
  -41.7566,
  -41.7684,
  -41.7803,
  -41.7928,
  -41.8057,
  -41.8189,
  -41.8324,
  -41.8457,
  -41.8589,
  -41.8722,
  -41.8851,
  -41.8972,
  -41.9071,
  -41.916,
  -41.9231,
  -41.9283,
  -41.9321,
  -41.9352,
  -41.9374,
  -41.9387,
  -41.9386,
  -41.9373,
  -41.9349,
  -41.9316,
  -41.9276,
  -41.9224,
  -41.9162,
  -41.9084,
  -41.8992,
  -41.8883,
  -41.8755,
  -41.8598,
  -41.8408,
  -41.8182,
  -41.7921,
  -41.7637,
  -41.7338,
  -41.7028,
  -41.6714,
  -41.6394,
  -41.6052,
  -41.568,
  -41.5264,
  -41.4795,
  -41.428,
  -41.3726,
  -41.3138,
  -41.2504,
  -41.1816,
  -41.1069,
  -41.0259,
  -40.9383,
  -40.8449,
  -40.7462,
  -40.6435,
  -40.5389,
  -40.4339,
  -36.1806,
  -36.2174,
  -36.2561,
  -36.2957,
  -36.3362,
  -36.3775,
  -36.4194,
  -36.4619,
  -36.5051,
  -36.5489,
  -36.593,
  -36.637,
  -36.6804,
  -36.7229,
  -36.7647,
  -36.8055,
  -36.8446,
  -36.8838,
  -36.9221,
  -36.959,
  -36.9947,
  -37.0297,
  -37.0645,
  -37.0993,
  -37.1338,
  -37.1684,
  -37.2024,
  -37.2359,
  -37.2689,
  -37.3016,
  -37.3341,
  -37.3657,
  -37.3986,
  -37.4321,
  -37.4661,
  -37.5006,
  -37.5351,
  -37.5699,
  -37.605,
  -37.6409,
  -37.6778,
  -37.7157,
  -37.7544,
  -37.7935,
  -37.8323,
  -37.8703,
  -37.9065,
  -37.9429,
  -37.9786,
  -38.0137,
  -38.0481,
  -38.082,
  -38.1153,
  -38.1482,
  -38.1805,
  -38.2119,
  -38.243,
  -38.2737,
  -38.3039,
  -38.3339,
  -38.3639,
  -38.3938,
  -38.424,
  -38.4533,
  -38.4844,
  -38.5163,
  -38.5497,
  -38.5846,
  -38.6213,
  -38.6591,
  -38.6978,
  -38.7366,
  -38.7748,
  -38.8122,
  -38.8485,
  -38.8837,
  -38.9177,
  -38.9509,
  -38.9837,
  -39.0167,
  -39.0491,
  -39.0832,
  -39.1176,
  -39.1517,
  -39.185,
  -39.2173,
  -39.248,
  -39.2777,
  -39.3071,
  -39.337,
  -39.3677,
  -39.3994,
  -39.4318,
  -39.4647,
  -39.4979,
  -39.5314,
  -39.5648,
  -39.5975,
  -39.6287,
  -39.6594,
  -39.6893,
  -39.7185,
  -39.7472,
  -39.7755,
  -39.8028,
  -39.8287,
  -39.8528,
  -39.8748,
  -39.8947,
  -39.9126,
  -39.9287,
  -39.9426,
  -39.9551,
  -39.9662,
  -39.9764,
  -39.9858,
  -39.9944,
  -40.0009,
  -40.0073,
  -40.0128,
  -40.0178,
  -40.0228,
  -40.0283,
  -40.0345,
  -40.0413,
  -40.0487,
  -40.0566,
  -40.0642,
  -40.0719,
  -40.0795,
  -40.0873,
  -40.0954,
  -40.1043,
  -40.1136,
  -40.1236,
  -40.1344,
  -40.1463,
  -40.1584,
  -40.1732,
  -40.1895,
  -40.2071,
  -40.2261,
  -40.2459,
  -40.2663,
  -40.2866,
  -40.3066,
  -40.326,
  -40.345,
  -40.3635,
  -40.382,
  -40.4005,
  -40.4196,
  -40.439,
  -40.4589,
  -40.4787,
  -40.4981,
  -40.5165,
  -40.5339,
  -40.5504,
  -40.5663,
  -40.5807,
  -40.5955,
  -40.6102,
  -40.625,
  -40.6401,
  -40.6554,
  -40.6708,
  -40.6861,
  -40.7016,
  -40.7174,
  -40.7329,
  -40.748,
  -40.7633,
  -40.7786,
  -40.7948,
  -40.8117,
  -40.8297,
  -40.8485,
  -40.8675,
  -40.8866,
  -40.9054,
  -40.9244,
  -40.9443,
  -40.9659,
  -40.9883,
  -41.0143,
  -41.0427,
  -41.0729,
  -41.1038,
  -41.1341,
  -41.1633,
  -41.1905,
  -41.2153,
  -41.2375,
  -41.2575,
  -41.2757,
  -41.293,
  -41.3095,
  -41.3243,
  -41.3378,
  -41.3489,
  -41.3577,
  -41.3641,
  -41.3675,
  -41.3685,
  -41.3682,
  -41.3677,
  -41.3677,
  -41.3689,
  -41.3709,
  -41.3739,
  -41.3773,
  -41.3802,
  -41.3843,
  -41.3884,
  -41.3921,
  -41.3954,
  -41.3987,
  -41.4025,
  -41.4078,
  -41.4154,
  -41.4246,
  -41.4352,
  -41.4464,
  -41.4582,
  -41.4694,
  -41.4801,
  -41.4904,
  -41.5,
  -41.5094,
  -41.5191,
  -41.5295,
  -41.5406,
  -41.5526,
  -41.5649,
  -41.5779,
  -41.5911,
  -41.6048,
  -41.6186,
  -41.6323,
  -41.6459,
  -41.6591,
  -41.6722,
  -41.6849,
  -41.6965,
  -41.7087,
  -41.7209,
  -41.7334,
  -41.7462,
  -41.7595,
  -41.7731,
  -41.7869,
  -41.8008,
  -41.8146,
  -41.8282,
  -41.8409,
  -41.8522,
  -41.8614,
  -41.8683,
  -41.8734,
  -41.8772,
  -41.8807,
  -41.8836,
  -41.886,
  -41.8872,
  -41.8871,
  -41.8858,
  -41.8833,
  -41.8796,
  -41.8748,
  -41.8686,
  -41.861,
  -41.8519,
  -41.8407,
  -41.8275,
  -41.8116,
  -41.7926,
  -41.7701,
  -41.7446,
  -41.7169,
  -41.6877,
  -41.6578,
  -41.6276,
  -41.5967,
  -41.5627,
  -41.5262,
  -41.4853,
  -41.4391,
  -41.3882,
  -41.3332,
  -41.2744,
  -41.2112,
  -41.1425,
  -41.0679,
  -40.9868,
  -40.8991,
  -40.805,
  -40.7052,
  -40.6007,
  -40.4936,
  -40.3866,
  -36.0342,
  -36.0716,
  -36.1099,
  -36.1494,
  -36.1901,
  -36.2319,
  -36.2744,
  -36.3176,
  -36.3613,
  -36.4055,
  -36.4496,
  -36.4922,
  -36.535,
  -36.5769,
  -36.6179,
  -36.6581,
  -36.6976,
  -36.7367,
  -36.7746,
  -36.8115,
  -36.8476,
  -36.883,
  -36.9182,
  -36.9536,
  -36.9889,
  -37.0241,
  -37.0579,
  -37.0925,
  -37.1264,
  -37.1597,
  -37.1925,
  -37.2254,
  -37.2588,
  -37.2929,
  -37.3279,
  -37.3633,
  -37.3988,
  -37.4345,
  -37.4704,
  -37.5069,
  -37.5443,
  -37.5816,
  -37.6204,
  -37.6593,
  -37.698,
  -37.736,
  -37.7732,
  -37.8096,
  -37.8455,
  -37.8808,
  -37.9156,
  -37.9498,
  -37.9834,
  -38.0165,
  -38.049,
  -38.0814,
  -38.1134,
  -38.1441,
  -38.1755,
  -38.2068,
  -38.2379,
  -38.269,
  -38.3004,
  -38.3319,
  -38.364,
  -38.3972,
  -38.4317,
  -38.4679,
  -38.5057,
  -38.5446,
  -38.5841,
  -38.6234,
  -38.6622,
  -38.7,
  -38.7356,
  -38.7711,
  -38.8054,
  -38.839,
  -38.8723,
  -38.9055,
  -38.9393,
  -38.9734,
  -39.0078,
  -39.0422,
  -39.0758,
  -39.1079,
  -39.1391,
  -39.1694,
  -39.1991,
  -39.2292,
  -39.2601,
  -39.2917,
  -39.3234,
  -39.3565,
  -39.3901,
  -39.4236,
  -39.4573,
  -39.4905,
  -39.5232,
  -39.5546,
  -39.5855,
  -39.6156,
  -39.6449,
  -39.6738,
  -39.7015,
  -39.7274,
  -39.7517,
  -39.7736,
  -39.7935,
  -39.8112,
  -39.8269,
  -39.8399,
  -39.8525,
  -39.8641,
  -39.8753,
  -39.8859,
  -39.8958,
  -39.9048,
  -39.9127,
  -39.92,
  -39.9268,
  -39.9333,
  -39.9398,
  -39.9468,
  -39.954,
  -39.9612,
  -39.9688,
  -39.9764,
  -39.9842,
  -39.9921,
  -40.0004,
  -40.0085,
  -40.0179,
  -40.0281,
  -40.0388,
  -40.0502,
  -40.0626,
  -40.076,
  -40.0908,
  -40.1073,
  -40.1252,
  -40.1447,
  -40.1648,
  -40.1854,
  -40.2059,
  -40.2262,
  -40.2457,
  -40.2645,
  -40.2831,
  -40.3015,
  -40.32,
  -40.3388,
  -40.3572,
  -40.3769,
  -40.3966,
  -40.4158,
  -40.4344,
  -40.4521,
  -40.4687,
  -40.4846,
  -40.4995,
  -40.5138,
  -40.5281,
  -40.5424,
  -40.5572,
  -40.5726,
  -40.5882,
  -40.6041,
  -40.62,
  -40.6359,
  -40.6517,
  -40.6666,
  -40.6812,
  -40.6956,
  -40.7105,
  -40.7263,
  -40.7423,
  -40.7602,
  -40.7787,
  -40.7978,
  -40.817,
  -40.8368,
  -40.8579,
  -40.8805,
  -40.9049,
  -40.9323,
  -40.9612,
  -40.9915,
  -41.0223,
  -41.0524,
  -41.0812,
  -41.1084,
  -41.1334,
  -41.1566,
  -41.1781,
  -41.1981,
  -41.217,
  -41.2349,
  -41.2511,
  -41.2651,
  -41.277,
  -41.2859,
  -41.2911,
  -41.2945,
  -41.2954,
  -41.295,
  -41.2945,
  -41.2942,
  -41.295,
  -41.2968,
  -41.2996,
  -41.303,
  -41.3068,
  -41.3108,
  -41.3146,
  -41.3184,
  -41.3219,
  -41.3257,
  -41.3303,
  -41.3365,
  -41.3445,
  -41.3542,
  -41.3651,
  -41.3761,
  -41.3875,
  -41.3986,
  -41.4091,
  -41.4193,
  -41.4292,
  -41.4394,
  -41.4502,
  -41.462,
  -41.4734,
  -41.4864,
  -41.4994,
  -41.5129,
  -41.5267,
  -41.5408,
  -41.555,
  -41.5693,
  -41.5833,
  -41.5971,
  -41.6106,
  -41.6241,
  -41.6371,
  -41.6498,
  -41.6623,
  -41.6749,
  -41.6878,
  -41.7012,
  -41.7151,
  -41.7293,
  -41.7437,
  -41.7582,
  -41.7725,
  -41.7859,
  -41.7976,
  -41.8072,
  -41.8142,
  -41.8192,
  -41.823,
  -41.8265,
  -41.8298,
  -41.8328,
  -41.8348,
  -41.8357,
  -41.8354,
  -41.8337,
  -41.8308,
  -41.8254,
  -41.8199,
  -41.8124,
  -41.8033,
  -41.792,
  -41.7787,
  -41.7626,
  -41.7438,
  -41.7218,
  -41.6969,
  -41.6699,
  -41.6418,
  -41.6132,
  -41.5841,
  -41.5539,
  -41.5221,
  -41.4866,
  -41.4465,
  -41.401,
  -41.3502,
  -41.2953,
  -41.2365,
  -41.1733,
  -41.1044,
  -41.0294,
  -40.9481,
  -40.8598,
  -40.7647,
  -40.6631,
  -40.5561,
  -40.4458,
  -40.3349,
  -35.89,
  -35.9269,
  -35.965,
  -36.0046,
  -36.0457,
  -36.0881,
  -36.1303,
  -36.1743,
  -36.2187,
  -36.2631,
  -36.3071,
  -36.3503,
  -36.3925,
  -36.4336,
  -36.4739,
  -36.5134,
  -36.5524,
  -36.5909,
  -36.6288,
  -36.666,
  -36.7024,
  -36.7377,
  -36.7737,
  -36.8095,
  -36.8454,
  -36.8813,
  -36.9169,
  -36.952,
  -36.9863,
  -37.02,
  -37.053,
  -37.086,
  -37.1196,
  -37.1542,
  -37.1897,
  -37.226,
  -37.2616,
  -37.2984,
  -37.3352,
  -37.3725,
  -37.4105,
  -37.4489,
  -37.4881,
  -37.5269,
  -37.5652,
  -37.603,
  -37.6399,
  -37.6764,
  -37.7123,
  -37.7478,
  -37.7831,
  -37.818,
  -37.8512,
  -37.8849,
  -37.918,
  -37.951,
  -37.9837,
  -38.0162,
  -38.0486,
  -38.0809,
  -38.1132,
  -38.1455,
  -38.1778,
  -38.2106,
  -38.2439,
  -38.2783,
  -38.3143,
  -38.3518,
  -38.3897,
  -38.4297,
  -38.47,
  -38.5098,
  -38.5488,
  -38.5869,
  -38.6236,
  -38.6592,
  -38.6939,
  -38.7277,
  -38.7613,
  -38.7951,
  -38.8293,
  -38.8638,
  -38.8984,
  -38.9328,
  -38.9664,
  -38.9992,
  -39.0297,
  -39.0602,
  -39.0906,
  -39.1209,
  -39.152,
  -39.1843,
  -39.2171,
  -39.2504,
  -39.2839,
  -39.3177,
  -39.3513,
  -39.3847,
  -39.4176,
  -39.4498,
  -39.4815,
  -39.5124,
  -39.5424,
  -39.5715,
  -39.5983,
  -39.6244,
  -39.6488,
  -39.6711,
  -39.691,
  -39.7088,
  -39.7247,
  -39.739,
  -39.7523,
  -39.765,
  -39.7769,
  -39.7887,
  -39.7997,
  -39.81,
  -39.8192,
  -39.8278,
  -39.8359,
  -39.8437,
  -39.8516,
  -39.8592,
  -39.8656,
  -39.8731,
  -39.8806,
  -39.8879,
  -39.8957,
  -39.9038,
  -39.9126,
  -39.9222,
  -39.9324,
  -39.9435,
  -39.9553,
  -39.9677,
  -39.9808,
  -39.9949,
  -40.0102,
  -40.0271,
  -40.0454,
  -40.0652,
  -40.0858,
  -40.1068,
  -40.1276,
  -40.1469,
  -40.1665,
  -40.1855,
  -40.2039,
  -40.2221,
  -40.2403,
  -40.259,
  -40.278,
  -40.2973,
  -40.3165,
  -40.3355,
  -40.354,
  -40.3717,
  -40.3884,
  -40.4041,
  -40.4187,
  -40.4327,
  -40.4464,
  -40.4604,
  -40.4749,
  -40.4901,
  -40.5057,
  -40.5219,
  -40.5373,
  -40.5533,
  -40.5689,
  -40.5838,
  -40.5977,
  -40.6113,
  -40.6252,
  -40.6401,
  -40.6561,
  -40.6732,
  -40.6912,
  -40.7103,
  -40.73,
  -40.7506,
  -40.7728,
  -40.7964,
  -40.8223,
  -40.8501,
  -40.8799,
  -40.9102,
  -40.941,
  -40.9706,
  -40.999,
  -41.0263,
  -41.0517,
  -41.0749,
  -41.0978,
  -41.1196,
  -41.14,
  -41.1593,
  -41.1768,
  -41.1919,
  -41.204,
  -41.2133,
  -41.2192,
  -41.2225,
  -41.2236,
  -41.2238,
  -41.2232,
  -41.2226,
  -41.2232,
  -41.2248,
  -41.2273,
  -41.2304,
  -41.234,
  -41.2378,
  -41.2417,
  -41.2456,
  -41.2496,
  -41.254,
  -41.2593,
  -41.2662,
  -41.2747,
  -41.2849,
  -41.2948,
  -41.3062,
  -41.3174,
  -41.3278,
  -41.338,
  -41.348,
  -41.358,
  -41.3687,
  -41.3804,
  -41.3932,
  -41.4067,
  -41.4208,
  -41.4348,
  -41.4489,
  -41.4631,
  -41.4778,
  -41.4923,
  -41.5071,
  -41.5214,
  -41.5356,
  -41.5499,
  -41.5638,
  -41.5774,
  -41.5906,
  -41.6035,
  -41.6162,
  -41.6294,
  -41.643,
  -41.6572,
  -41.672,
  -41.6871,
  -41.7022,
  -41.7171,
  -41.7312,
  -41.7426,
  -41.7526,
  -41.7599,
  -41.7648,
  -41.7685,
  -41.7719,
  -41.7753,
  -41.7785,
  -41.7809,
  -41.7824,
  -41.7828,
  -41.7819,
  -41.7797,
  -41.776,
  -41.7711,
  -41.7643,
  -41.7556,
  -41.7444,
  -41.7308,
  -41.7152,
  -41.6964,
  -41.6749,
  -41.651,
  -41.625,
  -41.5979,
  -41.5705,
  -41.5424,
  -41.5132,
  -41.4817,
  -41.447,
  -41.4078,
  -41.3631,
  -41.3133,
  -41.2587,
  -41.1998,
  -41.1362,
  -41.067,
  -40.9917,
  -40.9099,
  -40.8208,
  -40.7243,
  -40.6204,
  -40.5104,
  -40.3962,
  -40.2809,
  -35.747,
  -35.7836,
  -35.8207,
  -35.8606,
  -35.9022,
  -35.9453,
  -35.9893,
  -36.034,
  -36.0789,
  -36.1235,
  -36.1674,
  -36.21,
  -36.2514,
  -36.2917,
  -36.3312,
  -36.3702,
  -36.4077,
  -36.446,
  -36.4839,
  -36.5214,
  -36.5585,
  -36.5955,
  -36.6321,
  -36.6686,
  -36.7051,
  -36.7415,
  -36.7776,
  -36.813,
  -36.8476,
  -36.8813,
  -36.9144,
  -36.9464,
  -36.9801,
  -37.015,
  -37.0512,
  -37.0883,
  -37.1259,
  -37.1636,
  -37.2014,
  -37.2396,
  -37.2782,
  -37.3172,
  -37.3562,
  -37.3948,
  -37.4329,
  -37.4702,
  -37.5069,
  -37.5422,
  -37.5784,
  -37.6144,
  -37.6504,
  -37.6859,
  -37.7209,
  -37.7553,
  -37.7892,
  -37.8228,
  -37.8562,
  -37.8894,
  -37.9225,
  -37.9557,
  -37.9888,
  -38.022,
  -38.0555,
  -38.0885,
  -38.1231,
  -38.1589,
  -38.1961,
  -38.2349,
  -38.2749,
  -38.3158,
  -38.3566,
  -38.3971,
  -38.4364,
  -38.4744,
  -38.5112,
  -38.547,
  -38.5817,
  -38.6158,
  -38.6497,
  -38.684,
  -38.7177,
  -38.7526,
  -38.7876,
  -38.8223,
  -38.8563,
  -38.8894,
  -38.9216,
  -38.9529,
  -38.9839,
  -39.0149,
  -39.0463,
  -39.0785,
  -39.1114,
  -39.1448,
  -39.1785,
  -39.2123,
  -39.2461,
  -39.2798,
  -39.312,
  -39.3448,
  -39.3769,
  -39.4082,
  -39.4387,
  -39.4678,
  -39.4956,
  -39.5218,
  -39.5464,
  -39.5689,
  -39.5891,
  -39.6075,
  -39.6241,
  -39.6392,
  -39.6533,
  -39.6668,
  -39.6802,
  -39.6931,
  -39.7053,
  -39.7153,
  -39.7256,
  -39.7354,
  -39.7448,
  -39.7541,
  -39.763,
  -39.7714,
  -39.7791,
  -39.7864,
  -39.7936,
  -39.8006,
  -39.8081,
  -39.8163,
  -39.8254,
  -39.8353,
  -39.8462,
  -39.8581,
  -39.8707,
  -39.884,
  -39.8984,
  -39.9137,
  -39.9289,
  -39.9464,
  -39.9653,
  -39.9854,
  -40.0062,
  -40.0274,
  -40.0485,
  -40.069,
  -40.0889,
  -40.1082,
  -40.1268,
  -40.1449,
  -40.1628,
  -40.1809,
  -40.1994,
  -40.218,
  -40.2369,
  -40.2553,
  -40.2734,
  -40.2906,
  -40.3071,
  -40.3225,
  -40.336,
  -40.3498,
  -40.3633,
  -40.3772,
  -40.3915,
  -40.4066,
  -40.4225,
  -40.439,
  -40.4556,
  -40.472,
  -40.4878,
  -40.5023,
  -40.516,
  -40.5289,
  -40.5422,
  -40.5562,
  -40.5714,
  -40.5877,
  -40.605,
  -40.6236,
  -40.6434,
  -40.6646,
  -40.6875,
  -40.7124,
  -40.7382,
  -40.7669,
  -40.7969,
  -40.8275,
  -40.8581,
  -40.8877,
  -40.9161,
  -40.9432,
  -40.9693,
  -40.9945,
  -41.0187,
  -41.0419,
  -41.0639,
  -41.0844,
  -41.1031,
  -41.119,
  -41.132,
  -41.1415,
  -41.1479,
  -41.1517,
  -41.1532,
  -41.1535,
  -41.1532,
  -41.1529,
  -41.1531,
  -41.1542,
  -41.156,
  -41.1587,
  -41.1611,
  -41.165,
  -41.1691,
  -41.1733,
  -41.1775,
  -41.1825,
  -41.1884,
  -41.1959,
  -41.2051,
  -41.2156,
  -41.2267,
  -41.2379,
  -41.2489,
  -41.2592,
  -41.2689,
  -41.2786,
  -41.2886,
  -41.2996,
  -41.3119,
  -41.3256,
  -41.3401,
  -41.3549,
  -41.3698,
  -41.3844,
  -41.399,
  -41.4138,
  -41.4288,
  -41.4439,
  -41.4589,
  -41.4739,
  -41.4887,
  -41.5034,
  -41.5166,
  -41.5303,
  -41.5435,
  -41.5566,
  -41.57,
  -41.584,
  -41.5988,
  -41.614,
  -41.6297,
  -41.6454,
  -41.661,
  -41.6757,
  -41.6889,
  -41.6994,
  -41.7071,
  -41.7122,
  -41.7157,
  -41.7187,
  -41.7219,
  -41.7251,
  -41.7278,
  -41.7297,
  -41.7307,
  -41.7307,
  -41.7293,
  -41.7266,
  -41.7223,
  -41.7162,
  -41.708,
  -41.6974,
  -41.6841,
  -41.6682,
  -41.6498,
  -41.6289,
  -41.6057,
  -41.5809,
  -41.5551,
  -41.5288,
  -41.5016,
  -41.4732,
  -41.4412,
  -41.407,
  -41.3682,
  -41.3247,
  -41.2759,
  -41.2222,
  -41.1634,
  -41.0996,
  -41.0303,
  -40.9545,
  -40.8722,
  -40.7823,
  -40.6843,
  -40.5781,
  -40.4647,
  -40.3463,
  -40.2258,
  -35.6049,
  -35.6414,
  -35.6795,
  -35.7197,
  -35.7617,
  -35.8054,
  -35.8502,
  -35.8955,
  -35.9408,
  -35.9854,
  -36.0288,
  -36.0698,
  -36.1105,
  -36.15,
  -36.1889,
  -36.2274,
  -36.2658,
  -36.3039,
  -36.342,
  -36.38,
  -36.4178,
  -36.4553,
  -36.4928,
  -36.5299,
  -36.5668,
  -36.6036,
  -36.6388,
  -36.6744,
  -36.709,
  -36.7426,
  -36.7759,
  -36.8093,
  -36.8433,
  -36.8785,
  -36.9151,
  -36.9528,
  -36.9911,
  -37.0296,
  -37.0684,
  -37.1073,
  -37.1465,
  -37.1847,
  -37.2238,
  -37.2623,
  -37.3001,
  -37.3371,
  -37.3736,
  -37.4098,
  -37.4463,
  -37.4829,
  -37.5198,
  -37.5564,
  -37.5924,
  -37.6276,
  -37.6622,
  -37.6963,
  -37.7302,
  -37.7627,
  -37.7963,
  -37.83,
  -37.864,
  -37.8982,
  -37.9328,
  -37.9679,
  -38.0039,
  -38.041,
  -38.0793,
  -38.1192,
  -38.16,
  -38.2016,
  -38.2431,
  -38.2838,
  -38.3233,
  -38.3616,
  -38.3976,
  -38.4334,
  -38.4683,
  -38.5025,
  -38.5368,
  -38.5714,
  -38.6065,
  -38.6419,
  -38.6773,
  -38.7125,
  -38.747,
  -38.7807,
  -38.8137,
  -38.8462,
  -38.8782,
  -38.9098,
  -38.9415,
  -38.9737,
  -39.0055,
  -39.039,
  -39.0728,
  -39.1069,
  -39.1411,
  -39.1749,
  -39.2084,
  -39.242,
  -39.2746,
  -39.3063,
  -39.3368,
  -39.3657,
  -39.3934,
  -39.4194,
  -39.4438,
  -39.4666,
  -39.4873,
  -39.5066,
  -39.5242,
  -39.5392,
  -39.5543,
  -39.5692,
  -39.5834,
  -39.5971,
  -39.61,
  -39.6218,
  -39.6328,
  -39.6435,
  -39.6543,
  -39.6649,
  -39.6751,
  -39.6844,
  -39.6926,
  -39.6998,
  -39.7065,
  -39.7134,
  -39.7208,
  -39.729,
  -39.7383,
  -39.7475,
  -39.7586,
  -39.7708,
  -39.784,
  -39.7984,
  -39.8137,
  -39.83,
  -39.8472,
  -39.8655,
  -39.8851,
  -39.9057,
  -39.9269,
  -39.9483,
  -39.9695,
  -39.9903,
  -40.0104,
  -40.0298,
  -40.0486,
  -40.0671,
  -40.0851,
  -40.103,
  -40.12,
  -40.1383,
  -40.1566,
  -40.1746,
  -40.1919,
  -40.2085,
  -40.2243,
  -40.2391,
  -40.2533,
  -40.2671,
  -40.2808,
  -40.2948,
  -40.3093,
  -40.3245,
  -40.3405,
  -40.3572,
  -40.3742,
  -40.391,
  -40.4069,
  -40.4214,
  -40.4348,
  -40.4475,
  -40.4601,
  -40.4733,
  -40.4866,
  -40.502,
  -40.5186,
  -40.5367,
  -40.5564,
  -40.5779,
  -40.6015,
  -40.6272,
  -40.655,
  -40.6843,
  -40.7147,
  -40.7454,
  -40.776,
  -40.8057,
  -40.8342,
  -40.8617,
  -40.8885,
  -40.9146,
  -40.9399,
  -40.9644,
  -40.9876,
  -41.0092,
  -41.0287,
  -41.0455,
  -41.0592,
  -41.0694,
  -41.0755,
  -41.0802,
  -41.0825,
  -41.0835,
  -41.0836,
  -41.0832,
  -41.0832,
  -41.0837,
  -41.0851,
  -41.0875,
  -41.0908,
  -41.0945,
  -41.0987,
  -41.1029,
  -41.1075,
  -41.113,
  -41.1193,
  -41.1274,
  -41.1369,
  -41.1479,
  -41.1591,
  -41.1703,
  -41.1811,
  -41.1911,
  -41.2005,
  -41.2098,
  -41.2197,
  -41.2311,
  -41.244,
  -41.2583,
  -41.2734,
  -41.2877,
  -41.3029,
  -41.3177,
  -41.3327,
  -41.3478,
  -41.3632,
  -41.3788,
  -41.3946,
  -41.4103,
  -41.4261,
  -41.4416,
  -41.4567,
  -41.471,
  -41.4848,
  -41.4982,
  -41.512,
  -41.5263,
  -41.5415,
  -41.5573,
  -41.5734,
  -41.5898,
  -41.6059,
  -41.6212,
  -41.635,
  -41.6463,
  -41.6545,
  -41.6597,
  -41.6632,
  -41.6659,
  -41.6688,
  -41.6717,
  -41.6746,
  -41.677,
  -41.6787,
  -41.6795,
  -41.679,
  -41.6773,
  -41.6728,
  -41.6672,
  -41.6594,
  -41.6493,
  -41.6363,
  -41.6207,
  -41.6025,
  -41.5821,
  -41.56,
  -41.5365,
  -41.5121,
  -41.4869,
  -41.4608,
  -41.4327,
  -41.4021,
  -41.368,
  -41.3301,
  -41.2874,
  -41.2402,
  -41.1877,
  -41.1297,
  -41.0659,
  -40.9965,
  -40.9207,
  -40.838,
  -40.7475,
  -40.6482,
  -40.5397,
  -40.4231,
  -40.3005,
  -40.1749,
  -35.4659,
  -35.5026,
  -35.5409,
  -35.5812,
  -35.6236,
  -35.6676,
  -35.7128,
  -35.7575,
  -35.8029,
  -35.8473,
  -35.8903,
  -35.9317,
  -35.9717,
  -36.0107,
  -36.0492,
  -36.0875,
  -36.1256,
  -36.1639,
  -36.2022,
  -36.2405,
  -36.2786,
  -36.3157,
  -36.3538,
  -36.3914,
  -36.4286,
  -36.4654,
  -36.5018,
  -36.5374,
  -36.5723,
  -36.6061,
  -36.6396,
  -36.6736,
  -36.7083,
  -36.7436,
  -36.7806,
  -36.8187,
  -36.8565,
  -36.8957,
  -36.9352,
  -36.9748,
  -37.0146,
  -37.0543,
  -37.0934,
  -37.1318,
  -37.1691,
  -37.2058,
  -37.2422,
  -37.2789,
  -37.3157,
  -37.3532,
  -37.391,
  -37.4286,
  -37.4644,
  -37.5005,
  -37.5359,
  -37.5706,
  -37.6048,
  -37.6387,
  -37.6727,
  -37.7069,
  -37.7415,
  -37.7764,
  -37.8119,
  -37.8479,
  -37.885,
  -37.9232,
  -37.9627,
  -38.0033,
  -38.0448,
  -38.0859,
  -38.128,
  -38.1691,
  -38.2091,
  -38.2476,
  -38.2848,
  -38.3208,
  -38.3559,
  -38.3906,
  -38.425,
  -38.4598,
  -38.4954,
  -38.5313,
  -38.5672,
  -38.6029,
  -38.638,
  -38.6727,
  -38.7058,
  -38.7394,
  -38.7724,
  -38.8048,
  -38.8369,
  -38.8693,
  -38.902,
  -38.9353,
  -38.9692,
  -39.0032,
  -39.0374,
  -39.0721,
  -39.1059,
  -39.1394,
  -39.1726,
  -39.2048,
  -39.2355,
  -39.2646,
  -39.2911,
  -39.317,
  -39.3416,
  -39.3647,
  -39.386,
  -39.4062,
  -39.4246,
  -39.4416,
  -39.4577,
  -39.4731,
  -39.4881,
  -39.5021,
  -39.5154,
  -39.5276,
  -39.5392,
  -39.5508,
  -39.5626,
  -39.5743,
  -39.5855,
  -39.5956,
  -39.6034,
  -39.611,
  -39.618,
  -39.6249,
  -39.6323,
  -39.6405,
  -39.6497,
  -39.6601,
  -39.6712,
  -39.6835,
  -39.6974,
  -39.7124,
  -39.7287,
  -39.7461,
  -39.7645,
  -39.7837,
  -39.8036,
  -39.8244,
  -39.8458,
  -39.8677,
  -39.8894,
  -39.9096,
  -39.9302,
  -39.95,
  -39.9693,
  -39.9879,
  -40.0062,
  -40.0243,
  -40.0423,
  -40.0601,
  -40.0777,
  -40.0951,
  -40.1117,
  -40.1274,
  -40.1425,
  -40.1572,
  -40.1714,
  -40.1851,
  -40.1991,
  -40.2134,
  -40.2281,
  -40.2435,
  -40.2598,
  -40.2766,
  -40.2928,
  -40.3097,
  -40.3258,
  -40.3405,
  -40.3536,
  -40.3659,
  -40.378,
  -40.3904,
  -40.4041,
  -40.4185,
  -40.4343,
  -40.452,
  -40.4716,
  -40.4935,
  -40.5179,
  -40.5444,
  -40.5729,
  -40.6027,
  -40.6335,
  -40.6646,
  -40.6952,
  -40.7251,
  -40.7539,
  -40.7819,
  -40.8093,
  -40.8351,
  -40.8611,
  -40.8862,
  -40.91,
  -40.9323,
  -40.9525,
  -40.9703,
  -40.9851,
  -40.9964,
  -41.0047,
  -41.0103,
  -41.0133,
  -41.015,
  -41.0155,
  -41.0154,
  -41.0152,
  -41.0156,
  -41.0165,
  -41.0187,
  -41.0217,
  -41.0253,
  -41.0294,
  -41.0339,
  -41.0388,
  -41.0444,
  -41.0512,
  -41.0599,
  -41.0697,
  -41.0805,
  -41.0905,
  -41.1016,
  -41.1123,
  -41.1219,
  -41.1315,
  -41.1408,
  -41.1511,
  -41.1626,
  -41.1758,
  -41.1904,
  -41.2058,
  -41.2214,
  -41.2367,
  -41.2518,
  -41.2668,
  -41.2822,
  -41.298,
  -41.3144,
  -41.331,
  -41.3478,
  -41.3646,
  -41.3812,
  -41.3972,
  -41.4121,
  -41.4264,
  -41.4402,
  -41.4542,
  -41.4689,
  -41.4844,
  -41.5007,
  -41.5174,
  -41.5341,
  -41.5507,
  -41.5665,
  -41.5808,
  -41.5915,
  -41.6003,
  -41.6057,
  -41.6092,
  -41.6119,
  -41.6145,
  -41.6173,
  -41.6203,
  -41.6232,
  -41.6257,
  -41.6274,
  -41.628,
  -41.6275,
  -41.6245,
  -41.6194,
  -41.6124,
  -41.6026,
  -41.5901,
  -41.5749,
  -41.5571,
  -41.5374,
  -41.5163,
  -41.4941,
  -41.4711,
  -41.4473,
  -41.4219,
  -41.3945,
  -41.3642,
  -41.3302,
  -41.2926,
  -41.2509,
  -41.2048,
  -41.1536,
  -41.0969,
  -41.0337,
  -40.9646,
  -40.8893,
  -40.8068,
  -40.716,
  -40.6159,
  -40.5057,
  -40.3865,
  -40.2601,
  -40.1299,
  -35.3292,
  -35.3663,
  -35.4039,
  -35.4443,
  -35.4866,
  -35.5308,
  -35.576,
  -35.6218,
  -35.667,
  -35.7112,
  -35.7536,
  -35.7944,
  -35.834,
  -35.8727,
  -35.911,
  -35.9494,
  -35.9867,
  -36.0251,
  -36.0635,
  -36.1019,
  -36.1403,
  -36.1787,
  -36.2169,
  -36.2549,
  -36.2924,
  -36.3295,
  -36.3662,
  -36.402,
  -36.437,
  -36.4715,
  -36.5057,
  -36.5393,
  -36.5745,
  -36.6103,
  -36.6473,
  -36.6855,
  -36.7245,
  -36.7641,
  -36.8041,
  -36.8445,
  -36.885,
  -36.9251,
  -36.9643,
  -37.0025,
  -37.0398,
  -37.0765,
  -37.113,
  -37.1489,
  -37.1864,
  -37.2249,
  -37.2635,
  -37.3018,
  -37.3397,
  -37.3766,
  -37.4126,
  -37.4477,
  -37.4823,
  -37.5165,
  -37.5506,
  -37.5852,
  -37.6204,
  -37.6559,
  -37.6921,
  -37.7281,
  -37.7661,
  -37.8051,
  -37.8452,
  -37.8865,
  -37.9286,
  -37.9712,
  -38.0136,
  -38.0551,
  -38.0955,
  -38.1345,
  -38.1721,
  -38.2086,
  -38.2442,
  -38.2792,
  -38.314,
  -38.3494,
  -38.3843,
  -38.4205,
  -38.457,
  -38.4932,
  -38.5291,
  -38.5647,
  -38.5998,
  -38.6345,
  -38.6684,
  -38.7016,
  -38.7342,
  -38.7668,
  -38.7996,
  -38.8329,
  -38.8668,
  -38.9009,
  -38.9351,
  -38.9695,
  -39.0029,
  -39.037,
  -39.0707,
  -39.1034,
  -39.1343,
  -39.1634,
  -39.1909,
  -39.2171,
  -39.2419,
  -39.2653,
  -39.2874,
  -39.3082,
  -39.3274,
  -39.3454,
  -39.3621,
  -39.3782,
  -39.3934,
  -39.4079,
  -39.4213,
  -39.4329,
  -39.4448,
  -39.4569,
  -39.4692,
  -39.4815,
  -39.4933,
  -39.5041,
  -39.5137,
  -39.5221,
  -39.5297,
  -39.537,
  -39.5447,
  -39.5531,
  -39.5626,
  -39.5731,
  -39.5845,
  -39.597,
  -39.6114,
  -39.6271,
  -39.6442,
  -39.6626,
  -39.6807,
  -39.7004,
  -39.7209,
  -39.7419,
  -39.7634,
  -39.7854,
  -39.8074,
  -39.8291,
  -39.8504,
  -39.871,
  -39.8909,
  -39.9099,
  -39.928,
  -39.9459,
  -39.9636,
  -39.9812,
  -39.9984,
  -40.0152,
  -40.0314,
  -40.0467,
  -40.0612,
  -40.0756,
  -40.0887,
  -40.1029,
  -40.1174,
  -40.1321,
  -40.1472,
  -40.1628,
  -40.1792,
  -40.1963,
  -40.2134,
  -40.2304,
  -40.2466,
  -40.2613,
  -40.2746,
  -40.2868,
  -40.2986,
  -40.3105,
  -40.3233,
  -40.337,
  -40.3525,
  -40.3699,
  -40.3896,
  -40.412,
  -40.4369,
  -40.4644,
  -40.4936,
  -40.5226,
  -40.5535,
  -40.5847,
  -40.6152,
  -40.645,
  -40.6743,
  -40.7029,
  -40.7305,
  -40.7577,
  -40.7841,
  -40.8094,
  -40.8334,
  -40.8562,
  -40.8772,
  -40.8958,
  -40.9114,
  -40.9237,
  -40.9331,
  -40.9397,
  -40.9441,
  -40.9467,
  -40.9479,
  -40.948,
  -40.9481,
  -40.9482,
  -40.9489,
  -40.9508,
  -40.9526,
  -40.956,
  -40.96,
  -40.9646,
  -40.9697,
  -40.9757,
  -40.9829,
  -40.9914,
  -41.0009,
  -41.0115,
  -41.0224,
  -41.0329,
  -41.0437,
  -41.0538,
  -41.0634,
  -41.0733,
  -41.0841,
  -41.0961,
  -41.1096,
  -41.1243,
  -41.1398,
  -41.1554,
  -41.1706,
  -41.1856,
  -41.2007,
  -41.2164,
  -41.2329,
  -41.2501,
  -41.2679,
  -41.2858,
  -41.3038,
  -41.3214,
  -41.3372,
  -41.3528,
  -41.3674,
  -41.3815,
  -41.3958,
  -41.4107,
  -41.4265,
  -41.4431,
  -41.46,
  -41.4772,
  -41.494,
  -41.51,
  -41.5246,
  -41.5369,
  -41.5461,
  -41.5522,
  -41.5561,
  -41.5587,
  -41.5613,
  -41.5642,
  -41.5674,
  -41.5706,
  -41.5739,
  -41.5767,
  -41.5783,
  -41.5783,
  -41.5762,
  -41.572,
  -41.5653,
  -41.5559,
  -41.5443,
  -41.5294,
  -41.5124,
  -41.4934,
  -41.4732,
  -41.4525,
  -41.4311,
  -41.4089,
  -41.3845,
  -41.3575,
  -41.3274,
  -41.2928,
  -41.2555,
  -41.2144,
  -41.1693,
  -41.1195,
  -41.0639,
  -41.002,
  -40.9336,
  -40.8594,
  -40.7776,
  -40.6872,
  -40.587,
  -40.4761,
  -40.3551,
  -40.226,
  -40.0922,
  -35.1935,
  -35.2312,
  -35.2701,
  -35.3106,
  -35.3529,
  -35.3968,
  -35.4418,
  -35.4873,
  -35.5323,
  -35.576,
  -35.618,
  -35.6574,
  -35.6968,
  -35.7355,
  -35.774,
  -35.8124,
  -35.8509,
  -35.8894,
  -35.9279,
  -35.9662,
  -36.0046,
  -36.0429,
  -36.0812,
  -36.1193,
  -36.1571,
  -36.1945,
  -36.2305,
  -36.2668,
  -36.3025,
  -36.3378,
  -36.3731,
  -36.4087,
  -36.4442,
  -36.4804,
  -36.5172,
  -36.5551,
  -36.5942,
  -36.6343,
  -36.6749,
  -36.7159,
  -36.7569,
  -36.7973,
  -36.8358,
  -36.874,
  -36.9113,
  -36.9483,
  -36.9852,
  -37.0225,
  -37.0606,
  -37.0996,
  -37.1389,
  -37.1781,
  -37.2167,
  -37.2544,
  -37.291,
  -37.3266,
  -37.3615,
  -37.3959,
  -37.4295,
  -37.4644,
  -37.4998,
  -37.5359,
  -37.5726,
  -37.6101,
  -37.6485,
  -37.6881,
  -37.7289,
  -37.7708,
  -37.8133,
  -37.8561,
  -37.8988,
  -37.941,
  -37.982,
  -38.0216,
  -38.0598,
  -38.0958,
  -38.132,
  -38.1677,
  -38.2034,
  -38.2394,
  -38.2754,
  -38.312,
  -38.3489,
  -38.3861,
  -38.4227,
  -38.4591,
  -38.4952,
  -38.5307,
  -38.5654,
  -38.5993,
  -38.6325,
  -38.6654,
  -38.6973,
  -38.7307,
  -38.7644,
  -38.7984,
  -38.8327,
  -38.8673,
  -38.902,
  -38.9366,
  -38.9707,
  -39.0038,
  -39.0352,
  -39.0646,
  -39.0923,
  -39.1185,
  -39.1437,
  -39.1678,
  -39.1905,
  -39.2118,
  -39.2318,
  -39.2493,
  -39.2666,
  -39.2831,
  -39.2988,
  -39.3133,
  -39.3269,
  -39.3395,
  -39.3517,
  -39.3639,
  -39.3766,
  -39.3892,
  -39.4014,
  -39.4127,
  -39.4229,
  -39.4321,
  -39.4405,
  -39.4486,
  -39.4569,
  -39.4658,
  -39.4755,
  -39.4851,
  -39.4966,
  -39.5096,
  -39.5242,
  -39.5406,
  -39.5587,
  -39.5779,
  -39.5979,
  -39.6183,
  -39.6391,
  -39.6604,
  -39.682,
  -39.704,
  -39.7263,
  -39.7482,
  -39.7701,
  -39.7913,
  -39.8116,
  -39.8309,
  -39.8494,
  -39.8673,
  -39.8848,
  -39.9009,
  -39.9175,
  -39.9338,
  -39.9498,
  -39.965,
  -39.9796,
  -39.9941,
  -40.0085,
  -40.0229,
  -40.0377,
  -40.0527,
  -40.0682,
  -40.084,
  -40.1007,
  -40.1177,
  -40.1349,
  -40.1521,
  -40.1684,
  -40.1832,
  -40.1967,
  -40.2089,
  -40.2205,
  -40.232,
  -40.2433,
  -40.2566,
  -40.272,
  -40.2896,
  -40.3098,
  -40.3327,
  -40.3583,
  -40.3862,
  -40.4155,
  -40.4461,
  -40.4771,
  -40.5079,
  -40.5383,
  -40.5682,
  -40.5974,
  -40.6264,
  -40.6545,
  -40.6819,
  -40.7083,
  -40.7337,
  -40.7578,
  -40.7805,
  -40.8017,
  -40.8208,
  -40.8374,
  -40.8509,
  -40.8616,
  -40.8682,
  -40.8736,
  -40.8773,
  -40.8792,
  -40.88,
  -40.8803,
  -40.8805,
  -40.8812,
  -40.8826,
  -40.885,
  -40.8882,
  -40.8921,
  -40.8966,
  -40.9019,
  -40.9081,
  -40.9154,
  -40.9237,
  -40.9329,
  -40.9429,
  -40.9534,
  -40.9639,
  -40.9744,
  -40.985,
  -40.9953,
  -41.0061,
  -41.0177,
  -41.0303,
  -41.0441,
  -41.0588,
  -41.0742,
  -41.0885,
  -41.1037,
  -41.1187,
  -41.134,
  -41.1502,
  -41.1674,
  -41.1858,
  -41.2047,
  -41.2241,
  -41.2432,
  -41.2617,
  -41.2791,
  -41.2951,
  -41.3101,
  -41.3243,
  -41.3387,
  -41.3538,
  -41.3697,
  -41.3864,
  -41.4035,
  -41.4206,
  -41.4374,
  -41.4535,
  -41.4682,
  -41.4809,
  -41.4908,
  -41.4978,
  -41.5024,
  -41.5055,
  -41.5083,
  -41.5113,
  -41.5147,
  -41.5184,
  -41.5224,
  -41.526,
  -41.5286,
  -41.5294,
  -41.527,
  -41.5232,
  -41.5171,
  -41.5087,
  -41.4973,
  -41.4834,
  -41.4671,
  -41.4491,
  -41.4302,
  -41.411,
  -41.3913,
  -41.3704,
  -41.3473,
  -41.3209,
  -41.2911,
  -41.258,
  -41.2214,
  -41.1809,
  -41.1366,
  -41.0876,
  -41.0332,
  -40.9727,
  -40.9056,
  -40.8325,
  -40.7519,
  -40.6625,
  -40.5632,
  -40.4526,
  -40.3312,
  -40.2009,
  -40.0651,
  -35.0604,
  -35.0989,
  -35.1382,
  -35.1788,
  -35.2209,
  -35.2644,
  -35.3091,
  -35.3532,
  -35.3977,
  -35.4409,
  -35.4826,
  -35.5229,
  -35.5623,
  -35.6013,
  -35.64,
  -35.6786,
  -35.7172,
  -35.7556,
  -35.794,
  -35.8321,
  -35.8702,
  -35.9073,
  -35.9454,
  -35.9835,
  -36.0215,
  -36.0593,
  -36.0967,
  -36.1339,
  -36.1706,
  -36.2072,
  -36.2438,
  -36.2802,
  -36.3166,
  -36.3528,
  -36.3894,
  -36.427,
  -36.4662,
  -36.5056,
  -36.5468,
  -36.5884,
  -36.6299,
  -36.6706,
  -36.7101,
  -36.7486,
  -36.7862,
  -36.8234,
  -36.8608,
  -36.8986,
  -36.9372,
  -36.9766,
  -37.0164,
  -37.0561,
  -37.0943,
  -37.1326,
  -37.17,
  -37.2062,
  -37.2414,
  -37.2762,
  -37.311,
  -37.346,
  -37.3817,
  -37.4179,
  -37.455,
  -37.4929,
  -37.5317,
  -37.5718,
  -37.6131,
  -37.6553,
  -37.6981,
  -37.7402,
  -37.7833,
  -37.8257,
  -37.8674,
  -37.9076,
  -37.9464,
  -37.9842,
  -38.0213,
  -38.0581,
  -38.0944,
  -38.1311,
  -38.1683,
  -38.2053,
  -38.2428,
  -38.2805,
  -38.3181,
  -38.3551,
  -38.3911,
  -38.4273,
  -38.4628,
  -38.4971,
  -38.5307,
  -38.5639,
  -38.5972,
  -38.6305,
  -38.6642,
  -38.698,
  -38.7322,
  -38.7667,
  -38.8018,
  -38.8369,
  -38.8716,
  -38.9052,
  -38.9371,
  -38.9669,
  -38.9949,
  -39.0206,
  -39.0463,
  -39.0708,
  -39.0941,
  -39.1159,
  -39.1362,
  -39.1548,
  -39.1728,
  -39.1896,
  -39.2053,
  -39.2206,
  -39.2343,
  -39.2471,
  -39.2594,
  -39.2718,
  -39.2844,
  -39.297,
  -39.3094,
  -39.321,
  -39.3307,
  -39.3407,
  -39.35,
  -39.3588,
  -39.3678,
  -39.3772,
  -39.3873,
  -39.3981,
  -39.4099,
  -39.423,
  -39.4381,
  -39.4552,
  -39.474,
  -39.4941,
  -39.5149,
  -39.536,
  -39.5572,
  -39.5786,
  -39.6005,
  -39.6226,
  -39.645,
  -39.6664,
  -39.6886,
  -39.7102,
  -39.7309,
  -39.7507,
  -39.7695,
  -39.7875,
  -39.8049,
  -39.8216,
  -39.838,
  -39.8539,
  -39.8696,
  -39.8849,
  -39.8997,
  -39.9143,
  -39.929,
  -39.9437,
  -39.9588,
  -39.9742,
  -39.9898,
  -40.0061,
  -40.0227,
  -40.0401,
  -40.0565,
  -40.0736,
  -40.0896,
  -40.1046,
  -40.1181,
  -40.1305,
  -40.1423,
  -40.1538,
  -40.1659,
  -40.1797,
  -40.1952,
  -40.2134,
  -40.2341,
  -40.2576,
  -40.2837,
  -40.3121,
  -40.3419,
  -40.3727,
  -40.4038,
  -40.4344,
  -40.4643,
  -40.494,
  -40.5233,
  -40.5522,
  -40.5805,
  -40.6079,
  -40.6334,
  -40.6587,
  -40.6826,
  -40.7052,
  -40.7262,
  -40.7457,
  -40.7628,
  -40.7771,
  -40.7887,
  -40.7978,
  -40.8043,
  -40.8088,
  -40.8116,
  -40.8131,
  -40.8136,
  -40.8139,
  -40.8146,
  -40.816,
  -40.818,
  -40.8207,
  -40.8243,
  -40.8287,
  -40.8339,
  -40.8403,
  -40.8475,
  -40.8557,
  -40.8646,
  -40.8741,
  -40.884,
  -40.8932,
  -40.9037,
  -40.9145,
  -40.9257,
  -40.9376,
  -40.9502,
  -40.9636,
  -40.978,
  -40.9928,
  -41.0081,
  -41.0234,
  -41.0385,
  -41.0536,
  -41.0694,
  -41.0861,
  -41.1043,
  -41.1238,
  -41.1441,
  -41.1648,
  -41.1851,
  -41.2043,
  -41.2221,
  -41.2383,
  -41.2535,
  -41.2678,
  -41.2822,
  -41.2973,
  -41.3131,
  -41.3297,
  -41.3466,
  -41.3635,
  -41.3799,
  -41.3956,
  -41.4103,
  -41.4223,
  -41.4331,
  -41.4411,
  -41.4467,
  -41.4507,
  -41.4541,
  -41.4577,
  -41.4615,
  -41.4659,
  -41.4703,
  -41.4745,
  -41.4778,
  -41.4793,
  -41.4786,
  -41.4755,
  -41.4701,
  -41.4624,
  -41.4519,
  -41.4389,
  -41.4238,
  -41.4069,
  -41.3895,
  -41.3718,
  -41.3536,
  -41.3339,
  -41.3118,
  -41.2865,
  -41.2573,
  -41.225,
  -41.1894,
  -41.1497,
  -41.106,
  -41.058,
  -41.0043,
  -40.9449,
  -40.8793,
  -40.8074,
  -40.7282,
  -40.6405,
  -40.5426,
  -40.4335,
  -40.3131,
  -40.1831,
  -40.047,
  -34.9288,
  -34.9678,
  -35.0065,
  -35.0473,
  -35.0894,
  -35.1327,
  -35.1771,
  -35.2214,
  -35.2654,
  -35.3082,
  -35.3498,
  -35.3903,
  -35.4299,
  -35.4693,
  -35.5081,
  -35.5467,
  -35.5851,
  -35.6224,
  -35.6604,
  -35.6983,
  -35.7359,
  -35.7737,
  -35.8116,
  -35.8496,
  -35.8878,
  -35.9258,
  -35.964,
  -36.0021,
  -36.0405,
  -36.0788,
  -36.1167,
  -36.1532,
  -36.1901,
  -36.2263,
  -36.2628,
  -36.3005,
  -36.3396,
  -36.3804,
  -36.4221,
  -36.464,
  -36.5057,
  -36.5466,
  -36.5864,
  -36.6252,
  -36.6632,
  -36.7009,
  -36.7388,
  -36.776,
  -36.8149,
  -36.8546,
  -36.8948,
  -36.9349,
  -36.9746,
  -37.0135,
  -37.0513,
  -37.088,
  -37.1237,
  -37.1589,
  -37.1939,
  -37.229,
  -37.2647,
  -37.3012,
  -37.3384,
  -37.3756,
  -37.4149,
  -37.4556,
  -37.4973,
  -37.5398,
  -37.5826,
  -37.6257,
  -37.6689,
  -37.7118,
  -37.7538,
  -37.7946,
  -37.8341,
  -37.8729,
  -37.911,
  -37.9488,
  -37.9863,
  -38.024,
  -38.0618,
  -38.099,
  -38.1372,
  -38.1757,
  -38.2141,
  -38.2521,
  -38.2898,
  -38.3266,
  -38.3624,
  -38.3971,
  -38.4311,
  -38.4647,
  -38.4982,
  -38.5316,
  -38.5651,
  -38.5988,
  -38.633,
  -38.6677,
  -38.7031,
  -38.7376,
  -38.7729,
  -38.8067,
  -38.8387,
  -38.8688,
  -38.8971,
  -38.9242,
  -38.9503,
  -38.9754,
  -38.9991,
  -39.0212,
  -39.0419,
  -39.0612,
  -39.0793,
  -39.0965,
  -39.1128,
  -39.1281,
  -39.1423,
  -39.1552,
  -39.1668,
  -39.1794,
  -39.1919,
  -39.2046,
  -39.2168,
  -39.2287,
  -39.2398,
  -39.2503,
  -39.2605,
  -39.2703,
  -39.2801,
  -39.29,
  -39.3003,
  -39.3113,
  -39.3232,
  -39.3369,
  -39.3524,
  -39.3702,
  -39.3898,
  -39.4107,
  -39.4312,
  -39.453,
  -39.4747,
  -39.4965,
  -39.5186,
  -39.5409,
  -39.5635,
  -39.5863,
  -39.6087,
  -39.6308,
  -39.6519,
  -39.6719,
  -39.6907,
  -39.7088,
  -39.726,
  -39.7427,
  -39.7589,
  -39.7747,
  -39.7902,
  -39.8054,
  -39.8204,
  -39.8352,
  -39.85,
  -39.864,
  -39.8793,
  -39.895,
  -39.9113,
  -39.928,
  -39.945,
  -39.9625,
  -39.9798,
  -39.9966,
  -40.0125,
  -40.0274,
  -40.0411,
  -40.0537,
  -40.0657,
  -40.0777,
  -40.0905,
  -40.1048,
  -40.1212,
  -40.1398,
  -40.1614,
  -40.1855,
  -40.2124,
  -40.2412,
  -40.2715,
  -40.3012,
  -40.332,
  -40.3624,
  -40.3924,
  -40.4219,
  -40.451,
  -40.4797,
  -40.5079,
  -40.5354,
  -40.5616,
  -40.5868,
  -40.6106,
  -40.6328,
  -40.6535,
  -40.6728,
  -40.69,
  -40.7049,
  -40.7174,
  -40.7272,
  -40.7348,
  -40.7405,
  -40.7443,
  -40.7464,
  -40.7474,
  -40.7478,
  -40.7484,
  -40.7495,
  -40.751,
  -40.7521,
  -40.7552,
  -40.7591,
  -40.7645,
  -40.7709,
  -40.7784,
  -40.7864,
  -40.7953,
  -40.8043,
  -40.8136,
  -40.8232,
  -40.8334,
  -40.8446,
  -40.8567,
  -40.8698,
  -40.8835,
  -40.898,
  -40.9131,
  -40.9284,
  -40.9437,
  -40.959,
  -40.9743,
  -40.9898,
  -41.0062,
  -41.0239,
  -41.0431,
  -41.0636,
  -41.0848,
  -41.1066,
  -41.1278,
  -41.1476,
  -41.1657,
  -41.1812,
  -41.1965,
  -41.211,
  -41.2255,
  -41.2405,
  -41.2562,
  -41.2724,
  -41.2889,
  -41.3052,
  -41.321,
  -41.3362,
  -41.3507,
  -41.3639,
  -41.3754,
  -41.3845,
  -41.3913,
  -41.3966,
  -41.401,
  -41.4054,
  -41.41,
  -41.4148,
  -41.4198,
  -41.4243,
  -41.428,
  -41.4299,
  -41.4297,
  -41.4274,
  -41.423,
  -41.4162,
  -41.407,
  -41.3951,
  -41.3811,
  -41.3657,
  -41.3497,
  -41.3336,
  -41.3167,
  -41.2982,
  -41.2771,
  -41.2527,
  -41.2248,
  -41.1926,
  -41.158,
  -41.1196,
  -41.0766,
  -41.0289,
  -40.9759,
  -40.9174,
  -40.8533,
  -40.7827,
  -40.7052,
  -40.6194,
  -40.5237,
  -40.4169,
  -40.2987,
  -40.1706,
  -40.036,
  -34.7974,
  -34.8369,
  -34.877,
  -34.9181,
  -34.9602,
  -35.0034,
  -35.0473,
  -35.091,
  -35.1344,
  -35.1767,
  -35.2182,
  -35.2589,
  -35.2981,
  -35.3375,
  -35.3766,
  -35.4152,
  -35.4533,
  -35.4911,
  -35.5288,
  -35.5663,
  -35.604,
  -35.6415,
  -35.679,
  -35.717,
  -35.7553,
  -35.7937,
  -35.8331,
  -35.8718,
  -35.9116,
  -35.9512,
  -35.9909,
  -36.0293,
  -36.0667,
  -36.1032,
  -36.1398,
  -36.1772,
  -36.2167,
  -36.2575,
  -36.2994,
  -36.3413,
  -36.3831,
  -36.4241,
  -36.4632,
  -36.5024,
  -36.5409,
  -36.5792,
  -36.6174,
  -36.656,
  -36.6954,
  -36.7355,
  -36.7761,
  -36.8166,
  -36.8567,
  -36.896,
  -36.9341,
  -36.9711,
  -37.0072,
  -37.0427,
  -37.0771,
  -37.1124,
  -37.1484,
  -37.1849,
  -37.2223,
  -37.2608,
  -37.3007,
  -37.3418,
  -37.3839,
  -37.4266,
  -37.4695,
  -37.5124,
  -37.5553,
  -37.5983,
  -37.6406,
  -37.6818,
  -37.7223,
  -37.761,
  -37.8001,
  -37.8389,
  -37.8775,
  -37.9163,
  -37.9551,
  -37.9943,
  -38.0336,
  -38.0732,
  -38.1127,
  -38.1517,
  -38.19,
  -38.2272,
  -38.2632,
  -38.2982,
  -38.3325,
  -38.3664,
  -38.4001,
  -38.433,
  -38.4668,
  -38.5007,
  -38.535,
  -38.5703,
  -38.6062,
  -38.6421,
  -38.6774,
  -38.7111,
  -38.7431,
  -38.773,
  -38.8011,
  -38.8282,
  -38.8545,
  -38.8797,
  -38.9037,
  -38.9262,
  -38.9473,
  -38.966,
  -38.9847,
  -39.0024,
  -39.0192,
  -39.0351,
  -39.0493,
  -39.0629,
  -39.0757,
  -39.0882,
  -39.1008,
  -39.1131,
  -39.1255,
  -39.1376,
  -39.1494,
  -39.1608,
  -39.1719,
  -39.1825,
  -39.1931,
  -39.2035,
  -39.214,
  -39.2245,
  -39.2367,
  -39.2509,
  -39.267,
  -39.2855,
  -39.306,
  -39.3277,
  -39.3498,
  -39.3722,
  -39.3944,
  -39.4168,
  -39.4394,
  -39.462,
  -39.4848,
  -39.5078,
  -39.5306,
  -39.5528,
  -39.574,
  -39.594,
  -39.6127,
  -39.6306,
  -39.6476,
  -39.6631,
  -39.6791,
  -39.6948,
  -39.7103,
  -39.7257,
  -39.7409,
  -39.7559,
  -39.7711,
  -39.7863,
  -39.8017,
  -39.8179,
  -39.8343,
  -39.8513,
  -39.8685,
  -39.886,
  -39.9028,
  -39.9195,
  -39.9354,
  -39.9503,
  -39.9642,
  -39.9775,
  -39.9905,
  -40.0037,
  -40.0176,
  -40.0322,
  -40.0497,
  -40.0697,
  -40.092,
  -40.1168,
  -40.1442,
  -40.173,
  -40.2033,
  -40.2338,
  -40.2644,
  -40.2945,
  -40.324,
  -40.3532,
  -40.3821,
  -40.4107,
  -40.4388,
  -40.4663,
  -40.4925,
  -40.517,
  -40.5404,
  -40.5622,
  -40.5825,
  -40.6012,
  -40.6183,
  -40.6334,
  -40.6465,
  -40.6563,
  -40.6649,
  -40.6714,
  -40.6759,
  -40.6787,
  -40.6802,
  -40.6808,
  -40.6814,
  -40.682,
  -40.683,
  -40.6846,
  -40.6869,
  -40.6905,
  -40.6957,
  -40.7023,
  -40.7101,
  -40.7182,
  -40.727,
  -40.7351,
  -40.7437,
  -40.753,
  -40.7632,
  -40.7746,
  -40.7875,
  -40.8015,
  -40.8164,
  -40.832,
  -40.8479,
  -40.8638,
  -40.8796,
  -40.8953,
  -40.9101,
  -40.9264,
  -40.9437,
  -40.9624,
  -40.9829,
  -41.0043,
  -41.0266,
  -41.049,
  -41.0706,
  -41.0907,
  -41.109,
  -41.1257,
  -41.1412,
  -41.156,
  -41.1706,
  -41.1856,
  -41.2011,
  -41.2169,
  -41.2329,
  -41.2485,
  -41.2635,
  -41.278,
  -41.2921,
  -41.3054,
  -41.3176,
  -41.3278,
  -41.336,
  -41.3427,
  -41.3488,
  -41.3543,
  -41.3596,
  -41.3651,
  -41.3703,
  -41.3748,
  -41.3783,
  -41.3805,
  -41.3807,
  -41.3778,
  -41.3744,
  -41.3689,
  -41.361,
  -41.3507,
  -41.3381,
  -41.3242,
  -41.3096,
  -41.2947,
  -41.2791,
  -41.2616,
  -41.2416,
  -41.2185,
  -41.192,
  -41.1621,
  -41.1287,
  -41.0913,
  -41.0493,
  -41.0022,
  -40.9498,
  -40.8921,
  -40.8291,
  -40.7603,
  -40.6844,
  -40.6006,
  -40.5073,
  -40.4031,
  -40.288,
  -40.1628,
  -40.0308,
  -34.6679,
  -34.708,
  -34.7484,
  -34.7899,
  -34.8325,
  -34.8755,
  -34.9189,
  -34.9612,
  -35.0036,
  -35.0456,
  -35.087,
  -35.1279,
  -35.1683,
  -35.2081,
  -35.2472,
  -35.2855,
  -35.3232,
  -35.3606,
  -35.3979,
  -35.4352,
  -35.4724,
  -35.5099,
  -35.5467,
  -35.5849,
  -35.6236,
  -35.6631,
  -35.7033,
  -35.7441,
  -35.7857,
  -35.8271,
  -35.8678,
  -35.9072,
  -35.9451,
  -35.9818,
  -36.0185,
  -36.0562,
  -36.0955,
  -36.1354,
  -36.1771,
  -36.2191,
  -36.2607,
  -36.3018,
  -36.3422,
  -36.382,
  -36.4211,
  -36.4599,
  -36.4986,
  -36.5376,
  -36.5774,
  -36.6176,
  -36.6585,
  -36.6994,
  -36.74,
  -36.7785,
  -36.8169,
  -36.8541,
  -36.8906,
  -36.9267,
  -36.9626,
  -36.9985,
  -37.0348,
  -37.0715,
  -37.1092,
  -37.1481,
  -37.1884,
  -37.2299,
  -37.2723,
  -37.315,
  -37.3578,
  -37.3994,
  -37.4421,
  -37.4848,
  -37.5272,
  -37.569,
  -37.6102,
  -37.6508,
  -37.6911,
  -37.7309,
  -37.7705,
  -37.8103,
  -37.8503,
  -37.8907,
  -37.9312,
  -37.9721,
  -38.0125,
  -38.0523,
  -38.0911,
  -38.1277,
  -38.164,
  -38.1991,
  -38.2337,
  -38.2679,
  -38.3021,
  -38.3366,
  -38.3709,
  -38.4055,
  -38.4403,
  -38.476,
  -38.5122,
  -38.5483,
  -38.5834,
  -38.6168,
  -38.6483,
  -38.6776,
  -38.7054,
  -38.7313,
  -38.7573,
  -38.7827,
  -38.8069,
  -38.8297,
  -38.8513,
  -38.8718,
  -38.8913,
  -38.9097,
  -38.9272,
  -38.9433,
  -38.9582,
  -38.9721,
  -38.9852,
  -38.9977,
  -39.0101,
  -39.0223,
  -39.0346,
  -39.047,
  -39.0596,
  -39.0709,
  -39.083,
  -39.0945,
  -39.1057,
  -39.1164,
  -39.1275,
  -39.1392,
  -39.1521,
  -39.1666,
  -39.1834,
  -39.2027,
  -39.224,
  -39.2463,
  -39.269,
  -39.2919,
  -39.3148,
  -39.3379,
  -39.3609,
  -39.3842,
  -39.4075,
  -39.4308,
  -39.4528,
  -39.4751,
  -39.4963,
  -39.5161,
  -39.5345,
  -39.5518,
  -39.5684,
  -39.5845,
  -39.6003,
  -39.6159,
  -39.6316,
  -39.6473,
  -39.6628,
  -39.6783,
  -39.6939,
  -39.7094,
  -39.7254,
  -39.7416,
  -39.7583,
  -39.7754,
  -39.7926,
  -39.8096,
  -39.8263,
  -39.8417,
  -39.8573,
  -39.8721,
  -39.8866,
  -39.9006,
  -39.915,
  -39.9299,
  -39.9458,
  -39.9633,
  -39.9826,
  -40.0038,
  -40.0275,
  -40.053,
  -40.0804,
  -40.1092,
  -40.1392,
  -40.1694,
  -40.1994,
  -40.2292,
  -40.2581,
  -40.2868,
  -40.3152,
  -40.3435,
  -40.3715,
  -40.3988,
  -40.4239,
  -40.4484,
  -40.4713,
  -40.4925,
  -40.5121,
  -40.5302,
  -40.5468,
  -40.5621,
  -40.5754,
  -40.587,
  -40.5963,
  -40.6037,
  -40.609,
  -40.6124,
  -40.6142,
  -40.6152,
  -40.6156,
  -40.616,
  -40.6166,
  -40.6174,
  -40.6191,
  -40.6223,
  -40.6273,
  -40.6339,
  -40.6416,
  -40.65,
  -40.6581,
  -40.6662,
  -40.6746,
  -40.6823,
  -40.6922,
  -40.7039,
  -40.7171,
  -40.7319,
  -40.7479,
  -40.7645,
  -40.7815,
  -40.7984,
  -40.815,
  -40.8315,
  -40.8482,
  -40.8657,
  -40.8842,
  -40.9042,
  -40.9257,
  -40.9482,
  -40.9712,
  -40.9938,
  -41.0155,
  -41.0356,
  -41.0539,
  -41.0707,
  -41.0865,
  -41.1017,
  -41.1167,
  -41.1317,
  -41.1471,
  -41.1627,
  -41.1779,
  -41.1929,
  -41.2073,
  -41.2211,
  -41.2348,
  -41.2481,
  -41.2598,
  -41.2709,
  -41.2804,
  -41.2884,
  -41.2959,
  -41.3026,
  -41.309,
  -41.3148,
  -41.32,
  -41.3243,
  -41.3278,
  -41.3298,
  -41.3303,
  -41.3293,
  -41.3267,
  -41.3226,
  -41.3165,
  -41.3078,
  -41.2969,
  -41.2845,
  -41.2711,
  -41.2573,
  -41.2426,
  -41.2263,
  -41.2074,
  -41.1855,
  -41.1603,
  -41.132,
  -41.1,
  -41.0638,
  -41.0229,
  -40.9765,
  -40.9246,
  -40.8675,
  -40.8055,
  -40.7379,
  -40.6638,
  -40.5817,
  -40.4907,
  -40.3898,
  -40.278,
  -40.1567,
  -40.0285,
  -34.5392,
  -34.5797,
  -34.6197,
  -34.6616,
  -34.7046,
  -34.7477,
  -34.7907,
  -34.8332,
  -34.8751,
  -34.9167,
  -34.9579,
  -34.9989,
  -35.0395,
  -35.0793,
  -35.1183,
  -35.1563,
  -35.1936,
  -35.2295,
  -35.2664,
  -35.3035,
  -35.3408,
  -35.3786,
  -35.4168,
  -35.4555,
  -35.495,
  -35.5355,
  -35.577,
  -35.6193,
  -35.6621,
  -35.7047,
  -35.7462,
  -35.7863,
  -35.8236,
  -35.8605,
  -35.8972,
  -35.9352,
  -35.9746,
  -36.0153,
  -36.0568,
  -36.0984,
  -36.1399,
  -36.1812,
  -36.2221,
  -36.2625,
  -36.3023,
  -36.3415,
  -36.3806,
  -36.419,
  -36.4589,
  -36.4994,
  -36.5405,
  -36.5819,
  -36.6228,
  -36.6626,
  -36.7012,
  -36.7387,
  -36.7756,
  -36.8124,
  -36.8491,
  -36.8858,
  -36.9227,
  -36.9599,
  -36.998,
  -37.0374,
  -37.077,
  -37.1189,
  -37.1614,
  -37.2041,
  -37.2464,
  -37.2888,
  -37.3312,
  -37.3737,
  -37.4162,
  -37.4586,
  -37.5006,
  -37.5421,
  -37.5831,
  -37.6239,
  -37.6646,
  -37.7054,
  -37.7467,
  -37.7874,
  -37.8292,
  -37.871,
  -37.9123,
  -37.9528,
  -37.9922,
  -38.0299,
  -38.0663,
  -38.1016,
  -38.1364,
  -38.1712,
  -38.206,
  -38.241,
  -38.276,
  -38.3115,
  -38.3474,
  -38.3836,
  -38.4201,
  -38.4551,
  -38.49,
  -38.5228,
  -38.5534,
  -38.5819,
  -38.6091,
  -38.6358,
  -38.6616,
  -38.6868,
  -38.7112,
  -38.7346,
  -38.7567,
  -38.7781,
  -38.7987,
  -38.818,
  -38.8362,
  -38.8529,
  -38.8681,
  -38.8822,
  -38.8945,
  -38.907,
  -38.9192,
  -38.9314,
  -38.9439,
  -38.9567,
  -38.9699,
  -38.9833,
  -38.9963,
  -39.0088,
  -39.0205,
  -39.0318,
  -39.0431,
  -39.055,
  -39.0682,
  -39.0833,
  -39.1008,
  -39.1207,
  -39.1425,
  -39.1654,
  -39.1887,
  -39.2113,
  -39.2348,
  -39.2585,
  -39.2824,
  -39.3064,
  -39.3304,
  -39.3541,
  -39.3773,
  -39.3998,
  -39.4207,
  -39.4402,
  -39.4581,
  -39.4746,
  -39.4906,
  -39.5061,
  -39.5216,
  -39.5374,
  -39.5534,
  -39.5695,
  -39.5856,
  -39.6015,
  -39.6176,
  -39.6326,
  -39.6487,
  -39.6651,
  -39.682,
  -39.699,
  -39.7162,
  -39.7329,
  -39.7492,
  -39.7652,
  -39.7806,
  -39.7958,
  -39.8109,
  -39.8261,
  -39.8419,
  -39.8588,
  -39.8768,
  -39.8964,
  -39.9177,
  -39.9406,
  -39.9649,
  -39.9911,
  -40.0187,
  -40.0474,
  -40.0767,
  -40.1065,
  -40.1348,
  -40.1639,
  -40.1924,
  -40.2205,
  -40.2485,
  -40.2766,
  -40.3044,
  -40.3314,
  -40.3574,
  -40.3819,
  -40.4046,
  -40.4253,
  -40.4443,
  -40.4617,
  -40.478,
  -40.4929,
  -40.5066,
  -40.5186,
  -40.5287,
  -40.5369,
  -40.5429,
  -40.5469,
  -40.5492,
  -40.5502,
  -40.5506,
  -40.5507,
  -40.5508,
  -40.5501,
  -40.5514,
  -40.5542,
  -40.559,
  -40.5654,
  -40.5729,
  -40.5809,
  -40.5889,
  -40.5966,
  -40.6045,
  -40.6132,
  -40.6227,
  -40.6343,
  -40.6478,
  -40.6632,
  -40.68,
  -40.6979,
  -40.716,
  -40.7341,
  -40.7519,
  -40.7696,
  -40.7875,
  -40.8063,
  -40.8265,
  -40.8478,
  -40.8704,
  -40.8938,
  -40.9172,
  -40.94,
  -40.9615,
  -40.9813,
  -40.9996,
  -41.0155,
  -41.0315,
  -41.0471,
  -41.0625,
  -41.0778,
  -41.0931,
  -41.1083,
  -41.1234,
  -41.138,
  -41.1517,
  -41.165,
  -41.1783,
  -41.1915,
  -41.2042,
  -41.216,
  -41.2267,
  -41.2361,
  -41.2448,
  -41.2526,
  -41.2596,
  -41.2657,
  -41.2707,
  -41.2747,
  -41.2778,
  -41.2798,
  -41.2806,
  -41.2809,
  -41.2798,
  -41.2771,
  -41.2725,
  -41.2656,
  -41.2563,
  -41.2453,
  -41.2331,
  -41.2203,
  -41.2065,
  -41.1912,
  -41.1734,
  -41.1526,
  -41.1291,
  -41.1021,
  -41.0704,
  -41.0356,
  -40.9954,
  -40.9498,
  -40.8983,
  -40.8416,
  -40.7801,
  -40.7136,
  -40.641,
  -40.5606,
  -40.4719,
  -40.3738,
  -40.2659,
  -40.1487,
  -40.0248,
  -34.4102,
  -34.4511,
  -34.4926,
  -34.535,
  -34.5781,
  -34.6213,
  -34.6641,
  -34.7062,
  -34.7477,
  -34.7888,
  -34.8298,
  -34.8706,
  -34.9101,
  -34.9497,
  -34.9886,
  -35.0263,
  -35.0634,
  -35.1001,
  -35.1369,
  -35.174,
  -35.2116,
  -35.2498,
  -35.2888,
  -35.3285,
  -35.3691,
  -35.4109,
  -35.4536,
  -35.4961,
  -35.54,
  -35.5834,
  -35.6254,
  -35.6656,
  -35.7039,
  -35.7411,
  -35.7779,
  -35.8158,
  -35.8551,
  -35.8956,
  -35.9368,
  -35.9782,
  -36.0196,
  -36.0611,
  -36.1017,
  -36.1428,
  -36.1833,
  -36.2231,
  -36.2624,
  -36.3019,
  -36.342,
  -36.3828,
  -36.4243,
  -36.4659,
  -36.5071,
  -36.5471,
  -36.5859,
  -36.6237,
  -36.6612,
  -36.6988,
  -36.7355,
  -36.7732,
  -36.8109,
  -36.8489,
  -36.8876,
  -36.9274,
  -36.9685,
  -37.0106,
  -37.0531,
  -37.0955,
  -37.1376,
  -37.1797,
  -37.2219,
  -37.2645,
  -37.3074,
  -37.3504,
  -37.3931,
  -37.4342,
  -37.4761,
  -37.5176,
  -37.5592,
  -37.6012,
  -37.6435,
  -37.6863,
  -37.7292,
  -37.7718,
  -37.8139,
  -37.855,
  -37.8945,
  -37.9325,
  -37.9691,
  -38.0047,
  -38.04,
  -38.0752,
  -38.1107,
  -38.1455,
  -38.1814,
  -38.2177,
  -38.2544,
  -38.2913,
  -38.3281,
  -38.364,
  -38.3984,
  -38.4305,
  -38.4602,
  -38.488,
  -38.5146,
  -38.5406,
  -38.5662,
  -38.5917,
  -38.616,
  -38.6399,
  -38.6633,
  -38.6857,
  -38.7063,
  -38.727,
  -38.7456,
  -38.7629,
  -38.7786,
  -38.7928,
  -38.806,
  -38.8186,
  -38.8308,
  -38.8429,
  -38.8555,
  -38.8688,
  -38.8829,
  -38.8972,
  -38.9112,
  -38.9244,
  -38.9365,
  -38.9481,
  -38.9597,
  -38.972,
  -38.9846,
  -39.0002,
  -39.0183,
  -39.0388,
  -39.061,
  -39.0843,
  -39.1081,
  -39.132,
  -39.1564,
  -39.1809,
  -39.2055,
  -39.2302,
  -39.2548,
  -39.2793,
  -39.3029,
  -39.3252,
  -39.346,
  -39.3649,
  -39.3821,
  -39.398,
  -39.4132,
  -39.4273,
  -39.4428,
  -39.4587,
  -39.4751,
  -39.4917,
  -39.5085,
  -39.5252,
  -39.5416,
  -39.5579,
  -39.5742,
  -39.5906,
  -39.6073,
  -39.6241,
  -39.6409,
  -39.6574,
  -39.6737,
  -39.6895,
  -39.705,
  -39.7207,
  -39.7364,
  -39.7528,
  -39.7703,
  -39.7892,
  -39.8095,
  -39.8302,
  -39.8534,
  -39.8778,
  -39.9034,
  -39.93,
  -39.9576,
  -39.986,
  -40.0149,
  -40.0438,
  -40.0726,
  -40.1011,
  -40.129,
  -40.1565,
  -40.1841,
  -40.2118,
  -40.2393,
  -40.2663,
  -40.2923,
  -40.3168,
  -40.3391,
  -40.3596,
  -40.3779,
  -40.3949,
  -40.4106,
  -40.4254,
  -40.439,
  -40.4516,
  -40.4615,
  -40.4705,
  -40.4772,
  -40.4817,
  -40.4844,
  -40.4854,
  -40.4857,
  -40.4855,
  -40.4852,
  -40.4853,
  -40.4863,
  -40.489,
  -40.4936,
  -40.4996,
  -40.5065,
  -40.5137,
  -40.521,
  -40.5283,
  -40.5359,
  -40.5441,
  -40.5537,
  -40.5654,
  -40.5791,
  -40.595,
  -40.6127,
  -40.6315,
  -40.6509,
  -40.6703,
  -40.6895,
  -40.7086,
  -40.7271,
  -40.7474,
  -40.7689,
  -40.7915,
  -40.8152,
  -40.8394,
  -40.8632,
  -40.8861,
  -40.9073,
  -40.9271,
  -40.9452,
  -40.9621,
  -40.9784,
  -40.9944,
  -41.0101,
  -41.0256,
  -41.041,
  -41.0562,
  -41.0711,
  -41.0855,
  -41.099,
  -41.1119,
  -41.1248,
  -41.1376,
  -41.1504,
  -41.1626,
  -41.174,
  -41.1845,
  -41.194,
  -41.2026,
  -41.21,
  -41.2161,
  -41.221,
  -41.2248,
  -41.2278,
  -41.2302,
  -41.232,
  -41.2322,
  -41.2325,
  -41.2315,
  -41.2284,
  -41.223,
  -41.2151,
  -41.2053,
  -41.1942,
  -41.1824,
  -41.1696,
  -41.1552,
  -41.1386,
  -41.1193,
  -41.097,
  -41.0714,
  -41.0419,
  -41.0082,
  -40.9688,
  -40.9237,
  -40.8725,
  -40.816,
  -40.7546,
  -40.6887,
  -40.6172,
  -40.5387,
  -40.4521,
  -40.3566,
  -40.2523,
  -40.1396,
  -40.0205,
  -34.2828,
  -34.3242,
  -34.3661,
  -34.4088,
  -34.452,
  -34.4953,
  -34.5381,
  -34.579,
  -34.6202,
  -34.661,
  -34.7016,
  -34.7421,
  -34.7822,
  -34.8217,
  -34.8602,
  -34.898,
  -34.935,
  -34.9718,
  -35.0087,
  -35.0461,
  -35.0842,
  -35.1232,
  -35.1622,
  -35.2032,
  -35.2452,
  -35.2882,
  -35.3321,
  -35.3766,
  -35.421,
  -35.4646,
  -35.5066,
  -35.5467,
  -35.585,
  -35.6222,
  -35.6592,
  -35.6971,
  -35.7361,
  -35.7753,
  -35.8162,
  -35.8575,
  -35.8991,
  -35.941,
  -35.9831,
  -36.0249,
  -36.0659,
  -36.1062,
  -36.1459,
  -36.1856,
  -36.2258,
  -36.2668,
  -36.3085,
  -36.3505,
  -36.392,
  -36.4313,
  -36.4703,
  -36.5085,
  -36.5467,
  -36.5851,
  -36.6238,
  -36.6626,
  -36.7012,
  -36.74,
  -36.7794,
  -36.8197,
  -36.8611,
  -36.9034,
  -36.9458,
  -36.9881,
  -37.03,
  -37.0721,
  -37.1136,
  -37.1565,
  -37.1999,
  -37.2434,
  -37.2868,
  -37.3297,
  -37.3721,
  -37.4144,
  -37.4569,
  -37.4998,
  -37.5431,
  -37.5868,
  -37.6305,
  -37.6738,
  -37.7163,
  -37.7575,
  -37.7972,
  -37.8344,
  -37.8713,
  -37.9072,
  -37.9429,
  -37.9789,
  -38.0152,
  -38.0519,
  -38.0888,
  -38.1259,
  -38.1631,
  -38.2004,
  -38.2373,
  -38.2731,
  -38.3069,
  -38.3384,
  -38.3674,
  -38.3947,
  -38.4208,
  -38.4455,
  -38.4709,
  -38.4962,
  -38.5212,
  -38.5457,
  -38.5699,
  -38.5934,
  -38.616,
  -38.6373,
  -38.6569,
  -38.6748,
  -38.6907,
  -38.7052,
  -38.7184,
  -38.731,
  -38.7432,
  -38.7556,
  -38.7687,
  -38.7827,
  -38.7974,
  -38.8115,
  -38.8261,
  -38.8399,
  -38.8527,
  -38.8647,
  -38.8767,
  -38.8895,
  -38.9037,
  -38.9198,
  -38.9383,
  -38.9591,
  -38.9814,
  -39.0048,
  -39.0289,
  -39.0534,
  -39.0783,
  -39.1034,
  -39.1287,
  -39.1542,
  -39.1794,
  -39.2041,
  -39.2271,
  -39.2495,
  -39.2701,
  -39.2888,
  -39.3055,
  -39.3208,
  -39.3355,
  -39.3505,
  -39.366,
  -39.3822,
  -39.399,
  -39.4162,
  -39.4336,
  -39.4508,
  -39.4678,
  -39.4844,
  -39.5009,
  -39.5172,
  -39.5337,
  -39.5501,
  -39.5667,
  -39.583,
  -39.5992,
  -39.6142,
  -39.6301,
  -39.6461,
  -39.6628,
  -39.6802,
  -39.6991,
  -39.7197,
  -39.7418,
  -39.7655,
  -39.7904,
  -39.8163,
  -39.8428,
  -39.87,
  -39.8977,
  -39.9259,
  -39.9543,
  -39.9827,
  -40.0109,
  -40.0388,
  -40.0662,
  -40.0935,
  -40.1207,
  -40.1481,
  -40.1754,
  -40.2024,
  -40.2283,
  -40.2516,
  -40.2739,
  -40.294,
  -40.3119,
  -40.3283,
  -40.3438,
  -40.3583,
  -40.3723,
  -40.3853,
  -40.3968,
  -40.4066,
  -40.414,
  -40.4191,
  -40.4218,
  -40.423,
  -40.4231,
  -40.4228,
  -40.4223,
  -40.4224,
  -40.4235,
  -40.4261,
  -40.4303,
  -40.4356,
  -40.4416,
  -40.4477,
  -40.454,
  -40.4605,
  -40.4676,
  -40.4757,
  -40.4845,
  -40.4964,
  -40.5106,
  -40.5271,
  -40.5455,
  -40.5653,
  -40.5858,
  -40.6066,
  -40.6272,
  -40.6478,
  -40.6687,
  -40.6904,
  -40.7133,
  -40.7371,
  -40.7617,
  -40.7864,
  -40.8107,
  -40.8337,
  -40.8552,
  -40.875,
  -40.8931,
  -40.9102,
  -40.9266,
  -40.9427,
  -40.9586,
  -40.9742,
  -40.9897,
  -41.0049,
  -41.0198,
  -41.0341,
  -41.0476,
  -41.0605,
  -41.0731,
  -41.0857,
  -41.0972,
  -41.1095,
  -41.1213,
  -41.1323,
  -41.1423,
  -41.1512,
  -41.1587,
  -41.1648,
  -41.1696,
  -41.1735,
  -41.1768,
  -41.1798,
  -41.1828,
  -41.1854,
  -41.1873,
  -41.1878,
  -41.1861,
  -41.1819,
  -41.1752,
  -41.1663,
  -41.1562,
  -41.1453,
  -41.1336,
  -41.1203,
  -41.1049,
  -41.087,
  -41.066,
  -41.0418,
  -41.0135,
  -40.9803,
  -40.9417,
  -40.8966,
  -40.8456,
  -40.7891,
  -40.7278,
  -40.6618,
  -40.591,
  -40.5142,
  -40.4298,
  -40.337,
  -40.236,
  -40.1274,
  -40.0128,
  -34.1566,
  -34.1983,
  -34.2405,
  -34.2824,
  -34.3257,
  -34.369,
  -34.4117,
  -34.4535,
  -34.4947,
  -34.5353,
  -34.5756,
  -34.6158,
  -34.6553,
  -34.6945,
  -34.7327,
  -34.7707,
  -34.808,
  -34.8443,
  -34.8815,
  -34.9193,
  -34.9581,
  -34.9982,
  -35.0396,
  -35.0821,
  -35.1254,
  -35.1697,
  -35.2144,
  -35.2595,
  -35.3039,
  -35.3471,
  -35.3886,
  -35.4285,
  -35.4657,
  -35.503,
  -35.5402,
  -35.5781,
  -35.617,
  -35.6569,
  -35.6977,
  -35.7391,
  -35.7809,
  -35.8231,
  -35.8655,
  -35.9076,
  -35.949,
  -35.9897,
  -36.0299,
  -36.0701,
  -36.1096,
  -36.1511,
  -36.193,
  -36.2352,
  -36.277,
  -36.3174,
  -36.3568,
  -36.3957,
  -36.4345,
  -36.4739,
  -36.5134,
  -36.553,
  -36.5925,
  -36.6321,
  -36.6721,
  -36.7128,
  -36.7535,
  -36.7958,
  -36.8381,
  -36.8803,
  -36.9223,
  -36.9649,
  -37.008,
  -37.0518,
  -37.096,
  -37.1404,
  -37.1843,
  -37.2278,
  -37.2707,
  -37.3134,
  -37.3566,
  -37.4003,
  -37.4445,
  -37.4879,
  -37.5321,
  -37.5758,
  -37.6184,
  -37.6597,
  -37.6995,
  -37.7377,
  -37.7747,
  -37.8111,
  -37.8475,
  -37.8843,
  -37.9218,
  -37.9595,
  -37.997,
  -38.0348,
  -38.0722,
  -38.1097,
  -38.1464,
  -38.1809,
  -38.2143,
  -38.2453,
  -38.274,
  -38.301,
  -38.3271,
  -38.3531,
  -38.3787,
  -38.4041,
  -38.4295,
  -38.4547,
  -38.4794,
  -38.5038,
  -38.5272,
  -38.5493,
  -38.5694,
  -38.5875,
  -38.6039,
  -38.6184,
  -38.6309,
  -38.6435,
  -38.6559,
  -38.6688,
  -38.6825,
  -38.6973,
  -38.7127,
  -38.7283,
  -38.7435,
  -38.7576,
  -38.7708,
  -38.7833,
  -38.796,
  -38.8094,
  -38.8242,
  -38.841,
  -38.8597,
  -38.8803,
  -38.9025,
  -38.9258,
  -38.95,
  -38.9739,
  -38.9992,
  -39.0249,
  -39.0507,
  -39.0766,
  -39.1023,
  -39.1274,
  -39.1514,
  -39.174,
  -39.195,
  -39.2135,
  -39.2299,
  -39.2452,
  -39.2599,
  -39.2749,
  -39.2906,
  -39.3071,
  -39.3245,
  -39.3421,
  -39.36,
  -39.3777,
  -39.395,
  -39.4108,
  -39.4273,
  -39.4437,
  -39.46,
  -39.4763,
  -39.4927,
  -39.509,
  -39.5254,
  -39.5417,
  -39.5582,
  -39.5749,
  -39.5922,
  -39.6106,
  -39.6305,
  -39.6522,
  -39.6757,
  -39.7008,
  -39.7271,
  -39.7542,
  -39.7818,
  -39.8095,
  -39.8375,
  -39.8655,
  -39.8937,
  -39.9217,
  -39.9485,
  -39.9761,
  -40.0033,
  -40.0303,
  -40.0575,
  -40.0848,
  -40.1118,
  -40.1388,
  -40.1647,
  -40.1885,
  -40.2104,
  -40.2303,
  -40.248,
  -40.264,
  -40.2794,
  -40.2939,
  -40.3081,
  -40.3215,
  -40.3338,
  -40.3444,
  -40.3525,
  -40.3577,
  -40.3606,
  -40.3615,
  -40.3615,
  -40.3612,
  -40.361,
  -40.3614,
  -40.3618,
  -40.3643,
  -40.3681,
  -40.3725,
  -40.3772,
  -40.3819,
  -40.3869,
  -40.3925,
  -40.3991,
  -40.4071,
  -40.4171,
  -40.4295,
  -40.4445,
  -40.4619,
  -40.4813,
  -40.502,
  -40.5236,
  -40.5454,
  -40.5672,
  -40.5891,
  -40.6113,
  -40.6343,
  -40.6583,
  -40.6831,
  -40.7083,
  -40.7336,
  -40.7583,
  -40.7817,
  -40.8037,
  -40.824,
  -40.8425,
  -40.8599,
  -40.8754,
  -40.8916,
  -40.9075,
  -40.923,
  -40.9384,
  -40.9536,
  -40.9685,
  -40.983,
  -40.9967,
  -41.0097,
  -41.0221,
  -41.0344,
  -41.0466,
  -41.0587,
  -41.0704,
  -41.0815,
  -41.0916,
  -41.1004,
  -41.1078,
  -41.1138,
  -41.1187,
  -41.1228,
  -41.1267,
  -41.1309,
  -41.1353,
  -41.1395,
  -41.143,
  -41.1449,
  -41.1444,
  -41.1412,
  -41.1353,
  -41.1273,
  -41.118,
  -41.108,
  -41.0972,
  -41.0852,
  -41.0711,
  -41.0545,
  -41.0348,
  -41.0116,
  -40.9841,
  -40.9506,
  -40.912,
  -40.8667,
  -40.8161,
  -40.7595,
  -40.6982,
  -40.6326,
  -40.5622,
  -40.4864,
  -40.4039,
  -40.3134,
  -40.2152,
  -40.11,
  -39.9997,
  -34.0312,
  -34.0733,
  -34.1157,
  -34.1585,
  -34.2016,
  -34.2449,
  -34.2875,
  -34.3294,
  -34.3706,
  -34.4113,
  -34.4515,
  -34.4914,
  -34.5297,
  -34.5684,
  -34.6066,
  -34.6445,
  -34.6821,
  -34.7195,
  -34.7575,
  -34.7961,
  -34.836,
  -34.8774,
  -34.9201,
  -34.964,
  -35.0084,
  -35.0536,
  -35.0988,
  -35.1428,
  -35.1869,
  -35.2293,
  -35.2703,
  -35.3099,
  -35.3482,
  -35.3858,
  -35.4234,
  -35.4616,
  -35.5005,
  -35.5404,
  -35.5812,
  -35.6226,
  -35.6646,
  -35.7068,
  -35.7491,
  -35.79,
  -35.8316,
  -35.8726,
  -35.9135,
  -35.9544,
  -35.996,
  -36.0378,
  -36.0799,
  -36.1225,
  -36.1642,
  -36.205,
  -36.2449,
  -36.2843,
  -36.3239,
  -36.3639,
  -36.4043,
  -36.4437,
  -36.4839,
  -36.5241,
  -36.5647,
  -36.6058,
  -36.6475,
  -36.6897,
  -36.7319,
  -36.7739,
  -36.8165,
  -36.86,
  -36.9042,
  -36.9491,
  -36.9945,
  -37.0395,
  -37.0843,
  -37.127,
  -37.1703,
  -37.2137,
  -37.2574,
  -37.3017,
  -37.3465,
  -37.3913,
  -37.4359,
  -37.4797,
  -37.5225,
  -37.5638,
  -37.6036,
  -37.6419,
  -37.6791,
  -37.716,
  -37.7531,
  -37.7908,
  -37.8292,
  -37.8667,
  -37.9053,
  -37.943,
  -37.9806,
  -38.0181,
  -38.0543,
  -38.0894,
  -38.1223,
  -38.1531,
  -38.1818,
  -38.2091,
  -38.2356,
  -38.2617,
  -38.2877,
  -38.314,
  -38.34,
  -38.3658,
  -38.3914,
  -38.4163,
  -38.4391,
  -38.4615,
  -38.482,
  -38.5005,
  -38.517,
  -38.5318,
  -38.5453,
  -38.5582,
  -38.5712,
  -38.5847,
  -38.599,
  -38.6143,
  -38.6302,
  -38.6462,
  -38.6615,
  -38.676,
  -38.6895,
  -38.7028,
  -38.7162,
  -38.7303,
  -38.7448,
  -38.7618,
  -38.7806,
  -38.801,
  -38.8229,
  -38.846,
  -38.8704,
  -38.8956,
  -38.9214,
  -38.9473,
  -38.9733,
  -38.9994,
  -39.0253,
  -39.0507,
  -39.075,
  -39.0982,
  -39.1193,
  -39.1382,
  -39.155,
  -39.1705,
  -39.1854,
  -39.2005,
  -39.2155,
  -39.2324,
  -39.2501,
  -39.268,
  -39.2859,
  -39.3039,
  -39.3213,
  -39.3384,
  -39.3553,
  -39.3718,
  -39.3881,
  -39.4043,
  -39.4206,
  -39.437,
  -39.4537,
  -39.4705,
  -39.4876,
  -39.5051,
  -39.5232,
  -39.5423,
  -39.563,
  -39.5856,
  -39.6099,
  -39.6359,
  -39.6622,
  -39.6901,
  -39.7186,
  -39.7471,
  -39.7755,
  -39.8036,
  -39.8317,
  -39.8596,
  -39.8874,
  -39.915,
  -39.9423,
  -39.9694,
  -39.9964,
  -40.0237,
  -40.0508,
  -40.0774,
  -40.1027,
  -40.1263,
  -40.1479,
  -40.1673,
  -40.185,
  -40.2012,
  -40.2166,
  -40.2317,
  -40.2462,
  -40.2601,
  -40.2718,
  -40.2828,
  -40.291,
  -40.2964,
  -40.2993,
  -40.3003,
  -40.3002,
  -40.3,
  -40.3001,
  -40.3009,
  -40.3025,
  -40.3051,
  -40.3081,
  -40.3114,
  -40.3148,
  -40.3181,
  -40.3218,
  -40.3263,
  -40.3321,
  -40.3398,
  -40.3503,
  -40.3636,
  -40.3797,
  -40.3984,
  -40.419,
  -40.441,
  -40.4635,
  -40.4863,
  -40.509,
  -40.532,
  -40.5552,
  -40.5782,
  -40.603,
  -40.6285,
  -40.6542,
  -40.68,
  -40.7053,
  -40.7296,
  -40.7524,
  -40.7734,
  -40.7925,
  -40.8103,
  -40.8271,
  -40.8431,
  -40.8588,
  -40.8742,
  -40.8893,
  -40.9044,
  -40.9193,
  -40.9338,
  -40.9476,
  -40.9607,
  -40.9731,
  -40.9852,
  -40.9971,
  -41.0089,
  -41.0203,
  -41.0311,
  -41.0408,
  -41.0493,
  -41.0564,
  -41.0624,
  -41.0675,
  -41.0723,
  -41.077,
  -41.0824,
  -41.0883,
  -41.0942,
  -41.0982,
  -41.1013,
  -41.1018,
  -41.0995,
  -41.0944,
  -41.0872,
  -41.0786,
  -41.0694,
  -41.0595,
  -41.0486,
  -41.0358,
  -41.0206,
  -41.002,
  -40.9795,
  -40.9525,
  -40.9202,
  -40.8817,
  -40.8368,
  -40.7856,
  -40.7291,
  -40.6683,
  -40.603,
  -40.5332,
  -40.458,
  -40.3767,
  -40.2886,
  -40.1931,
  -40.0911,
  -39.9841,
  -33.9089,
  -33.9511,
  -33.9938,
  -34.0367,
  -34.0796,
  -34.1224,
  -34.165,
  -34.2069,
  -34.2472,
  -34.2881,
  -34.3285,
  -34.3684,
  -34.4076,
  -34.4462,
  -34.4843,
  -34.5221,
  -34.5598,
  -34.5977,
  -34.6362,
  -34.6761,
  -34.7171,
  -34.7598,
  -34.8028,
  -34.8477,
  -34.8931,
  -34.9386,
  -34.9839,
  -35.0285,
  -35.0718,
  -35.1137,
  -35.1542,
  -35.1935,
  -35.2321,
  -35.2704,
  -35.3086,
  -35.3472,
  -35.3865,
  -35.4254,
  -35.4661,
  -35.5075,
  -35.5493,
  -35.5913,
  -35.6331,
  -35.6746,
  -35.7161,
  -35.7575,
  -35.7992,
  -35.8412,
  -35.8834,
  -35.9259,
  -35.9687,
  -36.011,
  -36.0531,
  -36.0932,
  -36.1336,
  -36.1737,
  -36.2141,
  -36.2549,
  -36.2959,
  -36.3369,
  -36.3777,
  -36.4184,
  -36.4594,
  -36.5007,
  -36.5424,
  -36.5844,
  -36.6264,
  -36.6689,
  -36.7122,
  -36.7564,
  -36.8008,
  -36.847,
  -36.8935,
  -36.9396,
  -36.9848,
  -37.0291,
  -37.0729,
  -37.1168,
  -37.161,
  -37.2057,
  -37.2508,
  -37.2959,
  -37.3406,
  -37.3846,
  -37.4275,
  -37.469,
  -37.509,
  -37.5465,
  -37.5841,
  -37.6215,
  -37.6592,
  -37.6977,
  -37.7369,
  -37.7761,
  -37.8149,
  -37.8529,
  -37.8903,
  -37.9271,
  -37.963,
  -37.9975,
  -38.0302,
  -38.0612,
  -38.0904,
  -38.1184,
  -38.1456,
  -38.1725,
  -38.1983,
  -38.2252,
  -38.2519,
  -38.2783,
  -38.3044,
  -38.3297,
  -38.3538,
  -38.3763,
  -38.3969,
  -38.4155,
  -38.4321,
  -38.4471,
  -38.4611,
  -38.4744,
  -38.4881,
  -38.5023,
  -38.5173,
  -38.533,
  -38.549,
  -38.5639,
  -38.5791,
  -38.5935,
  -38.6075,
  -38.6214,
  -38.6358,
  -38.651,
  -38.6672,
  -38.6846,
  -38.7032,
  -38.7232,
  -38.7447,
  -38.7677,
  -38.7921,
  -38.8175,
  -38.8436,
  -38.8698,
  -38.8959,
  -38.922,
  -38.9479,
  -38.9732,
  -38.9978,
  -39.0203,
  -39.0421,
  -39.0617,
  -39.0794,
  -39.0956,
  -39.1109,
  -39.1265,
  -39.1427,
  -39.1596,
  -39.1771,
  -39.1952,
  -39.2132,
  -39.2312,
  -39.249,
  -39.2665,
  -39.2836,
  -39.3004,
  -39.3168,
  -39.3331,
  -39.3495,
  -39.3662,
  -39.3831,
  -39.4008,
  -39.4175,
  -39.4357,
  -39.4547,
  -39.4748,
  -39.4963,
  -39.5195,
  -39.5444,
  -39.5707,
  -39.5984,
  -39.627,
  -39.6559,
  -39.6853,
  -39.7141,
  -39.7427,
  -39.7707,
  -39.7988,
  -39.8267,
  -39.8546,
  -39.8821,
  -39.9097,
  -39.9371,
  -39.9644,
  -39.9913,
  -40.0172,
  -40.0417,
  -40.0638,
  -40.085,
  -40.1044,
  -40.1223,
  -40.1389,
  -40.1548,
  -40.1703,
  -40.1855,
  -40.1999,
  -40.213,
  -40.2238,
  -40.2318,
  -40.2371,
  -40.2399,
  -40.2409,
  -40.2409,
  -40.2409,
  -40.2412,
  -40.2423,
  -40.2441,
  -40.2461,
  -40.2483,
  -40.2503,
  -40.2524,
  -40.2542,
  -40.2566,
  -40.26,
  -40.265,
  -40.2728,
  -40.2827,
  -40.2971,
  -40.3148,
  -40.3352,
  -40.3575,
  -40.3808,
  -40.4046,
  -40.4284,
  -40.4521,
  -40.4757,
  -40.4998,
  -40.5247,
  -40.55,
  -40.5758,
  -40.6022,
  -40.6288,
  -40.6549,
  -40.6799,
  -40.7035,
  -40.7251,
  -40.7449,
  -40.7631,
  -40.78,
  -40.7961,
  -40.8118,
  -40.8269,
  -40.8417,
  -40.8565,
  -40.8712,
  -40.8855,
  -40.8993,
  -40.9123,
  -40.9247,
  -40.9367,
  -40.9484,
  -40.9589,
  -40.97,
  -40.9803,
  -40.9896,
  -40.9976,
  -41.0045,
  -41.0106,
  -41.0161,
  -41.0215,
  -41.0273,
  -41.034,
  -41.0411,
  -41.0482,
  -41.0543,
  -41.0584,
  -41.0598,
  -41.0582,
  -41.054,
  -41.0476,
  -41.0398,
  -41.0313,
  -41.0222,
  -41.0121,
  -41.0003,
  -40.9859,
  -40.9681,
  -40.9463,
  -40.9195,
  -40.8871,
  -40.8492,
  -40.8045,
  -40.7541,
  -40.6979,
  -40.6374,
  -40.5726,
  -40.5032,
  -40.4288,
  -40.3485,
  -40.2619,
  -40.1688,
  -40.0693,
  -39.9649,
  -33.7887,
  -33.8313,
  -33.8742,
  -33.9161,
  -33.9589,
  -34.0015,
  -34.0437,
  -34.0856,
  -34.1271,
  -34.1682,
  -34.2089,
  -34.2488,
  -34.2881,
  -34.3265,
  -34.3645,
  -34.4022,
  -34.4402,
  -34.4776,
  -34.517,
  -34.5577,
  -34.6,
  -34.6439,
  -34.689,
  -34.7348,
  -34.7806,
  -34.8262,
  -34.8713,
  -34.9152,
  -34.9579,
  -34.9994,
  -35.0396,
  -35.0791,
  -35.117,
  -35.1558,
  -35.1948,
  -35.234,
  -35.2737,
  -35.3139,
  -35.3545,
  -35.3958,
  -35.4373,
  -35.4787,
  -35.52,
  -35.5612,
  -35.6025,
  -35.6443,
  -35.6866,
  -35.7293,
  -35.7713,
  -35.8144,
  -35.8575,
  -35.9002,
  -35.9424,
  -35.9839,
  -36.0249,
  -36.0659,
  -36.107,
  -36.1485,
  -36.1901,
  -36.2317,
  -36.273,
  -36.3143,
  -36.3556,
  -36.3971,
  -36.4378,
  -36.4798,
  -36.5221,
  -36.5647,
  -36.6084,
  -36.6534,
  -36.6999,
  -36.7471,
  -36.7945,
  -36.8415,
  -36.8875,
  -36.9327,
  -36.9772,
  -37.0216,
  -37.0664,
  -37.1114,
  -37.1566,
  -37.2007,
  -37.2455,
  -37.2895,
  -37.3326,
  -37.3743,
  -37.4147,
  -37.4537,
  -37.4919,
  -37.5298,
  -37.568,
  -37.6069,
  -37.6463,
  -37.6859,
  -37.7249,
  -37.763,
  -37.8002,
  -37.8366,
  -37.8722,
  -37.9064,
  -37.9381,
  -37.9693,
  -37.9993,
  -38.0282,
  -38.0565,
  -38.0844,
  -38.112,
  -38.1395,
  -38.1668,
  -38.1938,
  -38.2201,
  -38.2457,
  -38.2697,
  -38.2923,
  -38.3128,
  -38.3315,
  -38.3484,
  -38.3637,
  -38.3782,
  -38.3914,
  -38.4058,
  -38.4206,
  -38.436,
  -38.4518,
  -38.4677,
  -38.4832,
  -38.4982,
  -38.5126,
  -38.5268,
  -38.5414,
  -38.5567,
  -38.5728,
  -38.5898,
  -38.6077,
  -38.6265,
  -38.6464,
  -38.6676,
  -38.6903,
  -38.7146,
  -38.7391,
  -38.7653,
  -38.7916,
  -38.8178,
  -38.8438,
  -38.8697,
  -38.8952,
  -38.92,
  -38.9439,
  -38.9663,
  -38.9868,
  -39.0054,
  -39.0224,
  -39.0383,
  -39.0541,
  -39.0704,
  -39.0872,
  -39.1045,
  -39.1222,
  -39.1403,
  -39.1584,
  -39.1766,
  -39.1945,
  -39.2112,
  -39.2285,
  -39.2453,
  -39.2618,
  -39.2785,
  -39.2956,
  -39.3131,
  -39.3311,
  -39.3498,
  -39.3689,
  -39.3888,
  -39.4099,
  -39.4324,
  -39.4563,
  -39.4816,
  -39.5082,
  -39.5358,
  -39.5645,
  -39.5936,
  -39.6233,
  -39.6528,
  -39.6815,
  -39.7102,
  -39.7385,
  -39.7659,
  -39.7942,
  -39.8224,
  -39.8502,
  -39.878,
  -39.9054,
  -39.9317,
  -39.9569,
  -39.9807,
  -40.0032,
  -40.0243,
  -40.0439,
  -40.0622,
  -40.0794,
  -40.0961,
  -40.1122,
  -40.128,
  -40.1429,
  -40.1557,
  -40.1663,
  -40.1741,
  -40.1791,
  -40.1819,
  -40.183,
  -40.1831,
  -40.1832,
  -40.1836,
  -40.1846,
  -40.1848,
  -40.1861,
  -40.1871,
  -40.1879,
  -40.1887,
  -40.1893,
  -40.1904,
  -40.1927,
  -40.1972,
  -40.2047,
  -40.216,
  -40.2317,
  -40.2511,
  -40.2736,
  -40.2979,
  -40.3232,
  -40.3487,
  -40.3739,
  -40.3986,
  -40.4233,
  -40.4482,
  -40.4734,
  -40.4993,
  -40.526,
  -40.5528,
  -40.5797,
  -40.6064,
  -40.632,
  -40.6561,
  -40.6782,
  -40.6983,
  -40.7168,
  -40.734,
  -40.7493,
  -40.765,
  -40.78,
  -40.7946,
  -40.8091,
  -40.8234,
  -40.8373,
  -40.8508,
  -40.8636,
  -40.8758,
  -40.8876,
  -40.8993,
  -40.9106,
  -40.9215,
  -40.9316,
  -40.9404,
  -40.9482,
  -40.955,
  -40.9613,
  -40.9673,
  -40.9733,
  -40.98,
  -40.9874,
  -40.9955,
  -41.0034,
  -41.0103,
  -41.0151,
  -41.0172,
  -41.0164,
  -41.013,
  -41.0074,
  -41.0003,
  -40.9923,
  -40.9837,
  -40.9741,
  -40.963,
  -40.9493,
  -40.9323,
  -40.9108,
  -40.8845,
  -40.8526,
  -40.8136,
  -40.77,
  -40.7204,
  -40.6653,
  -40.6056,
  -40.5411,
  -40.4721,
  -40.3979,
  -40.3184,
  -40.2331,
  -40.1419,
  -40.0447,
  -39.9423,
  -33.6696,
  -33.7127,
  -33.7557,
  -33.7987,
  -33.8413,
  -33.8837,
  -33.9257,
  -33.9674,
  -34.0089,
  -34.0501,
  -34.0909,
  -34.1311,
  -34.1703,
  -34.2079,
  -34.2458,
  -34.2837,
  -34.322,
  -34.3611,
  -34.4014,
  -34.4431,
  -34.4866,
  -34.5315,
  -34.5775,
  -34.6238,
  -34.6699,
  -34.7154,
  -34.76,
  -34.8024,
  -34.8445,
  -34.8856,
  -34.9259,
  -34.9654,
  -35.0048,
  -35.0445,
  -35.0844,
  -35.1241,
  -35.1645,
  -35.2047,
  -35.2455,
  -35.2865,
  -35.3276,
  -35.3687,
  -35.4094,
  -35.4494,
  -35.4907,
  -35.5326,
  -35.5753,
  -35.6185,
  -35.6621,
  -35.7057,
  -35.7492,
  -35.7923,
  -35.8348,
  -35.8768,
  -35.9184,
  -35.96,
  -36.0018,
  -36.0438,
  -36.086,
  -36.127,
  -36.1689,
  -36.2106,
  -36.2524,
  -36.2943,
  -36.3362,
  -36.3783,
  -36.4206,
  -36.4636,
  -36.5077,
  -36.5534,
  -36.6004,
  -36.6485,
  -36.6967,
  -36.7445,
  -36.7915,
  -36.8375,
  -36.8821,
  -36.9274,
  -36.9727,
  -37.018,
  -37.0634,
  -37.1084,
  -37.1529,
  -37.197,
  -37.2399,
  -37.282,
  -37.3228,
  -37.3625,
  -37.4013,
  -37.4398,
  -37.4783,
  -37.5175,
  -37.5571,
  -37.5968,
  -37.6349,
  -37.6731,
  -37.7102,
  -37.7465,
  -37.7818,
  -37.8159,
  -37.8488,
  -37.8805,
  -37.9113,
  -37.9413,
  -37.9707,
  -37.9997,
  -38.0283,
  -38.0564,
  -38.0839,
  -38.1109,
  -38.1376,
  -38.1631,
  -38.186,
  -38.2083,
  -38.2289,
  -38.2477,
  -38.2649,
  -38.2808,
  -38.2959,
  -38.3109,
  -38.3259,
  -38.3412,
  -38.3568,
  -38.3726,
  -38.3882,
  -38.4033,
  -38.4179,
  -38.4323,
  -38.4468,
  -38.4621,
  -38.4783,
  -38.4953,
  -38.5133,
  -38.5309,
  -38.5501,
  -38.5701,
  -38.5913,
  -38.6138,
  -38.6378,
  -38.6631,
  -38.6891,
  -38.7153,
  -38.7414,
  -38.7672,
  -38.793,
  -38.8186,
  -38.8436,
  -38.8678,
  -38.8908,
  -38.9121,
  -38.9316,
  -38.9493,
  -38.9659,
  -38.982,
  -38.9972,
  -39.0138,
  -39.0308,
  -39.0483,
  -39.0664,
  -39.0847,
  -39.1033,
  -39.1219,
  -39.1402,
  -39.1581,
  -39.1755,
  -39.1924,
  -39.2096,
  -39.2272,
  -39.2453,
  -39.264,
  -39.2833,
  -39.3035,
  -39.3245,
  -39.3467,
  -39.3701,
  -39.3947,
  -39.4204,
  -39.4472,
  -39.4739,
  -39.5023,
  -39.5315,
  -39.5612,
  -39.591,
  -39.6202,
  -39.6493,
  -39.6783,
  -39.7073,
  -39.7363,
  -39.7653,
  -39.7936,
  -39.8215,
  -39.8485,
  -39.8742,
  -39.8986,
  -39.9217,
  -39.9438,
  -39.9647,
  -39.9846,
  -40.0035,
  -40.0216,
  -40.039,
  -40.0559,
  -40.0722,
  -40.087,
  -40.0997,
  -40.1088,
  -40.1162,
  -40.121,
  -40.1237,
  -40.125,
  -40.1254,
  -40.1255,
  -40.1258,
  -40.1261,
  -40.1266,
  -40.1269,
  -40.1267,
  -40.1262,
  -40.1256,
  -40.1249,
  -40.1249,
  -40.1263,
  -40.1303,
  -40.1376,
  -40.1496,
  -40.1664,
  -40.1875,
  -40.2124,
  -40.2391,
  -40.2667,
  -40.2944,
  -40.3214,
  -40.3479,
  -40.3738,
  -40.3996,
  -40.4245,
  -40.4509,
  -40.4778,
  -40.505,
  -40.5322,
  -40.559,
  -40.5848,
  -40.609,
  -40.6313,
  -40.6516,
  -40.6703,
  -40.6877,
  -40.7042,
  -40.72,
  -40.7351,
  -40.7498,
  -40.764,
  -40.7779,
  -40.7913,
  -40.8042,
  -40.8166,
  -40.8286,
  -40.8403,
  -40.852,
  -40.8634,
  -40.8743,
  -40.8843,
  -40.893,
  -40.9009,
  -40.9079,
  -40.9144,
  -40.9207,
  -40.9273,
  -40.9346,
  -40.9424,
  -40.9509,
  -40.9591,
  -40.9663,
  -40.9705,
  -40.9731,
  -40.973,
  -40.9703,
  -40.9655,
  -40.959,
  -40.9515,
  -40.9432,
  -40.934,
  -40.9231,
  -40.9098,
  -40.8932,
  -40.8723,
  -40.8468,
  -40.8155,
  -40.7785,
  -40.7357,
  -40.6872,
  -40.6332,
  -40.5742,
  -40.5101,
  -40.4412,
  -40.3678,
  -40.289,
  -40.205,
  -40.1149,
  -40.0195,
  -39.9188,
  -33.5531,
  -33.5968,
  -33.6401,
  -33.683,
  -33.7255,
  -33.7675,
  -33.8093,
  -33.851,
  -33.8914,
  -33.9329,
  -33.9737,
  -34.014,
  -34.0533,
  -34.0919,
  -34.1301,
  -34.1683,
  -34.207,
  -34.2469,
  -34.2881,
  -34.3309,
  -34.3753,
  -34.421,
  -34.4675,
  -34.5133,
  -34.5594,
  -34.6047,
  -34.6488,
  -34.6917,
  -34.7335,
  -34.7745,
  -34.8149,
  -34.8549,
  -34.895,
  -34.9353,
  -34.9757,
  -35.0163,
  -35.057,
  -35.0977,
  -35.1374,
  -35.1783,
  -35.2191,
  -35.2599,
  -35.3005,
  -35.3414,
  -35.3827,
  -35.4248,
  -35.4677,
  -35.5112,
  -35.5551,
  -35.5992,
  -35.6431,
  -35.6865,
  -35.7294,
  -35.7718,
  -35.813,
  -35.855,
  -35.8973,
  -35.9397,
  -35.9823,
  -36.0247,
  -36.0671,
  -36.1094,
  -36.1516,
  -36.1941,
  -36.2364,
  -36.2789,
  -36.3215,
  -36.3648,
  -36.4093,
  -36.4553,
  -36.5016,
  -36.55,
  -36.5987,
  -36.6472,
  -36.6952,
  -36.7426,
  -36.7894,
  -36.8358,
  -36.8817,
  -36.9273,
  -36.9727,
  -37.0177,
  -37.0622,
  -37.1058,
  -37.149,
  -37.1912,
  -37.2325,
  -37.2729,
  -37.3115,
  -37.3506,
  -37.3895,
  -37.4287,
  -37.4683,
  -37.508,
  -37.5472,
  -37.5858,
  -37.6231,
  -37.6595,
  -37.6948,
  -37.729,
  -37.7622,
  -37.7945,
  -37.8261,
  -37.857,
  -37.8874,
  -37.9172,
  -37.9449,
  -37.9735,
  -38.0012,
  -38.0287,
  -38.0551,
  -38.0806,
  -38.1043,
  -38.1265,
  -38.147,
  -38.166,
  -38.1835,
  -38.1998,
  -38.2156,
  -38.231,
  -38.2465,
  -38.2622,
  -38.278,
  -38.2938,
  -38.3091,
  -38.3239,
  -38.3373,
  -38.3518,
  -38.3667,
  -38.3826,
  -38.3996,
  -38.4177,
  -38.4367,
  -38.4563,
  -38.4763,
  -38.4967,
  -38.518,
  -38.5403,
  -38.564,
  -38.5888,
  -38.6145,
  -38.6403,
  -38.6661,
  -38.6917,
  -38.7176,
  -38.743,
  -38.7681,
  -38.7915,
  -38.8151,
  -38.8371,
  -38.8572,
  -38.8757,
  -38.8928,
  -38.9091,
  -38.9252,
  -38.9416,
  -38.9584,
  -38.9758,
  -38.994,
  -39.0127,
  -39.0318,
  -39.051,
  -39.0699,
  -39.0884,
  -39.1063,
  -39.1238,
  -39.1415,
  -39.1596,
  -39.1783,
  -39.1978,
  -39.2168,
  -39.2381,
  -39.2604,
  -39.2838,
  -39.3083,
  -39.3339,
  -39.3601,
  -39.3871,
  -39.4145,
  -39.4428,
  -39.4719,
  -39.5015,
  -39.5312,
  -39.5609,
  -39.5904,
  -39.6201,
  -39.6499,
  -39.6796,
  -39.7091,
  -39.7378,
  -39.7657,
  -39.7923,
  -39.8174,
  -39.8411,
  -39.8636,
  -39.8852,
  -39.9051,
  -39.9254,
  -39.9449,
  -39.9637,
  -39.982,
  -39.9996,
  -40.0161,
  -40.0307,
  -40.0431,
  -40.0526,
  -40.0595,
  -40.0641,
  -40.0669,
  -40.0684,
  -40.0689,
  -40.0691,
  -40.0689,
  -40.0687,
  -40.0682,
  -40.0671,
  -40.0657,
  -40.064,
  -40.0622,
  -40.0602,
  -40.0591,
  -40.0597,
  -40.0633,
  -40.0709,
  -40.0835,
  -40.1006,
  -40.1238,
  -40.1509,
  -40.1802,
  -40.2106,
  -40.2407,
  -40.27,
  -40.2981,
  -40.3256,
  -40.3527,
  -40.3794,
  -40.4063,
  -40.4334,
  -40.4608,
  -40.488,
  -40.5147,
  -40.5405,
  -40.5645,
  -40.5865,
  -40.6066,
  -40.6252,
  -40.6426,
  -40.6594,
  -40.6756,
  -40.6911,
  -40.706,
  -40.7201,
  -40.7336,
  -40.7465,
  -40.7587,
  -40.7705,
  -40.7819,
  -40.7936,
  -40.8053,
  -40.8171,
  -40.8274,
  -40.8377,
  -40.8467,
  -40.855,
  -40.8622,
  -40.8691,
  -40.8759,
  -40.8829,
  -40.8904,
  -40.8984,
  -40.9066,
  -40.9147,
  -40.9216,
  -40.9268,
  -40.9298,
  -40.9302,
  -40.9282,
  -40.924,
  -40.918,
  -40.9108,
  -40.9027,
  -40.8936,
  -40.8827,
  -40.8697,
  -40.8535,
  -40.8334,
  -40.8085,
  -40.7784,
  -40.7424,
  -40.7008,
  -40.6533,
  -40.6003,
  -40.5421,
  -40.4787,
  -40.4103,
  -40.3373,
  -40.2594,
  -40.1765,
  -40.088,
  -39.9938,
  -39.8944,
  -33.438,
  -33.4824,
  -33.526,
  -33.568,
  -33.6103,
  -33.6521,
  -33.6936,
  -33.7351,
  -33.7763,
  -33.8177,
  -33.8587,
  -33.8987,
  -33.9383,
  -33.9773,
  -34.0158,
  -34.0544,
  -34.0939,
  -34.1347,
  -34.1759,
  -34.2198,
  -34.2651,
  -34.3117,
  -34.3587,
  -34.4054,
  -34.4514,
  -34.4962,
  -34.5398,
  -34.5823,
  -34.624,
  -34.665,
  -34.7056,
  -34.746,
  -34.7865,
  -34.8264,
  -34.8675,
  -34.9087,
  -34.9497,
  -34.9908,
  -35.0318,
  -35.0728,
  -35.1138,
  -35.1547,
  -35.1955,
  -35.2365,
  -35.278,
  -35.3202,
  -35.3632,
  -35.407,
  -35.4501,
  -35.4944,
  -35.5385,
  -35.5823,
  -35.6256,
  -35.6683,
  -35.7106,
  -35.7529,
  -35.7954,
  -35.8381,
  -35.8808,
  -35.9236,
  -35.9664,
  -36.0092,
  -36.0521,
  -36.0951,
  -36.1382,
  -36.18,
  -36.2233,
  -36.2672,
  -36.3119,
  -36.3579,
  -36.4054,
  -36.4538,
  -36.5029,
  -36.5522,
  -36.6013,
  -36.6502,
  -36.6984,
  -36.7458,
  -36.7925,
  -36.8385,
  -36.884,
  -36.9289,
  -36.9723,
  -37.0161,
  -37.0591,
  -37.1016,
  -37.1433,
  -37.1842,
  -37.2245,
  -37.2642,
  -37.3036,
  -37.3431,
  -37.3828,
  -37.4225,
  -37.4619,
  -37.5007,
  -37.5383,
  -37.5749,
  -37.6105,
  -37.645,
  -37.6777,
  -37.7105,
  -37.7428,
  -37.7746,
  -37.8056,
  -37.8356,
  -37.8649,
  -37.8933,
  -37.9214,
  -37.9484,
  -37.975,
  -38.0001,
  -38.0237,
  -38.0457,
  -38.0662,
  -38.0853,
  -38.103,
  -38.1198,
  -38.136,
  -38.151,
  -38.1669,
  -38.183,
  -38.1988,
  -38.2144,
  -38.2296,
  -38.2442,
  -38.2585,
  -38.2732,
  -38.2886,
  -38.3051,
  -38.323,
  -38.3422,
  -38.3623,
  -38.3831,
  -38.4041,
  -38.4253,
  -38.4467,
  -38.4689,
  -38.4922,
  -38.5165,
  -38.5405,
  -38.5659,
  -38.5913,
  -38.6166,
  -38.6417,
  -38.6668,
  -38.6918,
  -38.7166,
  -38.7407,
  -38.7633,
  -38.7842,
  -38.8034,
  -38.821,
  -38.8376,
  -38.8538,
  -38.8699,
  -38.8869,
  -38.9044,
  -38.9227,
  -38.9417,
  -38.9611,
  -38.9807,
  -38.9992,
  -39.0183,
  -39.0369,
  -39.0551,
  -39.0733,
  -39.092,
  -39.1112,
  -39.1313,
  -39.1524,
  -39.1746,
  -39.1981,
  -39.2228,
  -39.2484,
  -39.2749,
  -39.3018,
  -39.3289,
  -39.3564,
  -39.3846,
  -39.4135,
  -39.443,
  -39.4727,
  -39.5025,
  -39.5326,
  -39.5629,
  -39.5935,
  -39.623,
  -39.6529,
  -39.6817,
  -39.7094,
  -39.7355,
  -39.76,
  -39.783,
  -39.8052,
  -39.8265,
  -39.8473,
  -39.8678,
  -39.8878,
  -39.9072,
  -39.9261,
  -39.944,
  -39.9606,
  -39.975,
  -39.9868,
  -39.9958,
  -40.0023,
  -40.0067,
  -40.0095,
  -40.0113,
  -40.012,
  -40.0122,
  -40.0119,
  -40.0111,
  -40.0096,
  -40.0064,
  -40.0037,
  -40.0008,
  -39.9976,
  -39.9945,
  -39.9923,
  -39.9924,
  -39.9959,
  -40.0039,
  -40.0174,
  -40.0371,
  -40.0624,
  -40.0919,
  -40.1242,
  -40.1573,
  -40.1899,
  -40.2217,
  -40.2519,
  -40.281,
  -40.309,
  -40.3366,
  -40.3639,
  -40.3912,
  -40.4185,
  -40.4456,
  -40.4721,
  -40.4973,
  -40.5209,
  -40.5424,
  -40.5622,
  -40.5808,
  -40.5984,
  -40.6143,
  -40.6311,
  -40.647,
  -40.6622,
  -40.6764,
  -40.6898,
  -40.7022,
  -40.7137,
  -40.7248,
  -40.7358,
  -40.7471,
  -40.7588,
  -40.7707,
  -40.7824,
  -40.7931,
  -40.8029,
  -40.8117,
  -40.8196,
  -40.8271,
  -40.8343,
  -40.8416,
  -40.8491,
  -40.8568,
  -40.8646,
  -40.872,
  -40.8785,
  -40.8834,
  -40.8865,
  -40.8872,
  -40.8857,
  -40.8822,
  -40.8766,
  -40.8696,
  -40.8615,
  -40.8523,
  -40.8415,
  -40.8284,
  -40.8125,
  -40.7929,
  -40.769,
  -40.7398,
  -40.705,
  -40.6636,
  -40.617,
  -40.5653,
  -40.5079,
  -40.445,
  -40.3775,
  -40.3053,
  -40.2283,
  -40.1465,
  -40.0595,
  -39.9667,
  -39.8684,
  -33.3229,
  -33.3682,
  -33.4123,
  -33.4556,
  -33.4978,
  -33.5395,
  -33.5809,
  -33.6219,
  -33.663,
  -33.704,
  -33.7447,
  -33.785,
  -33.8249,
  -33.863,
  -33.902,
  -33.9413,
  -33.9816,
  -34.0233,
  -34.0666,
  -34.1116,
  -34.1579,
  -34.2049,
  -34.252,
  -34.2985,
  -34.344,
  -34.3885,
  -34.4318,
  -34.4741,
  -34.5148,
  -34.556,
  -34.5969,
  -34.6377,
  -34.6786,
  -34.7197,
  -34.7614,
  -34.8029,
  -34.844,
  -34.8856,
  -34.9272,
  -34.9687,
  -35.0103,
  -35.0518,
  -35.0931,
  -35.1336,
  -35.1753,
  -35.2177,
  -35.2607,
  -35.3044,
  -35.3486,
  -35.393,
  -35.4374,
  -35.4813,
  -35.5247,
  -35.5675,
  -35.61,
  -35.6524,
  -35.695,
  -35.7376,
  -35.7805,
  -35.8224,
  -35.8655,
  -35.9089,
  -35.9525,
  -35.9961,
  -36.0398,
  -36.0835,
  -36.1274,
  -36.1718,
  -36.2173,
  -36.2633,
  -36.3107,
  -36.3592,
  -36.4086,
  -36.4587,
  -36.5091,
  -36.5593,
  -36.6077,
  -36.6562,
  -36.7037,
  -36.7502,
  -36.7959,
  -36.841,
  -36.8854,
  -36.9293,
  -36.9725,
  -37.0151,
  -37.0571,
  -37.0984,
  -37.1392,
  -37.1794,
  -37.2193,
  -37.2589,
  -37.2989,
  -37.339,
  -37.3778,
  -37.417,
  -37.4551,
  -37.4921,
  -37.528,
  -37.563,
  -37.5971,
  -37.6306,
  -37.6634,
  -37.6957,
  -37.727,
  -37.7573,
  -37.7863,
  -37.8146,
  -37.8422,
  -37.8691,
  -37.8953,
  -37.9202,
  -37.9436,
  -37.9645,
  -37.985,
  -38.0042,
  -38.0222,
  -38.0392,
  -38.0557,
  -38.0722,
  -38.0885,
  -38.1048,
  -38.1209,
  -38.1365,
  -38.1515,
  -38.1661,
  -38.1807,
  -38.1958,
  -38.2117,
  -38.2287,
  -38.2474,
  -38.2677,
  -38.289,
  -38.31,
  -38.3322,
  -38.3541,
  -38.376,
  -38.3982,
  -38.4211,
  -38.4448,
  -38.4692,
  -38.494,
  -38.5189,
  -38.5436,
  -38.5684,
  -38.5929,
  -38.6179,
  -38.6432,
  -38.6673,
  -38.6904,
  -38.7119,
  -38.7317,
  -38.7498,
  -38.7668,
  -38.7834,
  -38.7988,
  -38.8159,
  -38.8335,
  -38.8521,
  -38.8713,
  -38.891,
  -38.9109,
  -38.9308,
  -38.9505,
  -38.9697,
  -38.9886,
  -39.0074,
  -39.0264,
  -39.0461,
  -39.0667,
  -39.0885,
  -39.1118,
  -39.1364,
  -39.1622,
  -39.189,
  -39.2163,
  -39.2438,
  -39.2714,
  -39.299,
  -39.3263,
  -39.3552,
  -39.3846,
  -39.4142,
  -39.444,
  -39.4743,
  -39.5052,
  -39.5364,
  -39.5673,
  -39.5974,
  -39.6261,
  -39.6533,
  -39.6788,
  -39.7028,
  -39.7256,
  -39.7475,
  -39.7687,
  -39.7897,
  -39.8103,
  -39.8306,
  -39.8505,
  -39.8697,
  -39.8877,
  -39.9041,
  -39.9181,
  -39.9294,
  -39.9369,
  -39.9431,
  -39.9473,
  -39.9502,
  -39.9521,
  -39.9531,
  -39.9534,
  -39.9531,
  -39.9519,
  -39.9495,
  -39.9463,
  -39.9426,
  -39.9384,
  -39.9341,
  -39.9301,
  -39.9274,
  -39.9272,
  -39.9308,
  -39.9393,
  -39.9543,
  -39.9757,
  -40.0031,
  -40.0351,
  -40.0699,
  -40.1057,
  -40.1409,
  -40.1748,
  -40.207,
  -40.2376,
  -40.2671,
  -40.2954,
  -40.3221,
  -40.3495,
  -40.3767,
  -40.4035,
  -40.4295,
  -40.4541,
  -40.4769,
  -40.4979,
  -40.5174,
  -40.5358,
  -40.5534,
  -40.5709,
  -40.5879,
  -40.6042,
  -40.6198,
  -40.6345,
  -40.6479,
  -40.6601,
  -40.6712,
  -40.6816,
  -40.692,
  -40.7028,
  -40.7142,
  -40.7261,
  -40.738,
  -40.7493,
  -40.7597,
  -40.7693,
  -40.7781,
  -40.7864,
  -40.7942,
  -40.8018,
  -40.8092,
  -40.8165,
  -40.8234,
  -40.83,
  -40.8356,
  -40.8401,
  -40.842,
  -40.8431,
  -40.842,
  -40.8389,
  -40.8338,
  -40.8271,
  -40.819,
  -40.8095,
  -40.7982,
  -40.7849,
  -40.7689,
  -40.7498,
  -40.7266,
  -40.6985,
  -40.665,
  -40.6256,
  -40.5805,
  -40.5296,
  -40.4731,
  -40.4113,
  -40.3445,
  -40.2734,
  -40.1977,
  -40.1175,
  -40.0319,
  -39.9407,
  -39.8437,
  -33.2102,
  -33.2561,
  -33.301,
  -33.3446,
  -33.387,
  -33.4286,
  -33.4697,
  -33.5105,
  -33.5504,
  -33.5912,
  -33.6318,
  -33.6721,
  -33.712,
  -33.7515,
  -33.7909,
  -33.8309,
  -33.8721,
  -33.9148,
  -33.9593,
  -34.0052,
  -34.0521,
  -34.0994,
  -34.1464,
  -34.1916,
  -34.2368,
  -34.281,
  -34.3241,
  -34.3665,
  -34.4083,
  -34.4498,
  -34.4911,
  -34.5322,
  -34.5733,
  -34.6146,
  -34.6562,
  -34.6978,
  -34.7393,
  -34.7815,
  -34.8227,
  -34.8651,
  -34.9075,
  -34.9498,
  -34.992,
  -35.0341,
  -35.0763,
  -35.1188,
  -35.1617,
  -35.2053,
  -35.2494,
  -35.2939,
  -35.3382,
  -35.382,
  -35.4253,
  -35.4682,
  -35.5097,
  -35.5522,
  -35.5948,
  -35.6375,
  -35.6803,
  -35.7234,
  -35.7669,
  -35.8107,
  -35.8547,
  -35.899,
  -35.9433,
  -35.9877,
  -36.0323,
  -36.0774,
  -36.1232,
  -36.1699,
  -36.2175,
  -36.2652,
  -36.315,
  -36.3658,
  -36.4172,
  -36.4685,
  -36.5191,
  -36.5685,
  -36.6167,
  -36.6638,
  -36.71,
  -36.7554,
  -36.8002,
  -36.8445,
  -36.8879,
  -36.9308,
  -36.973,
  -37.0147,
  -37.0548,
  -37.0954,
  -37.1355,
  -37.1755,
  -37.2157,
  -37.2562,
  -37.2965,
  -37.3362,
  -37.3748,
  -37.4123,
  -37.4487,
  -37.4841,
  -37.5189,
  -37.553,
  -37.5864,
  -37.619,
  -37.6505,
  -37.6805,
  -37.7091,
  -37.7357,
  -37.7627,
  -37.7892,
  -37.815,
  -37.8398,
  -37.863,
  -37.8848,
  -37.9054,
  -37.9246,
  -37.9427,
  -37.9599,
  -37.9767,
  -37.9934,
  -38.0101,
  -38.0268,
  -38.0431,
  -38.0588,
  -38.0739,
  -38.0887,
  -38.1025,
  -38.1179,
  -38.1343,
  -38.1522,
  -38.1718,
  -38.1929,
  -38.2154,
  -38.2386,
  -38.2619,
  -38.2848,
  -38.3073,
  -38.3296,
  -38.3523,
  -38.3755,
  -38.3993,
  -38.4234,
  -38.4475,
  -38.4715,
  -38.4957,
  -38.5201,
  -38.5451,
  -38.5691,
  -38.5938,
  -38.6175,
  -38.6396,
  -38.6599,
  -38.6787,
  -38.6963,
  -38.7133,
  -38.7303,
  -38.7476,
  -38.7655,
  -38.7843,
  -38.8036,
  -38.8236,
  -38.8439,
  -38.8641,
  -38.8843,
  -38.9041,
  -38.9237,
  -38.943,
  -38.9624,
  -38.9823,
  -39.0032,
  -39.0256,
  -39.0486,
  -39.0741,
  -39.1009,
  -39.1285,
  -39.1565,
  -39.1847,
  -39.2128,
  -39.241,
  -39.2698,
  -39.2989,
  -39.3281,
  -39.3575,
  -39.3873,
  -39.4177,
  -39.4487,
  -39.4801,
  -39.5112,
  -39.541,
  -39.5693,
  -39.5959,
  -39.6209,
  -39.6446,
  -39.6672,
  -39.689,
  -39.7104,
  -39.7304,
  -39.7514,
  -39.7719,
  -39.792,
  -39.8114,
  -39.8292,
  -39.8452,
  -39.8587,
  -39.8695,
  -39.8777,
  -39.8836,
  -39.888,
  -39.8909,
  -39.8929,
  -39.8943,
  -39.8948,
  -39.8944,
  -39.8929,
  -39.8902,
  -39.8862,
  -39.8815,
  -39.8762,
  -39.871,
  -39.8664,
  -39.8634,
  -39.8632,
  -39.8674,
  -39.8772,
  -39.8936,
  -39.9159,
  -39.9455,
  -39.9799,
  -40.017,
  -40.055,
  -40.0924,
  -40.1283,
  -40.1623,
  -40.1944,
  -40.2248,
  -40.2538,
  -40.2819,
  -40.3094,
  -40.3366,
  -40.3631,
  -40.3886,
  -40.4126,
  -40.4349,
  -40.4554,
  -40.4746,
  -40.4929,
  -40.5107,
  -40.5283,
  -40.5456,
  -40.5625,
  -40.5786,
  -40.5936,
  -40.6072,
  -40.6193,
  -40.6301,
  -40.6399,
  -40.6497,
  -40.6599,
  -40.6708,
  -40.6823,
  -40.6931,
  -40.7047,
  -40.7156,
  -40.726,
  -40.7359,
  -40.7451,
  -40.7536,
  -40.7616,
  -40.7689,
  -40.7756,
  -40.7818,
  -40.7872,
  -40.792,
  -40.7959,
  -40.7986,
  -40.7998,
  -40.7992,
  -40.7965,
  -40.7917,
  -40.785,
  -40.7767,
  -40.7668,
  -40.7548,
  -40.7409,
  -40.7247,
  -40.7057,
  -40.6831,
  -40.6561,
  -40.6238,
  -40.5859,
  -40.5421,
  -40.4923,
  -40.4369,
  -40.3761,
  -40.3103,
  -40.2403,
  -40.1661,
  -40.0876,
  -40.0042,
  -39.915,
  -39.8201,
  -33.0986,
  -33.1454,
  -33.191,
  -33.2351,
  -33.2769,
  -33.3185,
  -33.3594,
  -33.4,
  -33.4406,
  -33.4813,
  -33.5219,
  -33.5622,
  -33.6021,
  -33.6419,
  -33.6818,
  -33.7225,
  -33.7646,
  -33.8083,
  -33.8527,
  -33.8994,
  -33.9467,
  -33.9939,
  -34.0407,
  -34.0867,
  -34.1315,
  -34.1757,
  -34.219,
  -34.2617,
  -34.3039,
  -34.3458,
  -34.3873,
  -34.4286,
  -34.4698,
  -34.5098,
  -34.5509,
  -34.5925,
  -34.6346,
  -34.6774,
  -34.7205,
  -34.764,
  -34.8075,
  -34.851,
  -34.8941,
  -34.9369,
  -34.9796,
  -35.0223,
  -35.065,
  -35.1083,
  -35.1521,
  -35.1952,
  -35.2392,
  -35.2828,
  -35.3259,
  -35.3686,
  -35.4112,
  -35.4539,
  -35.4967,
  -35.5395,
  -35.5825,
  -35.6257,
  -35.6694,
  -35.7135,
  -35.7579,
  -35.8027,
  -35.8476,
  -35.8916,
  -35.937,
  -35.9828,
  -36.0293,
  -36.0767,
  -36.1249,
  -36.1741,
  -36.2243,
  -36.2757,
  -36.3278,
  -36.38,
  -36.4314,
  -36.4815,
  -36.5304,
  -36.5782,
  -36.6249,
  -36.671,
  -36.7155,
  -36.7603,
  -36.8043,
  -36.8475,
  -36.89,
  -36.932,
  -36.9734,
  -37.0143,
  -37.0546,
  -37.0947,
  -37.1353,
  -37.1761,
  -37.2168,
  -37.257,
  -37.2961,
  -37.334,
  -37.3709,
  -37.4068,
  -37.4413,
  -37.4761,
  -37.5102,
  -37.543,
  -37.5743,
  -37.6038,
  -37.6317,
  -37.6587,
  -37.6851,
  -37.711,
  -37.7363,
  -37.7608,
  -37.7839,
  -37.8057,
  -37.8265,
  -37.8457,
  -37.8638,
  -37.8811,
  -37.8979,
  -37.9148,
  -37.9309,
  -37.948,
  -37.9646,
  -37.9806,
  -37.996,
  -38.011,
  -38.0262,
  -38.0421,
  -38.0591,
  -38.0776,
  -38.0977,
  -38.1196,
  -38.1431,
  -38.1674,
  -38.1918,
  -38.2157,
  -38.2389,
  -38.2617,
  -38.2843,
  -38.3071,
  -38.3294,
  -38.3527,
  -38.3761,
  -38.3994,
  -38.4231,
  -38.4473,
  -38.4721,
  -38.4973,
  -38.5223,
  -38.5464,
  -38.5691,
  -38.5901,
  -38.6097,
  -38.6281,
  -38.6459,
  -38.6634,
  -38.6811,
  -38.6993,
  -38.7182,
  -38.7378,
  -38.758,
  -38.7784,
  -38.7992,
  -38.8189,
  -38.8395,
  -38.8597,
  -38.8795,
  -38.8992,
  -38.9192,
  -38.9402,
  -38.9627,
  -38.9871,
  -39.0133,
  -39.0407,
  -39.069,
  -39.0976,
  -39.1263,
  -39.1552,
  -39.1843,
  -39.2136,
  -39.243,
  -39.2722,
  -39.3015,
  -39.3311,
  -39.3614,
  -39.3923,
  -39.4237,
  -39.4544,
  -39.4826,
  -39.5102,
  -39.5361,
  -39.5605,
  -39.584,
  -39.6066,
  -39.6286,
  -39.6501,
  -39.6714,
  -39.6927,
  -39.7134,
  -39.7338,
  -39.7529,
  -39.7705,
  -39.7859,
  -39.7989,
  -39.8094,
  -39.8175,
  -39.8236,
  -39.828,
  -39.8312,
  -39.8335,
  -39.835,
  -39.8358,
  -39.8355,
  -39.834,
  -39.8309,
  -39.8252,
  -39.8196,
  -39.8136,
  -39.8078,
  -39.8027,
  -39.7997,
  -39.8001,
  -39.8053,
  -39.8168,
  -39.8351,
  -39.8607,
  -39.8923,
  -39.9287,
  -39.9678,
  -40.0075,
  -40.0467,
  -40.0842,
  -40.1194,
  -40.1526,
  -40.1838,
  -40.2134,
  -40.2418,
  -40.2695,
  -40.2968,
  -40.3234,
  -40.3486,
  -40.3722,
  -40.394,
  -40.4141,
  -40.433,
  -40.4512,
  -40.4691,
  -40.4869,
  -40.5035,
  -40.5207,
  -40.5372,
  -40.5525,
  -40.5663,
  -40.5783,
  -40.5889,
  -40.5984,
  -40.6076,
  -40.6172,
  -40.6273,
  -40.6381,
  -40.6494,
  -40.661,
  -40.6723,
  -40.6835,
  -40.6942,
  -40.7044,
  -40.7138,
  -40.722,
  -40.7292,
  -40.7355,
  -40.7409,
  -40.7455,
  -40.7496,
  -40.7529,
  -40.7553,
  -40.7565,
  -40.7561,
  -40.7534,
  -40.7487,
  -40.7419,
  -40.7332,
  -40.7225,
  -40.7099,
  -40.6953,
  -40.6786,
  -40.6595,
  -40.6373,
  -40.6113,
  -40.5804,
  -40.544,
  -40.5006,
  -40.4521,
  -40.3975,
  -40.3378,
  -40.2733,
  -40.2046,
  -40.1324,
  -40.056,
  -39.9752,
  -39.8889,
  -39.797,
  -32.9881,
  -33.0353,
  -33.0814,
  -33.126,
  -33.1691,
  -33.2108,
  -33.2516,
  -33.2921,
  -33.3325,
  -33.3731,
  -33.4137,
  -33.4542,
  -33.4944,
  -33.5336,
  -33.5741,
  -33.6156,
  -33.6584,
  -33.7029,
  -33.7489,
  -33.7959,
  -33.843,
  -33.8899,
  -33.9364,
  -33.9821,
  -34.0272,
  -34.0714,
  -34.1152,
  -34.1588,
  -34.2004,
  -34.2429,
  -34.285,
  -34.3267,
  -34.3679,
  -34.4089,
  -34.4498,
  -34.4914,
  -34.5335,
  -34.5766,
  -34.6206,
  -34.6649,
  -34.7094,
  -34.7536,
  -34.7976,
  -34.8412,
  -34.8834,
  -34.9261,
  -34.9688,
  -35.0118,
  -35.0552,
  -35.0988,
  -35.1424,
  -35.1856,
  -35.2284,
  -35.2709,
  -35.3135,
  -35.3563,
  -35.3993,
  -35.4424,
  -35.4856,
  -35.5292,
  -35.572,
  -35.6164,
  -35.6611,
  -35.7063,
  -35.7518,
  -35.7976,
  -35.8437,
  -35.8903,
  -35.9377,
  -35.9858,
  -36.0346,
  -36.0844,
  -36.1352,
  -36.1869,
  -36.2396,
  -36.2924,
  -36.3445,
  -36.3943,
  -36.4439,
  -36.4924,
  -36.5399,
  -36.5867,
  -36.6329,
  -36.6781,
  -36.7226,
  -36.7664,
  -36.8094,
  -36.8518,
  -36.8939,
  -36.9349,
  -36.9755,
  -37.0158,
  -37.0563,
  -37.0974,
  -37.1372,
  -37.1777,
  -37.2171,
  -37.2555,
  -37.2929,
  -37.3296,
  -37.3657,
  -37.4012,
  -37.4358,
  -37.4688,
  -37.4999,
  -37.5289,
  -37.5561,
  -37.5822,
  -37.6081,
  -37.6333,
  -37.6581,
  -37.6822,
  -37.7053,
  -37.7262,
  -37.7469,
  -37.7665,
  -37.7847,
  -37.8021,
  -37.819,
  -37.836,
  -37.8532,
  -37.8705,
  -37.8874,
  -37.9035,
  -37.919,
  -37.9343,
  -37.95,
  -37.9666,
  -37.9842,
  -38.0032,
  -38.024,
  -38.0467,
  -38.071,
  -38.0953,
  -38.1206,
  -38.1454,
  -38.1694,
  -38.1927,
  -38.2155,
  -38.2383,
  -38.2609,
  -38.2837,
  -38.3065,
  -38.3292,
  -38.3523,
  -38.376,
  -38.4007,
  -38.4259,
  -38.4512,
  -38.4758,
  -38.4992,
  -38.5213,
  -38.5419,
  -38.5614,
  -38.5801,
  -38.5974,
  -38.6155,
  -38.634,
  -38.6531,
  -38.6728,
  -38.6932,
  -38.7141,
  -38.7352,
  -38.7568,
  -38.778,
  -38.799,
  -38.8192,
  -38.839,
  -38.859,
  -38.8799,
  -38.9023,
  -38.9269,
  -38.9533,
  -38.9809,
  -39.0097,
  -39.0391,
  -39.0687,
  -39.0985,
  -39.1283,
  -39.1571,
  -39.1867,
  -39.2159,
  -39.2449,
  -39.2741,
  -39.3039,
  -39.3345,
  -39.3655,
  -39.3954,
  -39.4237,
  -39.4505,
  -39.4757,
  -39.4999,
  -39.5232,
  -39.5457,
  -39.5678,
  -39.5897,
  -39.6115,
  -39.6331,
  -39.6541,
  -39.6745,
  -39.6934,
  -39.7106,
  -39.7255,
  -39.7382,
  -39.7486,
  -39.7568,
  -39.7621,
  -39.767,
  -39.7706,
  -39.7732,
  -39.7751,
  -39.7761,
  -39.7759,
  -39.7743,
  -39.7711,
  -39.766,
  -39.7597,
  -39.753,
  -39.7466,
  -39.7417,
  -39.7391,
  -39.7405,
  -39.7473,
  -39.7607,
  -39.7811,
  -39.8086,
  -39.8423,
  -39.8802,
  -39.9208,
  -39.962,
  -40.0025,
  -40.0412,
  -40.0773,
  -40.1113,
  -40.1429,
  -40.1731,
  -40.2019,
  -40.229,
  -40.2563,
  -40.2828,
  -40.3079,
  -40.3315,
  -40.3531,
  -40.3732,
  -40.3921,
  -40.4104,
  -40.4283,
  -40.4462,
  -40.4639,
  -40.4814,
  -40.498,
  -40.5133,
  -40.527,
  -40.5389,
  -40.5492,
  -40.5584,
  -40.5673,
  -40.5762,
  -40.5858,
  -40.5959,
  -40.6067,
  -40.6179,
  -40.6295,
  -40.6411,
  -40.6526,
  -40.6635,
  -40.6734,
  -40.682,
  -40.6891,
  -40.6949,
  -40.6997,
  -40.7037,
  -40.707,
  -40.7096,
  -40.7119,
  -40.7117,
  -40.7109,
  -40.7081,
  -40.7033,
  -40.6963,
  -40.6871,
  -40.6758,
  -40.6624,
  -40.647,
  -40.6298,
  -40.6106,
  -40.5887,
  -40.5634,
  -40.5336,
  -40.4984,
  -40.4573,
  -40.4101,
  -40.357,
  -40.2987,
  -40.2362,
  -40.1696,
  -40.0993,
  -40.0259,
  -39.9477,
  -39.8647,
  -39.7759,
  -32.8808,
  -32.9282,
  -32.9746,
  -33.0194,
  -33.0628,
  -33.1046,
  -33.1455,
  -33.1859,
  -33.2264,
  -33.2659,
  -33.3066,
  -33.3473,
  -33.3879,
  -33.4286,
  -33.4697,
  -33.5119,
  -33.5555,
  -33.6005,
  -33.6467,
  -33.6936,
  -33.7404,
  -33.7867,
  -33.8327,
  -33.8774,
  -33.9226,
  -33.9675,
  -34.0122,
  -34.0564,
  -34.1002,
  -34.1436,
  -34.1863,
  -34.2283,
  -34.2696,
  -34.3104,
  -34.3513,
  -34.3927,
  -34.4351,
  -34.4786,
  -34.5222,
  -34.5673,
  -34.6125,
  -34.6574,
  -34.7021,
  -34.7461,
  -34.7895,
  -34.8323,
  -34.8748,
  -34.9174,
  -34.9602,
  -35.0032,
  -35.0462,
  -35.0889,
  -35.1314,
  -35.1738,
  -35.2153,
  -35.2582,
  -35.3014,
  -35.3449,
  -35.3885,
  -35.4323,
  -35.4766,
  -35.5212,
  -35.5663,
  -35.612,
  -35.6581,
  -35.7047,
  -35.7518,
  -35.7995,
  -35.848,
  -35.897,
  -35.9465,
  -35.9958,
  -36.0468,
  -36.099,
  -36.1521,
  -36.2052,
  -36.2577,
  -36.3092,
  -36.3596,
  -36.4088,
  -36.4572,
  -36.5048,
  -36.5517,
  -36.5974,
  -36.6424,
  -36.6867,
  -36.7304,
  -36.7735,
  -36.816,
  -36.8567,
  -36.8975,
  -36.9378,
  -36.9782,
  -37.0188,
  -37.0595,
  -37.1001,
  -37.1399,
  -37.1787,
  -37.2167,
  -37.254,
  -37.2908,
  -37.3268,
  -37.3617,
  -37.3948,
  -37.4257,
  -37.4542,
  -37.4809,
  -37.5054,
  -37.5305,
  -37.5552,
  -37.5794,
  -37.6032,
  -37.6263,
  -37.6484,
  -37.6694,
  -37.6891,
  -37.7076,
  -37.7251,
  -37.7421,
  -37.7591,
  -37.7764,
  -37.7938,
  -37.8106,
  -37.8268,
  -37.8424,
  -37.8581,
  -37.8743,
  -37.8904,
  -37.9088,
  -37.9285,
  -37.9499,
  -37.9732,
  -37.9982,
  -38.0241,
  -38.0501,
  -38.0757,
  -38.1004,
  -38.1244,
  -38.1477,
  -38.1706,
  -38.1931,
  -38.2154,
  -38.2377,
  -38.2596,
  -38.2822,
  -38.3057,
  -38.3302,
  -38.3555,
  -38.38,
  -38.405,
  -38.4291,
  -38.4522,
  -38.4741,
  -38.4949,
  -38.5146,
  -38.5336,
  -38.5523,
  -38.571,
  -38.5902,
  -38.6101,
  -38.6307,
  -38.6521,
  -38.6742,
  -38.6964,
  -38.7186,
  -38.7403,
  -38.7611,
  -38.7811,
  -38.801,
  -38.8218,
  -38.844,
  -38.8671,
  -38.8934,
  -38.9212,
  -38.9502,
  -38.9802,
  -39.0105,
  -39.0411,
  -39.0717,
  -39.1019,
  -39.1315,
  -39.1605,
  -39.1891,
  -39.2179,
  -39.2472,
  -39.2772,
  -39.3074,
  -39.3368,
  -39.3645,
  -39.3904,
  -39.4151,
  -39.4388,
  -39.462,
  -39.4847,
  -39.5071,
  -39.5295,
  -39.5516,
  -39.5724,
  -39.5938,
  -39.614,
  -39.6325,
  -39.6491,
  -39.6637,
  -39.6762,
  -39.6867,
  -39.6954,
  -39.7023,
  -39.7077,
  -39.7119,
  -39.715,
  -39.7171,
  -39.7182,
  -39.7182,
  -39.7166,
  -39.7132,
  -39.708,
  -39.7013,
  -39.6942,
  -39.6877,
  -39.683,
  -39.6812,
  -39.6841,
  -39.6928,
  -39.7084,
  -39.7311,
  -39.7605,
  -39.7946,
  -39.834,
  -39.8755,
  -39.9177,
  -39.9589,
  -39.9982,
  -40.035,
  -40.0693,
  -40.1016,
  -40.1322,
  -40.1614,
  -40.1898,
  -40.2173,
  -40.244,
  -40.2691,
  -40.2926,
  -40.3144,
  -40.3347,
  -40.3539,
  -40.3722,
  -40.3904,
  -40.4082,
  -40.426,
  -40.4432,
  -40.4598,
  -40.4748,
  -40.4883,
  -40.5,
  -40.5101,
  -40.5192,
  -40.5278,
  -40.5363,
  -40.5455,
  -40.5551,
  -40.5654,
  -40.5752,
  -40.5865,
  -40.5983,
  -40.61,
  -40.6212,
  -40.6314,
  -40.6399,
  -40.6468,
  -40.6524,
  -40.6566,
  -40.66,
  -40.6627,
  -40.665,
  -40.6665,
  -40.6669,
  -40.6657,
  -40.6627,
  -40.6574,
  -40.65,
  -40.6403,
  -40.6283,
  -40.6144,
  -40.5983,
  -40.5806,
  -40.5611,
  -40.5395,
  -40.5147,
  -40.4857,
  -40.4517,
  -40.4119,
  -40.3662,
  -40.3151,
  -40.2587,
  -40.1983,
  -40.134,
  -40.0664,
  -39.9954,
  -39.9204,
  -39.8405,
  -39.7552,
  -32.7761,
  -32.8232,
  -32.8696,
  -32.9146,
  -32.9571,
  -32.9992,
  -33.0402,
  -33.0808,
  -33.1214,
  -33.1622,
  -33.2031,
  -33.2441,
  -33.2851,
  -33.3262,
  -33.3678,
  -33.4106,
  -33.4547,
  -33.5,
  -33.5451,
  -33.5914,
  -33.6375,
  -33.6833,
  -33.7288,
  -33.7744,
  -33.8201,
  -33.8658,
  -33.9114,
  -33.9568,
  -34.0017,
  -34.0462,
  -34.0899,
  -34.1327,
  -34.1744,
  -34.2142,
  -34.2549,
  -34.2963,
  -34.3387,
  -34.3825,
  -34.4273,
  -34.4727,
  -34.5182,
  -34.5635,
  -34.6086,
  -34.653,
  -34.6966,
  -34.7393,
  -34.7815,
  -34.8236,
  -34.8658,
  -34.9072,
  -34.9496,
  -34.9919,
  -35.0341,
  -35.0763,
  -35.1189,
  -35.1618,
  -35.2053,
  -35.249,
  -35.293,
  -35.3373,
  -35.382,
  -35.4271,
  -35.4728,
  -35.5191,
  -35.566,
  -35.6134,
  -35.6605,
  -35.7092,
  -35.7587,
  -35.8087,
  -35.8591,
  -35.91,
  -35.9616,
  -36.0142,
  -36.0674,
  -36.1209,
  -36.1739,
  -36.226,
  -36.277,
  -36.327,
  -36.3761,
  -36.4243,
  -36.4716,
  -36.5169,
  -36.5623,
  -36.607,
  -36.6513,
  -36.695,
  -36.7382,
  -36.7804,
  -36.8216,
  -36.8619,
  -36.9021,
  -36.9424,
  -36.9829,
  -37.0234,
  -37.0634,
  -37.1027,
  -37.1413,
  -37.1793,
  -37.2165,
  -37.2519,
  -37.2868,
  -37.3197,
  -37.3503,
  -37.3785,
  -37.4047,
  -37.4297,
  -37.454,
  -37.4782,
  -37.5021,
  -37.5257,
  -37.5488,
  -37.5712,
  -37.5925,
  -37.6127,
  -37.6315,
  -37.6492,
  -37.6664,
  -37.6834,
  -37.6997,
  -37.7169,
  -37.7337,
  -37.7499,
  -37.7658,
  -37.7818,
  -37.7985,
  -37.8163,
  -37.8353,
  -37.8557,
  -37.8777,
  -37.9014,
  -37.9268,
  -37.9531,
  -37.9795,
  -38.0056,
  -38.031,
  -38.0555,
  -38.0795,
  -38.1028,
  -38.1255,
  -38.1468,
  -38.1686,
  -38.1905,
  -38.2128,
  -38.236,
  -38.2603,
  -38.2854,
  -38.3109,
  -38.3363,
  -38.361,
  -38.385,
  -38.408,
  -38.4299,
  -38.4507,
  -38.4705,
  -38.4897,
  -38.5089,
  -38.5284,
  -38.5486,
  -38.5697,
  -38.5918,
  -38.6148,
  -38.6372,
  -38.6604,
  -38.6828,
  -38.7041,
  -38.7244,
  -38.7442,
  -38.7646,
  -38.7863,
  -38.8101,
  -38.8358,
  -38.8635,
  -38.8926,
  -38.923,
  -38.954,
  -38.9853,
  -39.0165,
  -39.0469,
  -39.0764,
  -39.1051,
  -39.1333,
  -39.1616,
  -39.1905,
  -39.2198,
  -39.2492,
  -39.2779,
  -39.304,
  -39.3297,
  -39.354,
  -39.3775,
  -39.4005,
  -39.4233,
  -39.4461,
  -39.4688,
  -39.4912,
  -39.5133,
  -39.5346,
  -39.5545,
  -39.5726,
  -39.5888,
  -39.603,
  -39.6155,
  -39.6263,
  -39.6353,
  -39.6429,
  -39.6489,
  -39.6537,
  -39.6572,
  -39.6597,
  -39.6611,
  -39.6612,
  -39.6597,
  -39.6563,
  -39.6511,
  -39.6437,
  -39.6367,
  -39.6306,
  -39.6265,
  -39.6261,
  -39.6308,
  -39.6418,
  -39.6595,
  -39.6842,
  -39.7153,
  -39.7516,
  -39.7916,
  -39.8336,
  -39.8762,
  -39.9177,
  -39.9573,
  -39.9943,
  -40.0289,
  -40.0613,
  -40.0921,
  -40.1218,
  -40.1506,
  -40.1784,
  -40.2052,
  -40.2305,
  -40.2545,
  -40.2768,
  -40.2977,
  -40.3173,
  -40.336,
  -40.354,
  -40.3717,
  -40.3891,
  -40.405,
  -40.4211,
  -40.4358,
  -40.4489,
  -40.4604,
  -40.4704,
  -40.4794,
  -40.488,
  -40.4965,
  -40.5054,
  -40.5147,
  -40.5244,
  -40.5348,
  -40.5457,
  -40.557,
  -40.5685,
  -40.5794,
  -40.5892,
  -40.5976,
  -40.6042,
  -40.6094,
  -40.6133,
  -40.6163,
  -40.6186,
  -40.6203,
  -40.6215,
  -40.6214,
  -40.6197,
  -40.616,
  -40.6102,
  -40.6022,
  -40.5919,
  -40.5794,
  -40.5648,
  -40.5483,
  -40.5303,
  -40.5107,
  -40.4891,
  -40.4647,
  -40.4366,
  -40.4037,
  -40.3654,
  -40.3205,
  -40.2713,
  -40.2174,
  -40.1594,
  -40.0977,
  -40.0327,
  -39.9642,
  -39.8916,
  -39.8144,
  -39.732,
  -32.673,
  -32.7198,
  -32.7657,
  -32.8106,
  -32.8541,
  -32.8964,
  -32.9378,
  -32.9786,
  -33.0196,
  -33.0605,
  -33.1016,
  -33.1428,
  -33.1843,
  -33.2258,
  -33.2669,
  -33.3103,
  -33.3548,
  -33.4002,
  -33.446,
  -33.4917,
  -33.5369,
  -33.582,
  -33.6272,
  -33.6729,
  -33.719,
  -33.7657,
  -33.8124,
  -33.8588,
  -33.9049,
  -33.9495,
  -33.9943,
  -34.0379,
  -34.0801,
  -34.1213,
  -34.1622,
  -34.2035,
  -34.246,
  -34.2899,
  -34.3347,
  -34.3801,
  -34.4257,
  -34.4712,
  -34.5164,
  -34.5609,
  -34.6035,
  -34.6461,
  -34.688,
  -34.7295,
  -34.771,
  -34.8127,
  -34.8546,
  -34.8966,
  -34.9386,
  -34.9809,
  -35.0235,
  -35.0665,
  -35.1101,
  -35.1541,
  -35.1985,
  -35.2433,
  -35.2876,
  -35.3334,
  -35.3798,
  -35.4267,
  -35.4744,
  -35.5227,
  -35.5719,
  -35.6219,
  -35.6725,
  -35.7236,
  -35.775,
  -35.8266,
  -35.8786,
  -35.9315,
  -35.9851,
  -36.039,
  -36.0925,
  -36.1441,
  -36.1957,
  -36.2462,
  -36.2957,
  -36.3443,
  -36.3918,
  -36.4384,
  -36.4841,
  -36.5292,
  -36.574,
  -36.6185,
  -36.6623,
  -36.7051,
  -36.7467,
  -36.7872,
  -36.8273,
  -36.8673,
  -36.9075,
  -36.9469,
  -36.987,
  -37.0268,
  -37.0658,
  -37.1042,
  -37.1418,
  -37.1781,
  -37.2127,
  -37.2453,
  -37.2757,
  -37.3036,
  -37.3297,
  -37.3544,
  -37.3783,
  -37.4019,
  -37.4255,
  -37.4489,
  -37.4721,
  -37.4947,
  -37.5154,
  -37.5359,
  -37.5553,
  -37.5734,
  -37.5909,
  -37.608,
  -37.6251,
  -37.6423,
  -37.659,
  -37.6753,
  -37.6914,
  -37.7078,
  -37.725,
  -37.7434,
  -37.7629,
  -37.7838,
  -37.8061,
  -37.8302,
  -37.8558,
  -37.8822,
  -37.9077,
  -37.9341,
  -37.9599,
  -37.9852,
  -38.0099,
  -38.0338,
  -38.0569,
  -38.0793,
  -38.1013,
  -38.1231,
  -38.1455,
  -38.1687,
  -38.193,
  -38.2179,
  -38.2433,
  -38.2687,
  -38.2939,
  -38.3186,
  -38.3425,
  -38.3654,
  -38.387,
  -38.4077,
  -38.4266,
  -38.4463,
  -38.4662,
  -38.4869,
  -38.5086,
  -38.5315,
  -38.5554,
  -38.5799,
  -38.6042,
  -38.6276,
  -38.6496,
  -38.6702,
  -38.6901,
  -38.7103,
  -38.7316,
  -38.7547,
  -38.78,
  -38.8075,
  -38.8365,
  -38.867,
  -38.8987,
  -38.9303,
  -38.9618,
  -38.9923,
  -39.0205,
  -39.0488,
  -39.0767,
  -39.1047,
  -39.1331,
  -39.162,
  -39.1909,
  -39.2191,
  -39.246,
  -39.2715,
  -39.2958,
  -39.3192,
  -39.3422,
  -39.3651,
  -39.388,
  -39.4109,
  -39.4335,
  -39.4555,
  -39.4764,
  -39.4957,
  -39.5132,
  -39.5289,
  -39.5428,
  -39.5553,
  -39.5665,
  -39.5762,
  -39.5843,
  -39.59,
  -39.5954,
  -39.5995,
  -39.6024,
  -39.6041,
  -39.6044,
  -39.6031,
  -39.5999,
  -39.595,
  -39.5889,
  -39.5826,
  -39.5773,
  -39.5745,
  -39.576,
  -39.5828,
  -39.5959,
  -39.6158,
  -39.6423,
  -39.6749,
  -39.712,
  -39.7524,
  -39.7946,
  -39.8369,
  -39.8783,
  -39.9178,
  -39.9547,
  -39.9892,
  -40.0216,
  -40.0525,
  -40.0824,
  -40.1115,
  -40.1385,
  -40.1654,
  -40.1912,
  -40.2159,
  -40.239,
  -40.2607,
  -40.2809,
  -40.2998,
  -40.3177,
  -40.335,
  -40.352,
  -40.3681,
  -40.3835,
  -40.3977,
  -40.4104,
  -40.4218,
  -40.4319,
  -40.4412,
  -40.4499,
  -40.4586,
  -40.4673,
  -40.4763,
  -40.4858,
  -40.4955,
  -40.5059,
  -40.5167,
  -40.5274,
  -40.5374,
  -40.5464,
  -40.554,
  -40.5601,
  -40.5649,
  -40.5686,
  -40.5715,
  -40.5735,
  -40.575,
  -40.5756,
  -40.5749,
  -40.5715,
  -40.5671,
  -40.5606,
  -40.5518,
  -40.541,
  -40.5282,
  -40.5134,
  -40.4966,
  -40.4784,
  -40.4588,
  -40.4372,
  -40.4132,
  -40.3857,
  -40.3538,
  -40.317,
  -40.275,
  -40.2281,
  -40.1768,
  -40.1214,
  -40.0624,
  -39.9997,
  -39.9332,
  -39.8624,
  -39.7871,
  -39.707,
  -32.5729,
  -32.6192,
  -32.6648,
  -32.7094,
  -32.7528,
  -32.7955,
  -32.8373,
  -32.8788,
  -32.9202,
  -32.9605,
  -33.0017,
  -33.0429,
  -33.0846,
  -33.1263,
  -33.169,
  -33.2128,
  -33.2574,
  -33.3027,
  -33.348,
  -33.393,
  -33.4375,
  -33.4821,
  -33.5271,
  -33.5729,
  -33.6186,
  -33.6659,
  -33.7135,
  -33.761,
  -33.808,
  -33.8547,
  -33.9007,
  -33.9451,
  -33.9883,
  -34.0302,
  -34.0714,
  -34.113,
  -34.1556,
  -34.1993,
  -34.2439,
  -34.2881,
  -34.3336,
  -34.3789,
  -34.424,
  -34.4687,
  -34.5121,
  -34.5546,
  -34.5961,
  -34.637,
  -34.6778,
  -34.7189,
  -34.7602,
  -34.8019,
  -34.844,
  -34.8863,
  -34.9291,
  -34.9715,
  -35.0154,
  -35.0597,
  -35.1046,
  -35.15,
  -35.196,
  -35.2426,
  -35.2898,
  -35.3376,
  -35.386,
  -35.4352,
  -35.4853,
  -35.5362,
  -35.588,
  -35.6402,
  -35.6924,
  -35.7437,
  -35.7965,
  -35.8501,
  -35.9043,
  -35.9588,
  -36.0128,
  -36.0659,
  -36.1177,
  -36.1684,
  -36.2179,
  -36.2665,
  -36.3142,
  -36.3609,
  -36.4067,
  -36.4524,
  -36.4977,
  -36.5425,
  -36.5871,
  -36.6295,
  -36.6715,
  -36.7124,
  -36.7525,
  -36.7924,
  -36.8324,
  -36.8727,
  -36.9129,
  -36.9529,
  -36.9923,
  -37.0309,
  -37.0685,
  -37.1046,
  -37.1388,
  -37.1709,
  -37.2011,
  -37.229,
  -37.2549,
  -37.2794,
  -37.302,
  -37.3252,
  -37.3484,
  -37.3717,
  -37.3951,
  -37.4178,
  -37.4399,
  -37.4609,
  -37.4805,
  -37.4991,
  -37.5168,
  -37.5342,
  -37.5514,
  -37.5686,
  -37.5855,
  -37.6021,
  -37.6186,
  -37.6355,
  -37.6533,
  -37.671,
  -37.6909,
  -37.712,
  -37.7345,
  -37.7586,
  -37.7841,
  -37.8104,
  -37.8369,
  -37.8634,
  -37.8896,
  -37.9155,
  -37.9409,
  -37.9655,
  -37.9893,
  -38.0123,
  -38.0347,
  -38.0571,
  -38.0799,
  -38.1034,
  -38.1276,
  -38.1524,
  -38.1775,
  -38.2017,
  -38.227,
  -38.252,
  -38.2765,
  -38.3001,
  -38.3225,
  -38.3439,
  -38.3646,
  -38.3849,
  -38.4056,
  -38.427,
  -38.4492,
  -38.4729,
  -38.4977,
  -38.5232,
  -38.5485,
  -38.5728,
  -38.5956,
  -38.6169,
  -38.6372,
  -38.6573,
  -38.6782,
  -38.7007,
  -38.7244,
  -38.7513,
  -38.7806,
  -38.8112,
  -38.8431,
  -38.8753,
  -38.9068,
  -38.9369,
  -38.966,
  -38.994,
  -39.0216,
  -39.0493,
  -39.0776,
  -39.1062,
  -39.1347,
  -39.1627,
  -39.1898,
  -39.2155,
  -39.2399,
  -39.2634,
  -39.2864,
  -39.3092,
  -39.3321,
  -39.3549,
  -39.3773,
  -39.3989,
  -39.4182,
  -39.4368,
  -39.4536,
  -39.4688,
  -39.4826,
  -39.4952,
  -39.5066,
  -39.5167,
  -39.5255,
  -39.5327,
  -39.5387,
  -39.5435,
  -39.5469,
  -39.5489,
  -39.5496,
  -39.5486,
  -39.5458,
  -39.5415,
  -39.5362,
  -39.5309,
  -39.5269,
  -39.5259,
  -39.5294,
  -39.5384,
  -39.5538,
  -39.5758,
  -39.604,
  -39.6376,
  -39.6754,
  -39.715,
  -39.7569,
  -39.7989,
  -39.8396,
  -39.8784,
  -39.9149,
  -39.9491,
  -39.9816,
  -40.0126,
  -40.0424,
  -40.0713,
  -40.0995,
  -40.1266,
  -40.1529,
  -40.1785,
  -40.2025,
  -40.225,
  -40.2458,
  -40.265,
  -40.2827,
  -40.2995,
  -40.3157,
  -40.331,
  -40.3456,
  -40.3591,
  -40.3715,
  -40.3828,
  -40.3932,
  -40.4028,
  -40.4119,
  -40.4207,
  -40.4294,
  -40.4383,
  -40.4474,
  -40.4568,
  -40.4655,
  -40.4753,
  -40.485,
  -40.4938,
  -40.5017,
  -40.5084,
  -40.5139,
  -40.5183,
  -40.5218,
  -40.5245,
  -40.5265,
  -40.5277,
  -40.528,
  -40.5267,
  -40.5236,
  -40.5184,
  -40.5112,
  -40.5018,
  -40.4905,
  -40.4774,
  -40.4626,
  -40.4459,
  -40.4277,
  -40.4077,
  -40.3862,
  -40.3625,
  -40.3356,
  -40.3049,
  -40.2695,
  -40.2294,
  -40.1848,
  -40.1359,
  -40.0829,
  -40.0261,
  -39.9651,
  -39.9002,
  -39.8309,
  -39.7566,
  -39.6777,
  -32.4751,
  -32.5207,
  -32.5658,
  -32.6099,
  -32.6523,
  -32.6951,
  -32.7377,
  -32.78,
  -32.822,
  -32.8637,
  -32.9053,
  -32.9466,
  -32.9882,
  -33.0302,
  -33.0731,
  -33.1169,
  -33.1616,
  -33.2065,
  -33.2513,
  -33.2946,
  -33.3385,
  -33.3827,
  -33.4277,
  -33.4737,
  -33.5208,
  -33.5686,
  -33.6169,
  -33.665,
  -33.7129,
  -33.7606,
  -33.8075,
  -33.8532,
  -33.8972,
  -33.9401,
  -33.9811,
  -34.0231,
  -34.0658,
  -34.1094,
  -34.1537,
  -34.1985,
  -34.2435,
  -34.2887,
  -34.3337,
  -34.3779,
  -34.4214,
  -34.4637,
  -34.505,
  -34.5456,
  -34.5858,
  -34.6261,
  -34.666,
  -34.7075,
  -34.7496,
  -34.7921,
  -34.8353,
  -34.879,
  -34.9233,
  -34.9682,
  -35.0138,
  -35.06,
  -35.1068,
  -35.1543,
  -35.2023,
  -35.2509,
  -35.3,
  -35.3498,
  -35.3996,
  -35.4514,
  -35.5041,
  -35.5568,
  -35.6098,
  -35.6633,
  -35.7169,
  -35.7715,
  -35.8266,
  -35.882,
  -35.9366,
  -35.99,
  -36.0418,
  -36.0922,
  -36.1415,
  -36.1898,
  -36.2373,
  -36.283,
  -36.3292,
  -36.3751,
  -36.421,
  -36.4668,
  -36.5114,
  -36.5555,
  -36.5981,
  -36.6394,
  -36.6798,
  -36.7197,
  -36.7598,
  -36.7998,
  -36.8398,
  -36.8798,
  -36.9194,
  -36.9581,
  -36.9956,
  -37.0304,
  -37.0643,
  -37.0963,
  -37.1261,
  -37.1537,
  -37.1795,
  -37.2039,
  -37.2272,
  -37.2501,
  -37.2732,
  -37.2965,
  -37.3197,
  -37.3426,
  -37.3647,
  -37.386,
  -37.4059,
  -37.4249,
  -37.4431,
  -37.4608,
  -37.4784,
  -37.4949,
  -37.5121,
  -37.5292,
  -37.5463,
  -37.5639,
  -37.5822,
  -37.6014,
  -37.6214,
  -37.6425,
  -37.6649,
  -37.6888,
  -37.714,
  -37.74,
  -37.7664,
  -37.793,
  -37.8196,
  -37.8462,
  -37.8723,
  -37.8977,
  -37.9223,
  -37.945,
  -37.9682,
  -37.9914,
  -38.0148,
  -38.0387,
  -38.063,
  -38.0877,
  -38.1125,
  -38.1375,
  -38.1626,
  -38.1876,
  -38.2124,
  -38.2364,
  -38.2595,
  -38.2816,
  -38.3031,
  -38.3243,
  -38.3458,
  -38.3679,
  -38.3906,
  -38.4149,
  -38.4405,
  -38.4667,
  -38.4917,
  -38.5169,
  -38.5406,
  -38.5628,
  -38.5837,
  -38.6039,
  -38.6245,
  -38.6465,
  -38.6705,
  -38.6971,
  -38.7263,
  -38.7574,
  -38.7895,
  -38.8218,
  -38.8531,
  -38.8833,
  -38.9122,
  -38.94,
  -38.9674,
  -38.9949,
  -39.0231,
  -39.0515,
  -39.0798,
  -39.1079,
  -39.1353,
  -39.1605,
  -39.1853,
  -39.209,
  -39.2319,
  -39.2545,
  -39.277,
  -39.2993,
  -39.3213,
  -39.3421,
  -39.3615,
  -39.3793,
  -39.3955,
  -39.4104,
  -39.4242,
  -39.4369,
  -39.4486,
  -39.4592,
  -39.4682,
  -39.4761,
  -39.4828,
  -39.4881,
  -39.4923,
  -39.4948,
  -39.4958,
  -39.4953,
  -39.4931,
  -39.4895,
  -39.4852,
  -39.4803,
  -39.4782,
  -39.4794,
  -39.4852,
  -39.4966,
  -39.5141,
  -39.5377,
  -39.5671,
  -39.6015,
  -39.6398,
  -39.6805,
  -39.7222,
  -39.7635,
  -39.8033,
  -39.8412,
  -39.8771,
  -39.911,
  -39.9433,
  -39.9741,
  -40.0037,
  -40.0324,
  -40.0603,
  -40.0878,
  -40.1148,
  -40.1413,
  -40.1663,
  -40.1896,
  -40.2109,
  -40.2303,
  -40.2478,
  -40.2641,
  -40.2792,
  -40.2934,
  -40.306,
  -40.3189,
  -40.3311,
  -40.3425,
  -40.3532,
  -40.3631,
  -40.3725,
  -40.3815,
  -40.3904,
  -40.3992,
  -40.4082,
  -40.4171,
  -40.4261,
  -40.4349,
  -40.4433,
  -40.451,
  -40.4577,
  -40.4634,
  -40.4683,
  -40.4723,
  -40.4756,
  -40.4781,
  -40.4799,
  -40.4811,
  -40.481,
  -40.4792,
  -40.4755,
  -40.4696,
  -40.4616,
  -40.4516,
  -40.44,
  -40.4266,
  -40.4118,
  -40.3951,
  -40.3769,
  -40.3573,
  -40.3359,
  -40.3123,
  -40.286,
  -40.2562,
  -40.2222,
  -40.1838,
  -40.1401,
  -40.0934,
  -40.0423,
  -39.9871,
  -39.9276,
  -39.8635,
  -39.7946,
  -39.7211,
  -39.6429,
  -32.3782,
  -32.4233,
  -32.4677,
  -32.5115,
  -32.5548,
  -32.5978,
  -32.6409,
  -32.684,
  -32.7268,
  -32.7692,
  -32.811,
  -32.8526,
  -32.8943,
  -32.9364,
  -32.9783,
  -33.0222,
  -33.0665,
  -33.111,
  -33.1551,
  -33.1989,
  -33.2425,
  -33.2865,
  -33.3313,
  -33.3778,
  -33.4252,
  -33.4733,
  -33.522,
  -33.5707,
  -33.6191,
  -33.6664,
  -33.714,
  -33.7606,
  -33.8057,
  -33.8495,
  -33.8925,
  -33.935,
  -33.9779,
  -34.0215,
  -34.0655,
  -34.11,
  -34.1548,
  -34.1996,
  -34.2441,
  -34.2883,
  -34.3304,
  -34.3726,
  -34.4138,
  -34.4541,
  -34.494,
  -34.5339,
  -34.5745,
  -34.6157,
  -34.6578,
  -34.7006,
  -34.7441,
  -34.7883,
  -34.8332,
  -34.8789,
  -34.9253,
  -34.9724,
  -35.0201,
  -35.0675,
  -35.1162,
  -35.1654,
  -35.2151,
  -35.2655,
  -35.3167,
  -35.3689,
  -35.4222,
  -35.4755,
  -35.5296,
  -35.5838,
  -35.6385,
  -35.6944,
  -35.7506,
  -35.8067,
  -35.8618,
  -35.9142,
  -35.9659,
  -36.016,
  -36.0649,
  -36.1129,
  -36.1602,
  -36.2071,
  -36.2536,
  -36.2999,
  -36.3463,
  -36.3927,
  -36.4382,
  -36.4824,
  -36.526,
  -36.5677,
  -36.6083,
  -36.6484,
  -36.6883,
  -36.7269,
  -36.767,
  -36.8068,
  -36.846,
  -36.8845,
  -36.9219,
  -36.9575,
  -36.9913,
  -37.023,
  -37.0526,
  -37.0802,
  -37.1059,
  -37.1301,
  -37.1533,
  -37.176,
  -37.1988,
  -37.2219,
  -37.2451,
  -37.2679,
  -37.2891,
  -37.3102,
  -37.3306,
  -37.35,
  -37.3687,
  -37.387,
  -37.4051,
  -37.423,
  -37.4408,
  -37.4585,
  -37.4764,
  -37.4948,
  -37.5137,
  -37.5333,
  -37.5534,
  -37.5744,
  -37.5965,
  -37.6201,
  -37.645,
  -37.6707,
  -37.6971,
  -37.7228,
  -37.7497,
  -37.7768,
  -37.8037,
  -37.8299,
  -37.8554,
  -37.8799,
  -37.9038,
  -37.9277,
  -37.9517,
  -37.9761,
  -38.0007,
  -38.0254,
  -38.0501,
  -38.0749,
  -38.0999,
  -38.1249,
  -38.1497,
  -38.1741,
  -38.1977,
  -38.2206,
  -38.2419,
  -38.2639,
  -38.2859,
  -38.3087,
  -38.3321,
  -38.3564,
  -38.3824,
  -38.4088,
  -38.4354,
  -38.4614,
  -38.4862,
  -38.5094,
  -38.5311,
  -38.5519,
  -38.5724,
  -38.5938,
  -38.6174,
  -38.644,
  -38.6731,
  -38.7042,
  -38.7366,
  -38.7689,
  -38.8002,
  -38.8304,
  -38.8582,
  -38.8859,
  -38.9133,
  -38.9407,
  -38.9686,
  -38.9969,
  -39.0257,
  -39.0539,
  -39.0816,
  -39.1081,
  -39.1335,
  -39.1574,
  -39.1802,
  -39.2024,
  -39.2243,
  -39.2458,
  -39.2667,
  -39.2866,
  -39.3052,
  -39.3222,
  -39.338,
  -39.3526,
  -39.3662,
  -39.3791,
  -39.3909,
  -39.4018,
  -39.4115,
  -39.4191,
  -39.4265,
  -39.4326,
  -39.4374,
  -39.4407,
  -39.4423,
  -39.4423,
  -39.4408,
  -39.4383,
  -39.4354,
  -39.4332,
  -39.4332,
  -39.4367,
  -39.4449,
  -39.4586,
  -39.4779,
  -39.5028,
  -39.5331,
  -39.5681,
  -39.6066,
  -39.6472,
  -39.6884,
  -39.729,
  -39.768,
  -39.8051,
  -39.8404,
  -39.8739,
  -39.9058,
  -39.9364,
  -39.9657,
  -39.9941,
  -40.021,
  -40.0486,
  -40.0763,
  -40.1033,
  -40.1292,
  -40.1531,
  -40.1751,
  -40.1946,
  -40.2119,
  -40.2273,
  -40.2414,
  -40.2546,
  -40.2673,
  -40.2796,
  -40.2916,
  -40.3033,
  -40.3143,
  -40.3246,
  -40.3344,
  -40.3437,
  -40.3528,
  -40.3618,
  -40.3704,
  -40.3788,
  -40.387,
  -40.3947,
  -40.4021,
  -40.4086,
  -40.4143,
  -40.4191,
  -40.4234,
  -40.4269,
  -40.4299,
  -40.4322,
  -40.4339,
  -40.4348,
  -40.4345,
  -40.4322,
  -40.4276,
  -40.4199,
  -40.411,
  -40.4004,
  -40.3882,
  -40.3748,
  -40.3599,
  -40.3437,
  -40.326,
  -40.3066,
  -40.2855,
  -40.262,
  -40.2361,
  -40.207,
  -40.1742,
  -40.1371,
  -40.096,
  -40.0506,
  -40.001,
  -39.9468,
  -39.888,
  -39.8242,
  -39.7556,
  -39.6821,
  -39.6042,
  -32.2844,
  -32.329,
  -32.3727,
  -32.4159,
  -32.459,
  -32.5022,
  -32.5457,
  -32.5895,
  -32.6332,
  -32.6753,
  -32.7178,
  -32.7598,
  -32.8016,
  -32.844,
  -32.887,
  -32.9305,
  -32.9745,
  -33.0184,
  -33.0619,
  -33.1052,
  -33.1484,
  -33.1923,
  -33.2374,
  -33.2839,
  -33.3305,
  -33.3789,
  -33.4276,
  -33.4765,
  -33.5253,
  -33.5739,
  -33.6221,
  -33.6694,
  -33.7154,
  -33.7603,
  -33.8041,
  -33.8475,
  -33.8907,
  -33.9342,
  -33.9782,
  -34.0215,
  -34.0658,
  -34.1101,
  -34.154,
  -34.1977,
  -34.2406,
  -34.2829,
  -34.3242,
  -34.3647,
  -34.4045,
  -34.4444,
  -34.4848,
  -34.5261,
  -34.5682,
  -34.6112,
  -34.655,
  -34.6987,
  -34.7443,
  -34.7908,
  -34.8382,
  -34.8863,
  -34.935,
  -34.9839,
  -35.0333,
  -35.0831,
  -35.1333,
  -35.184,
  -35.2356,
  -35.288,
  -35.3414,
  -35.3955,
  -35.45,
  -35.5053,
  -35.5601,
  -35.6171,
  -35.6743,
  -35.7311,
  -35.7865,
  -35.8399,
  -35.8912,
  -35.941,
  -35.9896,
  -36.0374,
  -36.0846,
  -36.1316,
  -36.1782,
  -36.2251,
  -36.2722,
  -36.3191,
  -36.3655,
  -36.4098,
  -36.4537,
  -36.4962,
  -36.5372,
  -36.5772,
  -36.6168,
  -36.6562,
  -36.6958,
  -36.735,
  -36.7742,
  -36.8123,
  -36.8493,
  -36.885,
  -36.9186,
  -36.9503,
  -36.9799,
  -37.0075,
  -37.033,
  -37.0571,
  -37.079,
  -37.1016,
  -37.1243,
  -37.1473,
  -37.1702,
  -37.1929,
  -37.2148,
  -37.2361,
  -37.2566,
  -37.2767,
  -37.2962,
  -37.3152,
  -37.3338,
  -37.3522,
  -37.3705,
  -37.389,
  -37.4078,
  -37.427,
  -37.4466,
  -37.4665,
  -37.4858,
  -37.5067,
  -37.5286,
  -37.552,
  -37.5766,
  -37.6022,
  -37.6285,
  -37.6553,
  -37.6826,
  -37.7102,
  -37.7377,
  -37.7645,
  -37.7904,
  -37.8155,
  -37.8401,
  -37.8645,
  -37.8893,
  -37.9144,
  -37.9394,
  -37.9644,
  -37.9893,
  -38.0131,
  -38.038,
  -38.063,
  -38.088,
  -38.1127,
  -38.1368,
  -38.1604,
  -38.1835,
  -38.2062,
  -38.229,
  -38.2518,
  -38.2753,
  -38.2996,
  -38.3251,
  -38.3517,
  -38.3787,
  -38.4056,
  -38.4315,
  -38.4559,
  -38.4785,
  -38.4999,
  -38.5206,
  -38.5422,
  -38.5643,
  -38.5904,
  -38.6196,
  -38.651,
  -38.6836,
  -38.7158,
  -38.7471,
  -38.7772,
  -38.806,
  -38.8338,
  -38.861,
  -38.8883,
  -38.916,
  -38.9442,
  -38.9733,
  -39.002,
  -39.0301,
  -39.0571,
  -39.0826,
  -39.1066,
  -39.1291,
  -39.1508,
  -39.1719,
  -39.1924,
  -39.2119,
  -39.2306,
  -39.2471,
  -39.2638,
  -39.2791,
  -39.2936,
  -39.3072,
  -39.3201,
  -39.332,
  -39.3431,
  -39.3533,
  -39.3626,
  -39.371,
  -39.3782,
  -39.3841,
  -39.3882,
  -39.3907,
  -39.3914,
  -39.391,
  -39.3897,
  -39.3885,
  -39.3883,
  -39.3906,
  -39.3966,
  -39.4072,
  -39.4226,
  -39.4435,
  -39.4697,
  -39.5006,
  -39.5357,
  -39.5742,
  -39.6145,
  -39.6543,
  -39.6942,
  -39.7324,
  -39.7688,
  -39.8034,
  -39.8366,
  -39.8683,
  -39.8986,
  -39.9276,
  -39.9555,
  -39.9832,
  -40.0108,
  -40.0387,
  -40.0663,
  -40.0926,
  -40.1171,
  -40.1395,
  -40.1592,
  -40.1763,
  -40.1911,
  -40.2043,
  -40.2166,
  -40.2286,
  -40.2406,
  -40.2525,
  -40.2642,
  -40.2755,
  -40.2863,
  -40.2967,
  -40.3065,
  -40.3159,
  -40.3247,
  -40.3329,
  -40.3407,
  -40.348,
  -40.3541,
  -40.3604,
  -40.3659,
  -40.3709,
  -40.3751,
  -40.3787,
  -40.3817,
  -40.3842,
  -40.3862,
  -40.3877,
  -40.3882,
  -40.3873,
  -40.3845,
  -40.3795,
  -40.3721,
  -40.3625,
  -40.3511,
  -40.3384,
  -40.3248,
  -40.3101,
  -40.2943,
  -40.2771,
  -40.2581,
  -40.2372,
  -40.214,
  -40.1884,
  -40.1599,
  -40.1278,
  -40.0916,
  -40.0515,
  -40.0072,
  -39.9583,
  -39.9046,
  -39.846,
  -39.7822,
  -39.7134,
  -39.6396,
  -39.561,
  -32.1923,
  -32.2365,
  -32.2799,
  -32.3226,
  -32.3654,
  -32.4076,
  -32.4514,
  -32.4956,
  -32.5399,
  -32.5837,
  -32.6267,
  -32.6691,
  -32.7115,
  -32.7543,
  -32.7974,
  -32.8409,
  -32.8847,
  -32.9281,
  -32.9711,
  -33.0129,
  -33.0561,
  -33.1,
  -33.1452,
  -33.1917,
  -33.2393,
  -33.2877,
  -33.3365,
  -33.3854,
  -33.4342,
  -33.4829,
  -33.5313,
  -33.579,
  -33.6257,
  -33.6712,
  -33.7145,
  -33.7585,
  -33.8023,
  -33.8462,
  -33.8903,
  -33.9345,
  -33.9784,
  -34.0221,
  -34.0656,
  -34.1087,
  -34.1515,
  -34.1938,
  -34.2352,
  -34.276,
  -34.3162,
  -34.3563,
  -34.3959,
  -34.4372,
  -34.4795,
  -34.5228,
  -34.5671,
  -34.6123,
  -34.6586,
  -34.7059,
  -34.7542,
  -34.8033,
  -34.8526,
  -34.9021,
  -34.9521,
  -35.0023,
  -35.0529,
  -35.1042,
  -35.1552,
  -35.2082,
  -35.262,
  -35.3165,
  -35.3716,
  -35.4274,
  -35.4842,
  -35.5417,
  -35.5996,
  -35.6567,
  -35.7121,
  -35.7651,
  -35.8163,
  -35.866,
  -35.9147,
  -35.9624,
  -36.0096,
  -36.0567,
  -36.103,
  -36.1505,
  -36.1982,
  -36.2457,
  -36.2928,
  -36.339,
  -36.3838,
  -36.4268,
  -36.4681,
  -36.5081,
  -36.5475,
  -36.5866,
  -36.6255,
  -36.6643,
  -36.7028,
  -36.7407,
  -36.7776,
  -36.8132,
  -36.846,
  -36.8778,
  -36.9074,
  -36.9347,
  -36.9601,
  -36.9838,
  -37.0066,
  -37.0291,
  -37.0517,
  -37.0746,
  -37.0974,
  -37.1199,
  -37.1418,
  -37.1631,
  -37.184,
  -37.2046,
  -37.2249,
  -37.2446,
  -37.2639,
  -37.2818,
  -37.3007,
  -37.3198,
  -37.3393,
  -37.3593,
  -37.3795,
  -37.3998,
  -37.4203,
  -37.4413,
  -37.4634,
  -37.4866,
  -37.5113,
  -37.5368,
  -37.5631,
  -37.5902,
  -37.6176,
  -37.6455,
  -37.6732,
  -37.7003,
  -37.7266,
  -37.752,
  -37.7759,
  -37.801,
  -37.8265,
  -37.8523,
  -37.8781,
  -37.9035,
  -37.9286,
  -37.9537,
  -37.9788,
  -38.004,
  -38.0293,
  -38.0544,
  -38.0791,
  -38.1032,
  -38.127,
  -38.1502,
  -38.1731,
  -38.1959,
  -38.2191,
  -38.2431,
  -38.2685,
  -38.295,
  -38.3224,
  -38.3491,
  -38.3762,
  -38.4018,
  -38.4255,
  -38.4477,
  -38.4689,
  -38.4906,
  -38.5141,
  -38.5401,
  -38.5692,
  -38.6001,
  -38.6324,
  -38.6646,
  -38.6958,
  -38.7258,
  -38.7547,
  -38.7825,
  -38.8097,
  -38.8368,
  -38.8644,
  -38.8925,
  -38.9213,
  -38.9503,
  -38.9787,
  -39.005,
  -39.0306,
  -39.0544,
  -39.0767,
  -39.0978,
  -39.118,
  -39.1374,
  -39.1556,
  -39.1733,
  -39.1898,
  -39.2056,
  -39.2208,
  -39.2351,
  -39.2486,
  -39.2615,
  -39.2736,
  -39.2851,
  -39.296,
  -39.3063,
  -39.3159,
  -39.3244,
  -39.3314,
  -39.3366,
  -39.3401,
  -39.342,
  -39.3427,
  -39.3429,
  -39.3435,
  -39.3455,
  -39.3491,
  -39.3574,
  -39.3701,
  -39.3875,
  -39.4098,
  -39.4368,
  -39.4682,
  -39.5032,
  -39.5414,
  -39.5812,
  -39.6214,
  -39.6606,
  -39.6981,
  -39.7339,
  -39.7681,
  -39.801,
  -39.8325,
  -39.8625,
  -39.8912,
  -39.9189,
  -39.9463,
  -39.9738,
  -40.0015,
  -40.0289,
  -40.0554,
  -40.0803,
  -40.1029,
  -40.1227,
  -40.1397,
  -40.1541,
  -40.1667,
  -40.1785,
  -40.1901,
  -40.2008,
  -40.2128,
  -40.2246,
  -40.2362,
  -40.2476,
  -40.2585,
  -40.2688,
  -40.2784,
  -40.2872,
  -40.2951,
  -40.3022,
  -40.3087,
  -40.3146,
  -40.3202,
  -40.3251,
  -40.3293,
  -40.3329,
  -40.336,
  -40.3385,
  -40.3407,
  -40.3424,
  -40.3436,
  -40.3437,
  -40.3423,
  -40.339,
  -40.3334,
  -40.3253,
  -40.3151,
  -40.303,
  -40.2897,
  -40.2757,
  -40.2612,
  -40.2458,
  -40.2292,
  -40.2108,
  -40.1903,
  -40.1673,
  -40.1419,
  -40.1136,
  -40.082,
  -40.0463,
  -40.0067,
  -39.9618,
  -39.9132,
  -39.8598,
  -39.8011,
  -39.7371,
  -39.6677,
  -39.593,
  -39.5135,
  -32.1005,
  -32.1447,
  -32.1879,
  -32.2304,
  -32.273,
  -32.3161,
  -32.36,
  -32.4044,
  -32.449,
  -32.4932,
  -32.5367,
  -32.5797,
  -32.6226,
  -32.6659,
  -32.7094,
  -32.7521,
  -32.7956,
  -32.8389,
  -32.8817,
  -32.9245,
  -32.9677,
  -33.0117,
  -33.0569,
  -33.1032,
  -33.1507,
  -33.199,
  -33.2476,
  -33.2964,
  -33.3451,
  -33.3928,
  -33.4412,
  -33.4887,
  -33.5356,
  -33.5813,
  -33.6261,
  -33.6706,
  -33.7147,
  -33.759,
  -33.8035,
  -33.8477,
  -33.8914,
  -33.9347,
  -33.9777,
  -34.0204,
  -34.0629,
  -34.1042,
  -34.146,
  -34.1872,
  -34.2278,
  -34.2684,
  -34.3092,
  -34.351,
  -34.3937,
  -34.4374,
  -34.4821,
  -34.528,
  -34.5749,
  -34.6231,
  -34.6721,
  -34.7218,
  -34.7718,
  -34.8208,
  -34.871,
  -34.9216,
  -34.9728,
  -35.0247,
  -35.0776,
  -35.1312,
  -35.1858,
  -35.2409,
  -35.2965,
  -35.3529,
  -35.41,
  -35.4678,
  -35.5256,
  -35.5824,
  -35.6374,
  -35.6901,
  -35.7402,
  -35.7901,
  -35.839,
  -35.8871,
  -35.9347,
  -35.9822,
  -36.0299,
  -36.0781,
  -36.1262,
  -36.1743,
  -36.222,
  -36.2688,
  -36.3142,
  -36.3578,
  -36.3995,
  -36.4396,
  -36.4788,
  -36.5175,
  -36.555,
  -36.5934,
  -36.6315,
  -36.6691,
  -36.7059,
  -36.7417,
  -36.7756,
  -36.8074,
  -36.8366,
  -36.8639,
  -36.889,
  -36.9124,
  -36.935,
  -36.9575,
  -36.9801,
  -37.0029,
  -37.0257,
  -37.0482,
  -37.0701,
  -37.0907,
  -37.112,
  -37.1332,
  -37.1541,
  -37.1746,
  -37.1945,
  -37.2139,
  -37.2333,
  -37.253,
  -37.2731,
  -37.2937,
  -37.3145,
  -37.3354,
  -37.3563,
  -37.3777,
  -37.4001,
  -37.4237,
  -37.4483,
  -37.474,
  -37.5004,
  -37.5264,
  -37.554,
  -37.5817,
  -37.6092,
  -37.6364,
  -37.6628,
  -37.6884,
  -37.7138,
  -37.7395,
  -37.7658,
  -37.7923,
  -37.8188,
  -37.8448,
  -37.8705,
  -37.8959,
  -37.9213,
  -37.947,
  -37.9726,
  -37.9981,
  -38.0232,
  -38.0478,
  -38.072,
  -38.0945,
  -38.1174,
  -38.14,
  -38.1629,
  -38.1866,
  -38.2118,
  -38.2385,
  -38.2665,
  -38.2949,
  -38.3232,
  -38.3498,
  -38.3747,
  -38.3977,
  -38.4195,
  -38.4417,
  -38.4654,
  -38.4915,
  -38.5203,
  -38.551,
  -38.5827,
  -38.6146,
  -38.6455,
  -38.6753,
  -38.704,
  -38.7308,
  -38.7579,
  -38.785,
  -38.8124,
  -38.8405,
  -38.8691,
  -38.8979,
  -38.9262,
  -38.9532,
  -38.9785,
  -39.0022,
  -39.0241,
  -39.0447,
  -39.0641,
  -39.0824,
  -39.0996,
  -39.1162,
  -39.1319,
  -39.1472,
  -39.1619,
  -39.176,
  -39.1895,
  -39.2023,
  -39.2145,
  -39.2265,
  -39.2383,
  -39.2499,
  -39.2599,
  -39.2699,
  -39.2784,
  -39.285,
  -39.2899,
  -39.2932,
  -39.2954,
  -39.2972,
  -39.2995,
  -39.3037,
  -39.3105,
  -39.321,
  -39.3356,
  -39.3546,
  -39.378,
  -39.4056,
  -39.4372,
  -39.4724,
  -39.5099,
  -39.549,
  -39.5884,
  -39.6269,
  -39.6639,
  -39.6991,
  -39.7331,
  -39.7658,
  -39.7972,
  -39.8268,
  -39.8554,
  -39.8829,
  -39.91,
  -39.9362,
  -39.9634,
  -39.9905,
  -40.0167,
  -40.0414,
  -40.064,
  -40.0839,
  -40.1009,
  -40.1153,
  -40.1279,
  -40.1395,
  -40.1509,
  -40.1626,
  -40.1746,
  -40.1865,
  -40.1985,
  -40.2102,
  -40.2216,
  -40.2324,
  -40.2422,
  -40.2508,
  -40.2583,
  -40.2647,
  -40.2705,
  -40.2757,
  -40.2805,
  -40.2847,
  -40.2882,
  -40.2913,
  -40.2939,
  -40.296,
  -40.2978,
  -40.2994,
  -40.3003,
  -40.3001,
  -40.2982,
  -40.2944,
  -40.2883,
  -40.2798,
  -40.2681,
  -40.2554,
  -40.2415,
  -40.2273,
  -40.2129,
  -40.198,
  -40.182,
  -40.1641,
  -40.1437,
  -40.1208,
  -40.0952,
  -40.0668,
  -40.0351,
  -39.9997,
  -39.9602,
  -39.9164,
  -39.868,
  -39.8145,
  -39.7557,
  -39.6912,
  -39.6211,
  -39.5453,
  -39.4646,
  -32.0107,
  -32.0552,
  -32.0985,
  -32.1412,
  -32.1839,
  -32.227,
  -32.2708,
  -32.3152,
  -32.3598,
  -32.4042,
  -32.4471,
  -32.4906,
  -32.5341,
  -32.578,
  -32.622,
  -32.666,
  -32.7096,
  -32.7528,
  -32.7957,
  -32.8387,
  -32.882,
  -32.9261,
  -32.9713,
  -33.0174,
  -33.0646,
  -33.1116,
  -33.16,
  -33.2087,
  -33.2573,
  -33.3059,
  -33.3539,
  -33.4012,
  -33.4477,
  -33.4933,
  -33.5382,
  -33.5828,
  -33.6275,
  -33.6722,
  -33.7168,
  -33.761,
  -33.8037,
  -33.8468,
  -33.8895,
  -33.932,
  -33.9743,
  -34.0166,
  -34.0585,
  -34.1001,
  -34.1414,
  -34.1825,
  -34.2239,
  -34.2662,
  -34.3094,
  -34.3538,
  -34.3992,
  -34.4457,
  -34.4923,
  -34.5411,
  -34.5908,
  -34.641,
  -34.6914,
  -34.7417,
  -34.7923,
  -34.8434,
  -34.8952,
  -34.9479,
  -35.0016,
  -35.0562,
  -35.1117,
  -35.1677,
  -35.2241,
  -35.2808,
  -35.3369,
  -35.3947,
  -35.4518,
  -35.5078,
  -35.562,
  -35.6145,
  -35.6656,
  -35.7157,
  -35.7651,
  -35.814,
  -35.8622,
  -35.91,
  -35.9583,
  -36.0068,
  -36.0553,
  -36.1037,
  -36.1516,
  -36.1986,
  -36.2434,
  -36.2875,
  -36.3297,
  -36.3701,
  -36.4094,
  -36.448,
  -36.4863,
  -36.5245,
  -36.5624,
  -36.5997,
  -36.6364,
  -36.6722,
  -36.7061,
  -36.738,
  -36.7668,
  -36.7936,
  -36.8183,
  -36.8417,
  -36.8643,
  -36.8859,
  -36.9087,
  -36.9317,
  -36.9546,
  -36.9772,
  -36.9994,
  -37.0214,
  -37.0431,
  -37.0649,
  -37.0865,
  -37.1075,
  -37.128,
  -37.1478,
  -37.1677,
  -37.1878,
  -37.2084,
  -37.2296,
  -37.251,
  -37.2724,
  -37.293,
  -37.3151,
  -37.3382,
  -37.3622,
  -37.3874,
  -37.4133,
  -37.4397,
  -37.4665,
  -37.4937,
  -37.521,
  -37.5482,
  -37.575,
  -37.6012,
  -37.6272,
  -37.6532,
  -37.6796,
  -37.7066,
  -37.7339,
  -37.761,
  -37.7877,
  -37.8138,
  -37.8398,
  -37.8648,
  -37.8908,
  -37.9167,
  -37.9426,
  -37.968,
  -37.9928,
  -38.0171,
  -38.0409,
  -38.0637,
  -38.0862,
  -38.109,
  -38.1326,
  -38.1579,
  -38.1849,
  -38.2134,
  -38.2429,
  -38.272,
  -38.2999,
  -38.3255,
  -38.3491,
  -38.3718,
  -38.3946,
  -38.4187,
  -38.4438,
  -38.4722,
  -38.5024,
  -38.5334,
  -38.5645,
  -38.5949,
  -38.6245,
  -38.6531,
  -38.6808,
  -38.7079,
  -38.7348,
  -38.762,
  -38.7897,
  -38.818,
  -38.8462,
  -38.8741,
  -38.9005,
  -38.9254,
  -38.9485,
  -38.97,
  -38.9901,
  -39.0089,
  -39.0265,
  -39.0429,
  -39.0586,
  -39.0737,
  -39.0875,
  -39.1018,
  -39.1155,
  -39.1289,
  -39.1418,
  -39.1543,
  -39.167,
  -39.1799,
  -39.1928,
  -39.2055,
  -39.2173,
  -39.2275,
  -39.2359,
  -39.2423,
  -39.2472,
  -39.251,
  -39.2545,
  -39.2588,
  -39.2649,
  -39.2737,
  -39.2861,
  -39.3023,
  -39.3226,
  -39.3469,
  -39.3752,
  -39.4069,
  -39.4416,
  -39.4785,
  -39.5166,
  -39.555,
  -39.5918,
  -39.6281,
  -39.6631,
  -39.6969,
  -39.7295,
  -39.7607,
  -39.7902,
  -39.8186,
  -39.846,
  -39.873,
  -39.8997,
  -39.9264,
  -39.9527,
  -39.9781,
  -40.0022,
  -40.0246,
  -40.0446,
  -40.0618,
  -40.0766,
  -40.0895,
  -40.1014,
  -40.1131,
  -40.125,
  -40.137,
  -40.149,
  -40.161,
  -40.1731,
  -40.1849,
  -40.1959,
  -40.2058,
  -40.2142,
  -40.2211,
  -40.2268,
  -40.2317,
  -40.2362,
  -40.2393,
  -40.243,
  -40.2462,
  -40.2488,
  -40.2509,
  -40.2526,
  -40.2543,
  -40.2558,
  -40.2566,
  -40.2561,
  -40.2539,
  -40.2497,
  -40.2432,
  -40.2343,
  -40.2231,
  -40.2099,
  -40.1957,
  -40.1813,
  -40.1672,
  -40.1527,
  -40.1373,
  -40.1197,
  -40.0993,
  -40.076,
  -40.05,
  -40.0212,
  -39.9892,
  -39.9536,
  -39.9138,
  -39.8698,
  -39.8213,
  -39.7678,
  -39.7088,
  -39.644,
  -39.573,
  -39.4962,
  -39.4143,
  -31.9221,
  -31.9671,
  -32.011,
  -32.0541,
  -32.097,
  -32.1391,
  -32.1828,
  -32.227,
  -32.2714,
  -32.3159,
  -32.36,
  -32.404,
  -32.4481,
  -32.4924,
  -32.537,
  -32.5814,
  -32.6253,
  -32.6687,
  -32.7119,
  -32.755,
  -32.7975,
  -32.8416,
  -32.8866,
  -32.9326,
  -32.9795,
  -33.0273,
  -33.0756,
  -33.1241,
  -33.1725,
  -33.2207,
  -33.2684,
  -33.3153,
  -33.3613,
  -33.4066,
  -33.4515,
  -33.4952,
  -33.5401,
  -33.585,
  -33.6297,
  -33.6739,
  -33.7175,
  -33.7606,
  -33.8033,
  -33.8458,
  -33.8881,
  -33.9303,
  -33.9725,
  -34.0145,
  -34.0563,
  -34.0981,
  -34.1393,
  -34.1823,
  -34.2262,
  -34.2713,
  -34.3174,
  -34.3645,
  -34.4128,
  -34.4621,
  -34.5123,
  -34.5628,
  -34.6134,
  -34.6641,
  -34.715,
  -34.7665,
  -34.8189,
  -34.8724,
  -34.9271,
  -34.9818,
  -35.0384,
  -35.0954,
  -35.1525,
  -35.2098,
  -35.267,
  -35.324,
  -35.3804,
  -35.4355,
  -35.4889,
  -35.541,
  -35.5921,
  -35.6427,
  -35.6927,
  -35.7421,
  -35.7908,
  -35.8392,
  -35.8867,
  -35.9353,
  -35.9839,
  -36.0322,
  -36.0799,
  -36.1269,
  -36.1729,
  -36.2174,
  -36.2602,
  -36.3012,
  -36.3409,
  -36.3797,
  -36.4182,
  -36.4562,
  -36.4939,
  -36.531,
  -36.5673,
  -36.6027,
  -36.6356,
  -36.6672,
  -36.6962,
  -36.7228,
  -36.7474,
  -36.7707,
  -36.7936,
  -36.8166,
  -36.8397,
  -36.863,
  -36.8861,
  -36.909,
  -36.9316,
  -36.9539,
  -36.9762,
  -36.9985,
  -37.0206,
  -37.0421,
  -37.063,
  -37.0833,
  -37.1026,
  -37.1233,
  -37.1445,
  -37.1662,
  -37.1883,
  -37.2105,
  -37.2329,
  -37.2557,
  -37.2794,
  -37.3042,
  -37.3297,
  -37.3559,
  -37.3823,
  -37.4089,
  -37.4357,
  -37.4624,
  -37.489,
  -37.5153,
  -37.5415,
  -37.5677,
  -37.5942,
  -37.6204,
  -37.6482,
  -37.6762,
  -37.704,
  -37.7313,
  -37.7581,
  -37.7847,
  -37.8111,
  -37.8374,
  -37.8636,
  -37.8895,
  -37.915,
  -37.9401,
  -37.9645,
  -37.9882,
  -38.0111,
  -38.0338,
  -38.0567,
  -38.0806,
  -38.1063,
  -38.1337,
  -38.1628,
  -38.1918,
  -38.2215,
  -38.2499,
  -38.2763,
  -38.3008,
  -38.3243,
  -38.3479,
  -38.3727,
  -38.399,
  -38.4269,
  -38.4562,
  -38.4864,
  -38.5166,
  -38.5464,
  -38.5756,
  -38.604,
  -38.6315,
  -38.6585,
  -38.6851,
  -38.712,
  -38.7393,
  -38.7669,
  -38.7944,
  -38.8213,
  -38.847,
  -38.8702,
  -38.8928,
  -38.9139,
  -38.9336,
  -38.9521,
  -38.9692,
  -38.9851,
  -39.0001,
  -39.0146,
  -39.0289,
  -39.0428,
  -39.0563,
  -39.0694,
  -39.0823,
  -39.0955,
  -39.109,
  -39.1231,
  -39.1375,
  -39.1518,
  -39.1653,
  -39.1775,
  -39.1879,
  -39.1963,
  -39.203,
  -39.2086,
  -39.214,
  -39.22,
  -39.2279,
  -39.2376,
  -39.2515,
  -39.269,
  -39.2902,
  -39.3152,
  -39.3437,
  -39.3754,
  -39.4097,
  -39.4458,
  -39.4831,
  -39.5205,
  -39.5575,
  -39.5934,
  -39.6282,
  -39.6618,
  -39.6942,
  -39.7252,
  -39.7547,
  -39.783,
  -39.8103,
  -39.837,
  -39.8633,
  -39.8892,
  -39.9145,
  -39.9389,
  -39.9623,
  -39.9841,
  -40.0041,
  -40.0217,
  -40.037,
  -40.0507,
  -40.0633,
  -40.0755,
  -40.0875,
  -40.0986,
  -40.1105,
  -40.1225,
  -40.1345,
  -40.1464,
  -40.1576,
  -40.1676,
  -40.1758,
  -40.1825,
  -40.1878,
  -40.1922,
  -40.1961,
  -40.1996,
  -40.2027,
  -40.2052,
  -40.2072,
  -40.2089,
  -40.2104,
  -40.212,
  -40.2134,
  -40.2141,
  -40.2135,
  -40.2111,
  -40.2065,
  -40.1996,
  -40.1904,
  -40.1789,
  -40.1654,
  -40.151,
  -40.1367,
  -40.1228,
  -40.1088,
  -40.0936,
  -40.0758,
  -40.0549,
  -40.031,
  -40.0043,
  -39.9748,
  -39.9422,
  -39.906,
  -39.8659,
  -39.8216,
  -39.7729,
  -39.7183,
  -39.6592,
  -39.594,
  -39.5223,
  -39.4445,
  -39.3617,
  -31.8346,
  -31.8791,
  -31.9239,
  -31.9677,
  -32.0111,
  -32.0544,
  -32.0979,
  -32.1418,
  -32.1861,
  -32.2305,
  -32.2749,
  -32.3192,
  -32.3638,
  -32.4085,
  -32.4534,
  -32.4973,
  -32.5415,
  -32.5853,
  -32.6288,
  -32.6722,
  -32.716,
  -32.7601,
  -32.8048,
  -32.8506,
  -32.8972,
  -32.9448,
  -32.9931,
  -33.0416,
  -33.09,
  -33.138,
  -33.1842,
  -33.2306,
  -33.2762,
  -33.3212,
  -33.3659,
  -33.4106,
  -33.4554,
  -33.5001,
  -33.5444,
  -33.5885,
  -33.6322,
  -33.6755,
  -33.7185,
  -33.7611,
  -33.8036,
  -33.8449,
  -33.8871,
  -33.9293,
  -33.9716,
  -34.0143,
  -34.0575,
  -34.1014,
  -34.1462,
  -34.1919,
  -34.2387,
  -34.2865,
  -34.3354,
  -34.3852,
  -34.4357,
  -34.4864,
  -34.5371,
  -34.588,
  -34.6382,
  -34.6903,
  -34.7433,
  -34.7978,
  -34.8535,
  -34.9105,
  -34.9682,
  -35.0263,
  -35.0843,
  -35.1421,
  -35.1991,
  -35.2555,
  -35.311,
  -35.365,
  -35.4176,
  -35.4694,
  -35.5197,
  -35.5706,
  -35.6215,
  -35.6713,
  -35.7204,
  -35.7695,
  -35.8177,
  -35.8661,
  -35.9143,
  -35.9623,
  -36.0093,
  -36.0559,
  -36.1018,
  -36.1467,
  -36.1901,
  -36.232,
  -36.2724,
  -36.3118,
  -36.3495,
  -36.3879,
  -36.4253,
  -36.4622,
  -36.498,
  -36.5328,
  -36.5663,
  -36.5975,
  -36.6265,
  -36.6531,
  -36.6778,
  -36.7017,
  -36.7251,
  -36.7487,
  -36.7724,
  -36.7962,
  -36.8198,
  -36.8432,
  -36.8662,
  -36.8879,
  -36.9106,
  -36.9331,
  -36.9555,
  -36.9772,
  -36.9985,
  -37.0194,
  -37.0402,
  -37.0613,
  -37.0831,
  -37.1055,
  -37.1284,
  -37.1516,
  -37.175,
  -37.1988,
  -37.2233,
  -37.2486,
  -37.2746,
  -37.3009,
  -37.3273,
  -37.3538,
  -37.3791,
  -37.4051,
  -37.4309,
  -37.4566,
  -37.4826,
  -37.509,
  -37.5361,
  -37.564,
  -37.5924,
  -37.6211,
  -37.6495,
  -37.6774,
  -37.7049,
  -37.7321,
  -37.7589,
  -37.7853,
  -37.8114,
  -37.8372,
  -37.8628,
  -37.8879,
  -37.9122,
  -37.9358,
  -37.9583,
  -37.9814,
  -38.0049,
  -38.0296,
  -38.0559,
  -38.0839,
  -38.1135,
  -38.1438,
  -38.1739,
  -38.2025,
  -38.2293,
  -38.2545,
  -38.2789,
  -38.3034,
  -38.3288,
  -38.3553,
  -38.3829,
  -38.4114,
  -38.4404,
  -38.4697,
  -38.4988,
  -38.5274,
  -38.5555,
  -38.5829,
  -38.6087,
  -38.6351,
  -38.6616,
  -38.6883,
  -38.7152,
  -38.7419,
  -38.7677,
  -38.7924,
  -38.8161,
  -38.838,
  -38.8588,
  -38.8783,
  -38.8965,
  -38.9134,
  -38.929,
  -38.9436,
  -38.9577,
  -38.9714,
  -38.9848,
  -38.998,
  -39.011,
  -39.0241,
  -39.038,
  -39.0523,
  -39.0675,
  -39.0835,
  -39.0992,
  -39.1134,
  -39.1274,
  -39.14,
  -39.1504,
  -39.1592,
  -39.1669,
  -39.174,
  -39.1818,
  -39.1914,
  -39.2035,
  -39.2188,
  -39.2373,
  -39.2592,
  -39.2846,
  -39.3133,
  -39.3447,
  -39.3786,
  -39.4141,
  -39.4504,
  -39.4869,
  -39.5231,
  -39.5585,
  -39.5932,
  -39.6267,
  -39.659,
  -39.6899,
  -39.7192,
  -39.7474,
  -39.7747,
  -39.8013,
  -39.8273,
  -39.8514,
  -39.8755,
  -39.8989,
  -39.9211,
  -39.9422,
  -39.9619,
  -39.98,
  -39.9961,
  -40.0106,
  -40.0241,
  -40.0368,
  -40.0492,
  -40.0613,
  -40.0731,
  -40.0847,
  -40.0966,
  -40.1083,
  -40.1194,
  -40.1294,
  -40.1377,
  -40.1443,
  -40.1494,
  -40.1534,
  -40.1568,
  -40.1597,
  -40.1621,
  -40.1641,
  -40.1656,
  -40.1669,
  -40.1683,
  -40.1699,
  -40.1717,
  -40.1722,
  -40.1715,
  -40.1688,
  -40.1637,
  -40.1564,
  -40.1467,
  -40.1348,
  -40.1203,
  -40.1059,
  -40.0917,
  -40.0779,
  -40.064,
  -40.0485,
  -40.0303,
  -40.0087,
  -39.9839,
  -39.9562,
  -39.9259,
  -39.8925,
  -39.8556,
  -39.8148,
  -39.7702,
  -39.7211,
  -39.6672,
  -39.6081,
  -39.5425,
  -39.4704,
  -39.3919,
  -39.3087,
  -31.7474,
  -31.7936,
  -31.839,
  -31.8837,
  -31.9276,
  -31.9711,
  -32.0145,
  -32.0583,
  -32.1024,
  -32.1468,
  -32.1904,
  -32.2351,
  -32.2801,
  -32.3252,
  -32.3704,
  -32.4156,
  -32.4601,
  -32.5043,
  -32.5481,
  -32.5918,
  -32.6356,
  -32.6796,
  -32.7243,
  -32.7697,
  -32.8162,
  -32.8628,
  -32.911,
  -32.9596,
  -33.008,
  -33.0558,
  -33.1028,
  -33.1489,
  -33.1943,
  -33.2392,
  -33.284,
  -33.3286,
  -33.373,
  -33.4171,
  -33.4609,
  -33.5045,
  -33.5472,
  -33.5907,
  -33.6341,
  -33.6772,
  -33.7199,
  -33.7625,
  -33.8049,
  -33.8475,
  -33.8904,
  -33.9338,
  -33.9778,
  -34.0226,
  -34.0683,
  -34.1147,
  -34.1622,
  -34.2107,
  -34.2592,
  -34.3095,
  -34.3601,
  -34.4109,
  -34.4618,
  -34.5128,
  -34.5644,
  -34.6169,
  -34.6707,
  -34.7261,
  -34.7829,
  -34.8409,
  -34.8997,
  -34.9585,
  -35.0171,
  -35.0748,
  -35.132,
  -35.1869,
  -35.2415,
  -35.2948,
  -35.347,
  -35.3986,
  -35.4499,
  -35.5014,
  -35.5525,
  -35.603,
  -35.6527,
  -35.7017,
  -35.7501,
  -35.798,
  -35.8454,
  -35.8923,
  -35.9387,
  -35.9849,
  -36.0297,
  -36.075,
  -36.1191,
  -36.1618,
  -36.2031,
  -36.2434,
  -36.2826,
  -36.321,
  -36.3585,
  -36.3949,
  -36.4302,
  -36.4642,
  -36.4969,
  -36.5278,
  -36.5568,
  -36.5837,
  -36.6091,
  -36.6337,
  -36.6581,
  -36.6815,
  -36.706,
  -36.7305,
  -36.7549,
  -36.7788,
  -36.8022,
  -36.8252,
  -36.848,
  -36.8705,
  -36.8928,
  -36.9147,
  -36.9363,
  -36.9578,
  -36.9793,
  -37.0011,
  -37.0236,
  -37.0469,
  -37.0707,
  -37.095,
  -37.1194,
  -37.143,
  -37.1682,
  -37.1939,
  -37.2201,
  -37.2467,
  -37.2734,
  -37.2997,
  -37.3258,
  -37.3512,
  -37.3763,
  -37.4013,
  -37.4268,
  -37.4533,
  -37.4807,
  -37.5091,
  -37.5381,
  -37.5672,
  -37.5962,
  -37.6248,
  -37.6529,
  -37.6805,
  -37.7065,
  -37.733,
  -37.759,
  -37.7847,
  -37.81,
  -37.8349,
  -37.8592,
  -37.8831,
  -37.9066,
  -37.9304,
  -37.955,
  -37.9809,
  -38.0081,
  -38.0369,
  -38.0669,
  -38.0973,
  -38.1271,
  -38.1556,
  -38.1825,
  -38.2082,
  -38.2335,
  -38.2591,
  -38.2853,
  -38.3121,
  -38.3385,
  -38.3662,
  -38.3941,
  -38.4224,
  -38.4508,
  -38.4789,
  -38.5066,
  -38.5337,
  -38.5602,
  -38.5864,
  -38.6126,
  -38.6389,
  -38.6649,
  -38.6906,
  -38.7155,
  -38.7395,
  -38.7623,
  -38.784,
  -38.8045,
  -38.824,
  -38.842,
  -38.8589,
  -38.8743,
  -38.8887,
  -38.9024,
  -38.9157,
  -38.9276,
  -38.9404,
  -38.9532,
  -38.9666,
  -38.9808,
  -38.996,
  -39.0123,
  -39.0292,
  -39.0463,
  -39.063,
  -39.0788,
  -39.0933,
  -39.1061,
  -39.1171,
  -39.1268,
  -39.1359,
  -39.1456,
  -39.1567,
  -39.1703,
  -39.1868,
  -39.2062,
  -39.2286,
  -39.2541,
  -39.2827,
  -39.3141,
  -39.3477,
  -39.3826,
  -39.418,
  -39.4536,
  -39.489,
  -39.523,
  -39.5574,
  -39.5908,
  -39.6229,
  -39.6536,
  -39.6828,
  -39.7109,
  -39.7381,
  -39.7646,
  -39.7902,
  -39.8146,
  -39.8378,
  -39.8599,
  -39.8811,
  -39.9016,
  -39.9211,
  -39.9394,
  -39.9563,
  -39.9717,
  -39.9859,
  -39.9993,
  -40.012,
  -40.024,
  -40.0357,
  -40.0469,
  -40.0581,
  -40.0692,
  -40.0801,
  -40.09,
  -40.0984,
  -40.1052,
  -40.1106,
  -40.1146,
  -40.1176,
  -40.1198,
  -40.1205,
  -40.1217,
  -40.1228,
  -40.1239,
  -40.1253,
  -40.1272,
  -40.1288,
  -40.1297,
  -40.1288,
  -40.1255,
  -40.1199,
  -40.112,
  -40.1018,
  -40.0895,
  -40.0758,
  -40.0615,
  -40.0473,
  -40.0334,
  -40.0191,
  -40.0031,
  -39.9841,
  -39.9616,
  -39.9358,
  -39.9071,
  -39.8757,
  -39.8413,
  -39.8036,
  -39.7622,
  -39.717,
  -39.6675,
  -39.6134,
  -39.5537,
  -39.4878,
  -39.4152,
  -39.3367,
  -39.2537,
  -31.663,
  -31.7097,
  -31.7557,
  -31.8007,
  -31.8449,
  -31.8885,
  -31.931,
  -31.9747,
  -32.0188,
  -32.0634,
  -32.1084,
  -32.1536,
  -32.199,
  -32.2446,
  -32.2902,
  -32.3355,
  -32.3804,
  -32.4247,
  -32.4685,
  -32.5122,
  -32.5549,
  -32.5989,
  -32.6434,
  -32.6888,
  -32.7353,
  -32.7828,
  -32.8311,
  -32.8797,
  -32.9281,
  -32.9759,
  -33.0228,
  -33.0689,
  -33.1145,
  -33.1596,
  -33.2045,
  -33.248,
  -33.2921,
  -33.3357,
  -33.3789,
  -33.4219,
  -33.4652,
  -33.5087,
  -33.5524,
  -33.5959,
  -33.6391,
  -33.6821,
  -33.7251,
  -33.7682,
  -33.8117,
  -33.8557,
  -33.9005,
  -33.945,
  -33.9914,
  -34.0386,
  -34.0868,
  -34.136,
  -34.1861,
  -34.2369,
  -34.2879,
  -34.339,
  -34.39,
  -34.4413,
  -34.4931,
  -34.5461,
  -34.6004,
  -34.6564,
  -34.714,
  -34.7718,
  -34.8311,
  -34.8905,
  -34.9493,
  -35.0073,
  -35.0641,
  -35.1196,
  -35.1736,
  -35.2265,
  -35.2784,
  -35.33,
  -35.3815,
  -35.4331,
  -35.4845,
  -35.5354,
  -35.5855,
  -35.6346,
  -35.6829,
  -35.7293,
  -35.776,
  -35.8221,
  -35.8679,
  -35.9136,
  -35.9594,
  -36.0049,
  -36.0496,
  -36.0931,
  -36.1352,
  -36.176,
  -36.2157,
  -36.2542,
  -36.2915,
  -36.3275,
  -36.3623,
  -36.3958,
  -36.4281,
  -36.4579,
  -36.4871,
  -36.5147,
  -36.5409,
  -36.5666,
  -36.5919,
  -36.6171,
  -36.6425,
  -36.6678,
  -36.6929,
  -36.7173,
  -36.7411,
  -36.7643,
  -36.787,
  -36.8094,
  -36.8316,
  -36.8537,
  -36.8757,
  -36.8978,
  -36.919,
  -36.9417,
  -36.9651,
  -36.9893,
  -37.0141,
  -37.0394,
  -37.0647,
  -37.0901,
  -37.1158,
  -37.142,
  -37.1686,
  -37.1954,
  -37.2222,
  -37.2485,
  -37.2743,
  -37.2994,
  -37.324,
  -37.3485,
  -37.3736,
  -37.3997,
  -37.4271,
  -37.4546,
  -37.4839,
  -37.5135,
  -37.5431,
  -37.5722,
  -37.6007,
  -37.6286,
  -37.6556,
  -37.6819,
  -37.7077,
  -37.7332,
  -37.7583,
  -37.7831,
  -37.8074,
  -37.8315,
  -37.8556,
  -37.8804,
  -37.9063,
  -37.9332,
  -37.9614,
  -37.9908,
  -38.021,
  -38.0513,
  -38.0798,
  -38.1081,
  -38.135,
  -38.1612,
  -38.1871,
  -38.2135,
  -38.2403,
  -38.2675,
  -38.2948,
  -38.322,
  -38.3493,
  -38.3768,
  -38.4045,
  -38.432,
  -38.4592,
  -38.4857,
  -38.5119,
  -38.5377,
  -38.5635,
  -38.5892,
  -38.6145,
  -38.6393,
  -38.6634,
  -38.6868,
  -38.7092,
  -38.7297,
  -38.7501,
  -38.7695,
  -38.7876,
  -38.8044,
  -38.82,
  -38.8344,
  -38.8479,
  -38.8607,
  -38.8732,
  -38.8855,
  -38.8982,
  -38.9115,
  -38.926,
  -38.9417,
  -38.9587,
  -38.9764,
  -38.9946,
  -39.0127,
  -39.0302,
  -39.0467,
  -39.0616,
  -39.0749,
  -39.0869,
  -39.0981,
  -39.1097,
  -39.1226,
  -39.1377,
  -39.1543,
  -39.1745,
  -39.1975,
  -39.2233,
  -39.2519,
  -39.2832,
  -39.3163,
  -39.3505,
  -39.3851,
  -39.4197,
  -39.4542,
  -39.4885,
  -39.5224,
  -39.5555,
  -39.5875,
  -39.6181,
  -39.6473,
  -39.6753,
  -39.7024,
  -39.7287,
  -39.7538,
  -39.7776,
  -39.8,
  -39.8213,
  -39.8417,
  -39.8616,
  -39.881,
  -39.8996,
  -39.9171,
  -39.9332,
  -39.9481,
  -39.962,
  -39.975,
  -39.9872,
  -39.9975,
  -40.0081,
  -40.0183,
  -40.0287,
  -40.0389,
  -40.0485,
  -40.057,
  -40.0641,
  -40.0696,
  -40.0736,
  -40.0764,
  -40.0781,
  -40.0791,
  -40.0798,
  -40.0805,
  -40.0814,
  -40.0829,
  -40.0848,
  -40.0866,
  -40.0874,
  -40.0863,
  -40.0827,
  -40.0766,
  -40.0682,
  -40.0576,
  -40.0452,
  -40.0312,
  -40.0167,
  -40.0021,
  -39.9876,
  -39.9726,
  -39.9557,
  -39.9358,
  -39.9124,
  -39.8856,
  -39.8559,
  -39.8234,
  -39.7881,
  -39.7496,
  -39.7076,
  -39.6618,
  -39.6117,
  -39.5569,
  -39.4956,
  -39.4291,
  -39.3563,
  -39.278,
  -39.1964,
  -31.5801,
  -31.6262,
  -31.6724,
  -31.7177,
  -31.762,
  -31.8056,
  -31.849,
  -31.8928,
  -31.9371,
  -31.982,
  -32.0274,
  -32.0731,
  -32.119,
  -32.1651,
  -32.211,
  -32.2556,
  -32.3005,
  -32.3449,
  -32.3887,
  -32.4323,
  -32.4759,
  -32.5197,
  -32.5643,
  -32.6097,
  -32.6563,
  -32.7038,
  -32.7521,
  -32.8006,
  -32.849,
  -32.8967,
  -32.9427,
  -32.989,
  -33.0349,
  -33.0806,
  -33.1258,
  -33.1704,
  -33.2143,
  -33.2574,
  -33.2999,
  -33.3423,
  -33.3852,
  -33.4286,
  -33.4726,
  -33.5167,
  -33.5606,
  -33.6042,
  -33.6467,
  -33.6904,
  -33.7344,
  -33.7789,
  -33.8242,
  -33.8703,
  -33.9174,
  -33.9653,
  -34.0143,
  -34.0644,
  -34.1152,
  -34.1666,
  -34.218,
  -34.2694,
  -34.3208,
  -34.3724,
  -34.4235,
  -34.4768,
  -34.5314,
  -34.5879,
  -34.6458,
  -34.705,
  -34.7647,
  -34.8243,
  -34.8833,
  -34.9412,
  -34.9978,
  -35.053,
  -35.1067,
  -35.1593,
  -35.2112,
  -35.2627,
  -35.3143,
  -35.365,
  -35.4166,
  -35.4678,
  -35.5182,
  -35.5676,
  -35.6158,
  -35.6628,
  -35.7088,
  -35.7541,
  -35.7993,
  -35.8447,
  -35.8903,
  -35.9359,
  -35.981,
  -36.0251,
  -36.068,
  -36.1094,
  -36.1494,
  -36.187,
  -36.224,
  -36.2597,
  -36.2941,
  -36.3272,
  -36.3593,
  -36.3902,
  -36.4198,
  -36.4482,
  -36.4755,
  -36.502,
  -36.5282,
  -36.5543,
  -36.5804,
  -36.6065,
  -36.6322,
  -36.6573,
  -36.6814,
  -36.7047,
  -36.7263,
  -36.7484,
  -36.7705,
  -36.7927,
  -36.8152,
  -36.838,
  -36.8612,
  -36.8849,
  -36.9092,
  -36.9343,
  -36.9601,
  -36.9862,
  -37.0123,
  -37.0384,
  -37.0647,
  -37.0912,
  -37.1181,
  -37.145,
  -37.1718,
  -37.1983,
  -37.2231,
  -37.2481,
  -37.2725,
  -37.2968,
  -37.3215,
  -37.3472,
  -37.3742,
  -37.4026,
  -37.4319,
  -37.4618,
  -37.4916,
  -37.521,
  -37.5496,
  -37.5774,
  -37.6043,
  -37.6305,
  -37.6561,
  -37.6814,
  -37.7064,
  -37.7309,
  -37.7554,
  -37.7798,
  -37.8039,
  -37.8298,
  -37.8569,
  -37.885,
  -37.9142,
  -37.9441,
  -37.9743,
  -38.0043,
  -38.0333,
  -38.0612,
  -38.0882,
  -38.1146,
  -38.1412,
  -38.1683,
  -38.1958,
  -38.2234,
  -38.2507,
  -38.2777,
  -38.3046,
  -38.3315,
  -38.3585,
  -38.3854,
  -38.4119,
  -38.4379,
  -38.4636,
  -38.488,
  -38.5134,
  -38.5385,
  -38.5633,
  -38.5874,
  -38.6109,
  -38.6338,
  -38.6559,
  -38.6773,
  -38.6977,
  -38.717,
  -38.7352,
  -38.7522,
  -38.768,
  -38.7826,
  -38.796,
  -38.8086,
  -38.8207,
  -38.8326,
  -38.8451,
  -38.8584,
  -38.8729,
  -38.8889,
  -38.9062,
  -38.9245,
  -38.9435,
  -38.9627,
  -38.9806,
  -38.9989,
  -39.016,
  -39.0316,
  -39.0457,
  -39.0591,
  -39.0727,
  -39.0873,
  -39.1039,
  -39.1226,
  -39.1437,
  -39.1672,
  -39.1933,
  -39.2222,
  -39.2533,
  -39.2861,
  -39.3197,
  -39.3534,
  -39.3871,
  -39.4206,
  -39.4541,
  -39.4874,
  -39.5201,
  -39.5519,
  -39.5823,
  -39.6114,
  -39.6393,
  -39.6663,
  -39.6924,
  -39.7173,
  -39.7407,
  -39.7616,
  -39.7824,
  -39.8023,
  -39.8218,
  -39.841,
  -39.8598,
  -39.8777,
  -39.8944,
  -39.9098,
  -39.9241,
  -39.9373,
  -39.9493,
  -39.96,
  -39.9698,
  -39.9791,
  -39.9884,
  -39.9979,
  -40.0071,
  -40.0157,
  -40.023,
  -40.0288,
  -40.033,
  -40.0356,
  -40.0369,
  -40.0373,
  -40.0375,
  -40.0377,
  -40.0385,
  -40.04,
  -40.042,
  -40.0439,
  -40.0446,
  -40.0433,
  -40.0393,
  -40.0327,
  -40.0237,
  -40.0128,
  -40,
  -39.9857,
  -39.9706,
  -39.9544,
  -39.9388,
  -39.9227,
  -39.9046,
  -39.8838,
  -39.8595,
  -39.8318,
  -39.8011,
  -39.7676,
  -39.7313,
  -39.6922,
  -39.6496,
  -39.6031,
  -39.5522,
  -39.4965,
  -39.4351,
  -39.3678,
  -39.2949,
  -39.2174,
  -39.1376,
  -31.4975,
  -31.5448,
  -31.5913,
  -31.6366,
  -31.6808,
  -31.7244,
  -31.7679,
  -31.8118,
  -31.8563,
  -31.9014,
  -31.9472,
  -31.9925,
  -32.039,
  -32.0856,
  -32.1318,
  -32.1774,
  -32.2223,
  -32.2665,
  -32.3102,
  -32.3536,
  -32.3971,
  -32.4411,
  -32.4858,
  -32.5314,
  -32.5781,
  -32.6247,
  -32.673,
  -32.7215,
  -32.7696,
  -32.8172,
  -32.864,
  -32.9105,
  -32.9569,
  -33.0031,
  -33.0488,
  -33.0936,
  -33.1375,
  -33.1803,
  -33.2226,
  -33.2647,
  -33.3074,
  -33.3499,
  -33.3941,
  -33.4386,
  -33.4831,
  -33.5275,
  -33.5717,
  -33.6159,
  -33.6604,
  -33.7054,
  -33.7511,
  -33.7977,
  -33.8453,
  -33.8941,
  -33.944,
  -33.9949,
  -34.0464,
  -34.0974,
  -34.1494,
  -34.2013,
  -34.2531,
  -34.3051,
  -34.3576,
  -34.4109,
  -34.4658,
  -34.5221,
  -34.58,
  -34.6393,
  -34.6989,
  -34.7586,
  -34.8178,
  -34.8757,
  -34.9323,
  -34.9861,
  -35.0396,
  -35.0921,
  -35.144,
  -35.1955,
  -35.2471,
  -35.2988,
  -35.3505,
  -35.4018,
  -35.4523,
  -35.502,
  -35.5502,
  -35.597,
  -35.6425,
  -35.6873,
  -35.7321,
  -35.7772,
  -35.8228,
  -35.8675,
  -35.9128,
  -35.9574,
  -36.0007,
  -36.0425,
  -36.0827,
  -36.1211,
  -36.158,
  -36.1933,
  -36.2275,
  -36.2607,
  -36.2928,
  -36.3241,
  -36.3544,
  -36.3837,
  -36.4119,
  -36.4392,
  -36.466,
  -36.4925,
  -36.5181,
  -36.5447,
  -36.5711,
  -36.5968,
  -36.6214,
  -36.6448,
  -36.6675,
  -36.6896,
  -36.7117,
  -36.7342,
  -36.7572,
  -36.7808,
  -36.805,
  -36.8297,
  -36.855,
  -36.8808,
  -36.9073,
  -36.934,
  -36.9607,
  -36.9875,
  -37.0132,
  -37.0401,
  -37.0672,
  -37.0942,
  -37.1212,
  -37.1475,
  -37.1734,
  -37.1986,
  -37.2232,
  -37.2475,
  -37.2721,
  -37.2974,
  -37.3239,
  -37.3519,
  -37.3811,
  -37.4109,
  -37.4408,
  -37.4701,
  -37.4985,
  -37.5261,
  -37.5528,
  -37.5779,
  -37.6034,
  -37.6288,
  -37.6537,
  -37.6783,
  -37.7029,
  -37.7278,
  -37.7537,
  -37.7807,
  -37.8089,
  -37.838,
  -37.8679,
  -37.8981,
  -37.9282,
  -37.9578,
  -37.9864,
  -38.0141,
  -38.041,
  -38.068,
  -38.0951,
  -38.1227,
  -38.1507,
  -38.1785,
  -38.2049,
  -38.2318,
  -38.2583,
  -38.2849,
  -38.3114,
  -38.3377,
  -38.3634,
  -38.3888,
  -38.414,
  -38.4389,
  -38.4638,
  -38.4885,
  -38.5127,
  -38.5362,
  -38.5593,
  -38.5818,
  -38.6038,
  -38.6251,
  -38.6455,
  -38.6649,
  -38.6832,
  -38.7004,
  -38.7165,
  -38.7313,
  -38.7449,
  -38.7574,
  -38.7693,
  -38.7801,
  -38.7923,
  -38.8055,
  -38.82,
  -38.8359,
  -38.8533,
  -38.8719,
  -38.8915,
  -38.9116,
  -38.9318,
  -38.9519,
  -38.971,
  -38.9887,
  -39.0051,
  -39.0206,
  -39.0362,
  -39.0526,
  -39.0705,
  -39.0905,
  -39.1125,
  -39.1367,
  -39.1633,
  -39.1925,
  -39.2235,
  -39.2559,
  -39.2888,
  -39.3217,
  -39.3544,
  -39.387,
  -39.4186,
  -39.4512,
  -39.4834,
  -39.5148,
  -39.5451,
  -39.574,
  -39.6017,
  -39.6285,
  -39.6544,
  -39.6792,
  -39.7025,
  -39.7244,
  -39.7449,
  -39.7646,
  -39.7838,
  -39.8028,
  -39.8216,
  -39.8398,
  -39.8569,
  -39.8727,
  -39.8872,
  -39.9002,
  -39.9116,
  -39.9217,
  -39.9307,
  -39.9391,
  -39.9477,
  -39.9565,
  -39.9653,
  -39.9737,
  -39.9812,
  -39.9872,
  -39.9914,
  -39.994,
  -39.995,
  -39.9949,
  -39.9944,
  -39.9933,
  -39.9938,
  -39.9951,
  -39.9971,
  -39.999,
  -39.9997,
  -39.9982,
  -39.994,
  -39.9871,
  -39.9777,
  -39.9662,
  -39.953,
  -39.9382,
  -39.9222,
  -39.9057,
  -39.8889,
  -39.8712,
  -39.852,
  -39.8302,
  -39.8051,
  -39.7766,
  -39.7452,
  -39.7109,
  -39.6738,
  -39.6341,
  -39.5908,
  -39.5435,
  -39.4916,
  -39.4347,
  -39.3721,
  -39.3037,
  -39.2306,
  -39.1543,
  -39.0772,
  -31.4165,
  -31.4642,
  -31.511,
  -31.5564,
  -31.6007,
  -31.6443,
  -31.6869,
  -31.7309,
  -31.7755,
  -31.8209,
  -31.8671,
  -31.9139,
  -31.9609,
  -32.0079,
  -32.0542,
  -32.0997,
  -32.1444,
  -32.1883,
  -32.2317,
  -32.2751,
  -32.3187,
  -32.362,
  -32.4071,
  -32.4531,
  -32.5,
  -32.5478,
  -32.596,
  -32.6444,
  -32.6924,
  -32.7398,
  -32.7867,
  -32.8331,
  -32.8797,
  -32.926,
  -32.972,
  -33.0169,
  -33.0599,
  -33.103,
  -33.1454,
  -33.1877,
  -33.2306,
  -33.2742,
  -33.3186,
  -33.3635,
  -33.4085,
  -33.4534,
  -33.4984,
  -33.5433,
  -33.5885,
  -33.6339,
  -33.6801,
  -33.7263,
  -33.7745,
  -33.824,
  -33.8747,
  -33.9263,
  -33.9785,
  -34.0311,
  -34.0837,
  -34.1362,
  -34.1886,
  -34.241,
  -34.2938,
  -34.3473,
  -34.4021,
  -34.4584,
  -34.5163,
  -34.5752,
  -34.6338,
  -34.6936,
  -34.7526,
  -34.8102,
  -34.8668,
  -34.9215,
  -34.975,
  -35.0273,
  -35.0791,
  -35.1306,
  -35.182,
  -35.2337,
  -35.2852,
  -35.3365,
  -35.3869,
  -35.4366,
  -35.4848,
  -35.5304,
  -35.5756,
  -35.6203,
  -35.6649,
  -35.7101,
  -35.7557,
  -35.8015,
  -35.847,
  -35.8917,
  -35.9353,
  -35.9774,
  -36.0176,
  -36.0558,
  -36.0925,
  -36.1276,
  -36.1617,
  -36.1949,
  -36.2276,
  -36.2595,
  -36.2895,
  -36.3196,
  -36.3485,
  -36.3764,
  -36.4037,
  -36.4305,
  -36.4572,
  -36.4842,
  -36.5111,
  -36.5373,
  -36.5625,
  -36.5865,
  -36.6096,
  -36.632,
  -36.6545,
  -36.6774,
  -36.701,
  -36.7254,
  -36.7504,
  -36.775,
  -36.8009,
  -36.8275,
  -36.8544,
  -36.8817,
  -36.9091,
  -36.9364,
  -36.9636,
  -36.9908,
  -37.018,
  -37.045,
  -37.0719,
  -37.0983,
  -37.1243,
  -37.1497,
  -37.1743,
  -37.1986,
  -37.223,
  -37.2481,
  -37.2745,
  -37.3022,
  -37.3302,
  -37.3599,
  -37.3896,
  -37.4188,
  -37.4471,
  -37.4745,
  -37.5011,
  -37.5271,
  -37.5527,
  -37.5781,
  -37.6031,
  -37.6279,
  -37.6529,
  -37.6784,
  -37.705,
  -37.7328,
  -37.7618,
  -37.7915,
  -37.8217,
  -37.852,
  -37.882,
  -37.9115,
  -37.94,
  -37.9667,
  -37.9938,
  -38.0208,
  -38.0482,
  -38.076,
  -38.104,
  -38.1319,
  -38.1592,
  -38.1859,
  -38.2122,
  -38.2383,
  -38.2642,
  -38.2898,
  -38.3151,
  -38.34,
  -38.3646,
  -38.3892,
  -38.4138,
  -38.438,
  -38.4618,
  -38.4853,
  -38.5081,
  -38.5303,
  -38.5519,
  -38.5733,
  -38.5927,
  -38.612,
  -38.6302,
  -38.6475,
  -38.6637,
  -38.6788,
  -38.6926,
  -38.7052,
  -38.7171,
  -38.7289,
  -38.7411,
  -38.7541,
  -38.7685,
  -38.7843,
  -38.8018,
  -38.8206,
  -38.8409,
  -38.8618,
  -38.8833,
  -38.9049,
  -38.9259,
  -38.9455,
  -38.964,
  -38.9816,
  -38.999,
  -39.0172,
  -39.0364,
  -39.0576,
  -39.0795,
  -39.1045,
  -39.1316,
  -39.161,
  -39.192,
  -39.2239,
  -39.2562,
  -39.2883,
  -39.3202,
  -39.3519,
  -39.3837,
  -39.4155,
  -39.4472,
  -39.4781,
  -39.5081,
  -39.5369,
  -39.5645,
  -39.5911,
  -39.6167,
  -39.6415,
  -39.6648,
  -39.6866,
  -39.7072,
  -39.7267,
  -39.7458,
  -39.7647,
  -39.7837,
  -39.8021,
  -39.8195,
  -39.8355,
  -39.8498,
  -39.8622,
  -39.8729,
  -39.8821,
  -39.8894,
  -39.8972,
  -39.9052,
  -39.9136,
  -39.9221,
  -39.9302,
  -39.9374,
  -39.9434,
  -39.9477,
  -39.9501,
  -39.9509,
  -39.9505,
  -39.9496,
  -39.9491,
  -39.9493,
  -39.9505,
  -39.9522,
  -39.9542,
  -39.9548,
  -39.9534,
  -39.9491,
  -39.9419,
  -39.9321,
  -39.9201,
  -39.906,
  -39.8902,
  -39.873,
  -39.8551,
  -39.8367,
  -39.8176,
  -39.7971,
  -39.7744,
  -39.7487,
  -39.7197,
  -39.6876,
  -39.6528,
  -39.6152,
  -39.5746,
  -39.5306,
  -39.4823,
  -39.4291,
  -39.3707,
  -39.3066,
  -39.2375,
  -39.1633,
  -39.0886,
  -39.0145,
  -31.3364,
  -31.3844,
  -31.4304,
  -31.476,
  -31.5206,
  -31.5645,
  -31.6082,
  -31.6522,
  -31.697,
  -31.7426,
  -31.7891,
  -31.8363,
  -31.8837,
  -31.9309,
  -31.9772,
  -32.0224,
  -32.0655,
  -32.109,
  -32.1523,
  -32.1957,
  -32.2398,
  -32.2846,
  -32.3303,
  -32.3768,
  -32.4241,
  -32.4719,
  -32.5201,
  -32.5682,
  -32.616,
  -32.6631,
  -32.7098,
  -32.7552,
  -32.8017,
  -32.8481,
  -32.894,
  -32.9391,
  -32.9833,
  -33.0268,
  -33.0697,
  -33.1127,
  -33.156,
  -33.2001,
  -33.2449,
  -33.2902,
  -33.3357,
  -33.3813,
  -33.4259,
  -33.4716,
  -33.5174,
  -33.5636,
  -33.6104,
  -33.6581,
  -33.7071,
  -33.7573,
  -33.8086,
  -33.8607,
  -33.9134,
  -33.9664,
  -34.0196,
  -34.0727,
  -34.1257,
  -34.1786,
  -34.2317,
  -34.2844,
  -34.3393,
  -34.3955,
  -34.4531,
  -34.5118,
  -34.5711,
  -34.6305,
  -34.6893,
  -34.7471,
  -34.8034,
  -34.8581,
  -34.9114,
  -34.9637,
  -35.0154,
  -35.0669,
  -35.1183,
  -35.1697,
  -35.2198,
  -35.2706,
  -35.3207,
  -35.3699,
  -35.4178,
  -35.4642,
  -35.5095,
  -35.5544,
  -35.5993,
  -35.6447,
  -35.6906,
  -35.7365,
  -35.7821,
  -35.8269,
  -35.8705,
  -35.9126,
  -35.9528,
  -35.9911,
  -36.0266,
  -36.0617,
  -36.0959,
  -36.1295,
  -36.1625,
  -36.195,
  -36.2267,
  -36.2574,
  -36.2868,
  -36.3151,
  -36.3424,
  -36.3693,
  -36.3962,
  -36.4233,
  -36.4506,
  -36.4775,
  -36.5034,
  -36.5282,
  -36.5521,
  -36.5743,
  -36.5974,
  -36.6209,
  -36.6453,
  -36.6706,
  -36.6964,
  -36.7227,
  -36.7493,
  -36.7762,
  -36.8035,
  -36.8311,
  -36.8589,
  -36.8867,
  -36.9143,
  -36.9418,
  -36.969,
  -36.996,
  -37.0227,
  -37.0492,
  -37.0752,
  -37.0998,
  -37.1247,
  -37.1492,
  -37.1737,
  -37.1987,
  -37.2249,
  -37.2525,
  -37.2813,
  -37.3108,
  -37.3403,
  -37.3694,
  -37.3976,
  -37.425,
  -37.4517,
  -37.4779,
  -37.5038,
  -37.5293,
  -37.5546,
  -37.5797,
  -37.6051,
  -37.6311,
  -37.6583,
  -37.6856,
  -37.715,
  -37.7449,
  -37.7751,
  -37.8052,
  -37.8351,
  -37.8644,
  -37.893,
  -37.9209,
  -37.9483,
  -37.9755,
  -38.0028,
  -38.0304,
  -38.0581,
  -38.0856,
  -38.1126,
  -38.139,
  -38.1649,
  -38.1904,
  -38.2158,
  -38.2408,
  -38.2655,
  -38.2899,
  -38.3141,
  -38.3374,
  -38.3617,
  -38.3858,
  -38.4095,
  -38.4327,
  -38.4554,
  -38.4775,
  -38.4992,
  -38.5202,
  -38.5403,
  -38.5595,
  -38.5777,
  -38.595,
  -38.6113,
  -38.6265,
  -38.6403,
  -38.6531,
  -38.6651,
  -38.6771,
  -38.6894,
  -38.7026,
  -38.717,
  -38.7328,
  -38.7502,
  -38.7695,
  -38.7901,
  -38.8119,
  -38.8349,
  -38.8569,
  -38.8795,
  -38.901,
  -38.9213,
  -38.9408,
  -38.96,
  -38.9796,
  -39.0003,
  -39.0225,
  -39.0465,
  -39.0721,
  -39.0998,
  -39.1294,
  -39.1603,
  -39.1919,
  -39.2236,
  -39.2552,
  -39.2864,
  -39.3175,
  -39.3486,
  -39.3797,
  -39.4107,
  -39.4411,
  -39.4706,
  -39.4991,
  -39.5265,
  -39.5529,
  -39.5784,
  -39.6029,
  -39.6263,
  -39.6483,
  -39.6679,
  -39.6875,
  -39.7065,
  -39.7255,
  -39.7445,
  -39.763,
  -39.7805,
  -39.7963,
  -39.8101,
  -39.8218,
  -39.8316,
  -39.8399,
  -39.8475,
  -39.855,
  -39.8628,
  -39.8711,
  -39.8793,
  -39.8872,
  -39.8943,
  -39.9001,
  -39.9043,
  -39.9066,
  -39.9072,
  -39.9065,
  -39.9054,
  -39.9045,
  -39.9043,
  -39.9051,
  -39.9066,
  -39.9085,
  -39.9091,
  -39.9077,
  -39.9033,
  -39.8958,
  -39.8856,
  -39.8728,
  -39.8577,
  -39.8406,
  -39.8221,
  -39.8026,
  -39.7816,
  -39.7611,
  -39.7395,
  -39.716,
  -39.6897,
  -39.6603,
  -39.6278,
  -39.5924,
  -39.5542,
  -39.513,
  -39.468,
  -39.4185,
  -39.3639,
  -39.3038,
  -39.2383,
  -39.1682,
  -39.0954,
  -39.0222,
  -38.9513,
  -31.2566,
  -31.3047,
  -31.3518,
  -31.3978,
  -31.4428,
  -31.487,
  -31.5309,
  -31.575,
  -31.6197,
  -31.6655,
  -31.7123,
  -31.7588,
  -31.8065,
  -31.8536,
  -31.8997,
  -31.9444,
  -31.9881,
  -32.0312,
  -32.0744,
  -32.118,
  -32.1627,
  -32.2083,
  -32.2547,
  -32.3018,
  -32.3495,
  -32.3971,
  -32.4441,
  -32.4919,
  -32.5393,
  -32.5861,
  -32.6326,
  -32.679,
  -32.7253,
  -32.7713,
  -32.8171,
  -32.8622,
  -32.9068,
  -32.9508,
  -32.9945,
  -33.0382,
  -33.0824,
  -33.1262,
  -33.1715,
  -33.2175,
  -33.2636,
  -33.3098,
  -33.3561,
  -33.4025,
  -33.4491,
  -33.4961,
  -33.5438,
  -33.5924,
  -33.6419,
  -33.6927,
  -33.7445,
  -33.797,
  -33.8499,
  -33.9023,
  -33.9559,
  -34.0094,
  -34.063,
  -34.1164,
  -34.17,
  -34.2239,
  -34.2788,
  -34.335,
  -34.3924,
  -34.4506,
  -34.5095,
  -34.5685,
  -34.6271,
  -34.6848,
  -34.7411,
  -34.7957,
  -34.8479,
  -34.9002,
  -34.952,
  -35.0035,
  -35.0548,
  -35.1058,
  -35.1564,
  -35.2063,
  -35.2555,
  -35.3037,
  -35.3513,
  -35.3976,
  -35.443,
  -35.4882,
  -35.5337,
  -35.5795,
  -35.6257,
  -35.6717,
  -35.7164,
  -35.7612,
  -35.8048,
  -35.847,
  -35.8872,
  -35.9258,
  -35.9625,
  -35.9978,
  -36.0321,
  -36.066,
  -36.0994,
  -36.1323,
  -36.1644,
  -36.1954,
  -36.2251,
  -36.2535,
  -36.2809,
  -36.3077,
  -36.3337,
  -36.361,
  -36.3886,
  -36.4163,
  -36.4431,
  -36.469,
  -36.4939,
  -36.5181,
  -36.5423,
  -36.5666,
  -36.5918,
  -36.6179,
  -36.6446,
  -36.6715,
  -36.6987,
  -36.726,
  -36.7534,
  -36.7812,
  -36.8092,
  -36.8374,
  -36.8644,
  -36.8921,
  -36.9193,
  -36.9463,
  -36.9728,
  -36.9992,
  -37.0254,
  -37.0512,
  -37.0765,
  -37.1014,
  -37.1261,
  -37.1513,
  -37.1775,
  -37.2049,
  -37.2335,
  -37.2628,
  -37.2921,
  -37.3211,
  -37.3494,
  -37.3772,
  -37.4042,
  -37.4309,
  -37.456,
  -37.4818,
  -37.5076,
  -37.5331,
  -37.5587,
  -37.5854,
  -37.6129,
  -37.6415,
  -37.6709,
  -37.7007,
  -37.7306,
  -37.7603,
  -37.7899,
  -37.8192,
  -37.848,
  -37.8762,
  -37.904,
  -37.9312,
  -37.9585,
  -37.9855,
  -38.0123,
  -38.039,
  -38.0654,
  -38.0902,
  -38.1155,
  -38.1405,
  -38.1651,
  -38.1894,
  -38.2135,
  -38.2374,
  -38.2613,
  -38.2853,
  -38.3093,
  -38.3333,
  -38.3571,
  -38.3804,
  -38.4031,
  -38.4252,
  -38.4466,
  -38.4674,
  -38.4873,
  -38.5063,
  -38.5244,
  -38.5416,
  -38.5579,
  -38.573,
  -38.5869,
  -38.5998,
  -38.6121,
  -38.6233,
  -38.6359,
  -38.6494,
  -38.664,
  -38.68,
  -38.6976,
  -38.7172,
  -38.7384,
  -38.7612,
  -38.7854,
  -38.8098,
  -38.8337,
  -38.8569,
  -38.879,
  -38.9001,
  -38.9209,
  -38.9419,
  -38.9639,
  -38.9871,
  -39.0118,
  -39.0382,
  -39.0666,
  -39.0964,
  -39.1273,
  -39.1586,
  -39.19,
  -39.2213,
  -39.2523,
  -39.283,
  -39.3136,
  -39.3431,
  -39.3733,
  -39.4031,
  -39.4321,
  -39.4601,
  -39.4872,
  -39.5132,
  -39.5384,
  -39.5626,
  -39.5858,
  -39.6079,
  -39.6286,
  -39.6484,
  -39.6676,
  -39.6866,
  -39.7054,
  -39.724,
  -39.7414,
  -39.7569,
  -39.7701,
  -39.7808,
  -39.7896,
  -39.7972,
  -39.8042,
  -39.8115,
  -39.8193,
  -39.8276,
  -39.8358,
  -39.8436,
  -39.8506,
  -39.8563,
  -39.8603,
  -39.8626,
  -39.8631,
  -39.8623,
  -39.8609,
  -39.8596,
  -39.8581,
  -39.8585,
  -39.8598,
  -39.8611,
  -39.8614,
  -39.86,
  -39.8555,
  -39.8478,
  -39.8369,
  -39.8232,
  -39.8069,
  -39.7885,
  -39.7684,
  -39.7473,
  -39.7259,
  -39.704,
  -39.6815,
  -39.6573,
  -39.6307,
  -39.601,
  -39.5682,
  -39.5323,
  -39.4934,
  -39.4512,
  -39.405,
  -39.3541,
  -39.2979,
  -39.2361,
  -39.1693,
  -39.0986,
  -39.0262,
  -38.9547,
  -38.8869,
  -31.1797,
  -31.2277,
  -31.2749,
  -31.321,
  -31.3663,
  -31.4108,
  -31.4549,
  -31.4981,
  -31.5429,
  -31.5889,
  -31.636,
  -31.6837,
  -31.7314,
  -31.7783,
  -31.824,
  -31.8684,
  -31.9118,
  -31.9548,
  -31.9981,
  -32.042,
  -32.0872,
  -32.1325,
  -32.1795,
  -32.2271,
  -32.2747,
  -32.3223,
  -32.37,
  -32.4174,
  -32.4645,
  -32.5111,
  -32.5574,
  -32.6034,
  -32.6494,
  -32.6953,
  -32.7409,
  -32.786,
  -32.8299,
  -32.8744,
  -32.9189,
  -32.9635,
  -33.0085,
  -33.0541,
  -33.1004,
  -33.1471,
  -33.1939,
  -33.2408,
  -33.2877,
  -33.3349,
  -33.3824,
  -33.4305,
  -33.4791,
  -33.5285,
  -33.5778,
  -33.6291,
  -33.6813,
  -33.7341,
  -33.7874,
  -33.841,
  -33.8948,
  -33.9487,
  -34.0026,
  -34.0565,
  -34.1104,
  -34.1647,
  -34.2198,
  -34.2759,
  -34.3329,
  -34.3907,
  -34.4491,
  -34.5067,
  -34.5649,
  -34.6223,
  -34.6784,
  -34.733,
  -34.7863,
  -34.8387,
  -34.8906,
  -34.9422,
  -34.9934,
  -35.0442,
  -35.0941,
  -35.1431,
  -35.1912,
  -35.2385,
  -35.285,
  -35.3309,
  -35.3755,
  -35.421,
  -35.4668,
  -35.5129,
  -35.5593,
  -35.6055,
  -35.6511,
  -35.696,
  -35.7399,
  -35.7823,
  -35.823,
  -35.862,
  -35.8991,
  -35.9348,
  -35.9695,
  -36.0036,
  -36.0372,
  -36.0702,
  -36.1013,
  -36.1324,
  -36.162,
  -36.1904,
  -36.2177,
  -36.2447,
  -36.2719,
  -36.2996,
  -36.3278,
  -36.3561,
  -36.3839,
  -36.4108,
  -36.4368,
  -36.4622,
  -36.4875,
  -36.513,
  -36.5392,
  -36.566,
  -36.5935,
  -36.6212,
  -36.6478,
  -36.6754,
  -36.703,
  -36.7309,
  -36.7591,
  -36.7874,
  -36.8157,
  -36.8435,
  -36.8708,
  -36.8977,
  -36.9242,
  -36.9506,
  -36.9771,
  -37.0032,
  -37.0289,
  -37.0541,
  -37.0794,
  -37.1049,
  -37.1311,
  -37.1585,
  -37.1869,
  -37.2148,
  -37.244,
  -37.273,
  -37.3017,
  -37.33,
  -37.3575,
  -37.3849,
  -37.4113,
  -37.4374,
  -37.4633,
  -37.4894,
  -37.5157,
  -37.5425,
  -37.5704,
  -37.599,
  -37.6282,
  -37.6578,
  -37.6873,
  -37.7168,
  -37.7461,
  -37.7754,
  -37.8044,
  -37.8319,
  -37.8599,
  -37.887,
  -37.9138,
  -37.9397,
  -37.9658,
  -37.9913,
  -38.0168,
  -38.0418,
  -38.0664,
  -38.0905,
  -38.1142,
  -38.1377,
  -38.1612,
  -38.1846,
  -38.2082,
  -38.232,
  -38.2559,
  -38.28,
  -38.304,
  -38.3275,
  -38.3503,
  -38.3724,
  -38.3936,
  -38.414,
  -38.4336,
  -38.4514,
  -38.4693,
  -38.4864,
  -38.5025,
  -38.5176,
  -38.5316,
  -38.5446,
  -38.5571,
  -38.5697,
  -38.5827,
  -38.5966,
  -38.6117,
  -38.6281,
  -38.6462,
  -38.6661,
  -38.6882,
  -38.7121,
  -38.7373,
  -38.763,
  -38.7884,
  -38.813,
  -38.8363,
  -38.8586,
  -38.8806,
  -38.9028,
  -38.9257,
  -38.9498,
  -38.9754,
  -39.0016,
  -39.0305,
  -39.0606,
  -39.0916,
  -39.123,
  -39.1543,
  -39.1856,
  -39.2167,
  -39.2474,
  -39.2778,
  -39.3079,
  -39.3374,
  -39.3664,
  -39.3947,
  -39.4221,
  -39.4487,
  -39.4743,
  -39.4991,
  -39.5228,
  -39.5457,
  -39.5676,
  -39.5883,
  -39.6083,
  -39.6278,
  -39.6471,
  -39.666,
  -39.6842,
  -39.7014,
  -39.7163,
  -39.7288,
  -39.7387,
  -39.7466,
  -39.7534,
  -39.7599,
  -39.7659,
  -39.7738,
  -39.782,
  -39.7904,
  -39.7983,
  -39.8051,
  -39.8107,
  -39.8148,
  -39.8171,
  -39.8177,
  -39.8168,
  -39.8153,
  -39.8138,
  -39.813,
  -39.8131,
  -39.8138,
  -39.8147,
  -39.8146,
  -39.8127,
  -39.8077,
  -39.7994,
  -39.7877,
  -39.7729,
  -39.7555,
  -39.7358,
  -39.7144,
  -39.6919,
  -39.6692,
  -39.6463,
  -39.6228,
  -39.598,
  -39.5711,
  -39.5412,
  -39.5082,
  -39.4718,
  -39.4321,
  -39.3886,
  -39.3409,
  -39.2882,
  -39.2301,
  -39.1667,
  -39.0986,
  -39.0274,
  -38.9555,
  -38.8849,
  -38.8206,
  -31.1047,
  -31.1526,
  -31.1987,
  -31.2449,
  -31.2902,
  -31.3349,
  -31.3791,
  -31.4234,
  -31.4685,
  -31.5147,
  -31.5619,
  -31.6098,
  -31.6574,
  -31.7042,
  -31.7496,
  -31.7939,
  -31.8363,
  -31.8794,
  -31.9229,
  -31.9673,
  -32.0128,
  -32.0596,
  -32.107,
  -32.1548,
  -32.2024,
  -32.2498,
  -32.2971,
  -32.3441,
  -32.3909,
  -32.4373,
  -32.4833,
  -32.5283,
  -32.574,
  -32.6196,
  -32.665,
  -32.7103,
  -32.7555,
  -32.8006,
  -32.8458,
  -32.8912,
  -32.937,
  -32.9835,
  -33.0306,
  -33.0781,
  -33.1257,
  -33.1732,
  -33.2209,
  -33.268,
  -33.3165,
  -33.3656,
  -33.4152,
  -33.4654,
  -33.5165,
  -33.5683,
  -33.6209,
  -33.6741,
  -33.7277,
  -33.7815,
  -33.8355,
  -33.8896,
  -33.9437,
  -33.9979,
  -34.0522,
  -34.1058,
  -34.161,
  -34.2169,
  -34.2737,
  -34.331,
  -34.3889,
  -34.4469,
  -34.5046,
  -34.5615,
  -34.6173,
  -34.6719,
  -34.7254,
  -34.778,
  -34.8301,
  -34.8818,
  -34.9331,
  -34.9836,
  -35.0321,
  -35.0804,
  -35.1275,
  -35.1734,
  -35.2188,
  -35.264,
  -35.3092,
  -35.3548,
  -35.4008,
  -35.4472,
  -35.4936,
  -35.5398,
  -35.5855,
  -35.6305,
  -35.6746,
  -35.7174,
  -35.7587,
  -35.7983,
  -35.8351,
  -35.8714,
  -35.9067,
  -35.9411,
  -35.9748,
  -36.0078,
  -36.0398,
  -36.0706,
  -36.1,
  -36.1284,
  -36.1557,
  -36.1831,
  -36.2107,
  -36.239,
  -36.2679,
  -36.2968,
  -36.3254,
  -36.3531,
  -36.3801,
  -36.4057,
  -36.4321,
  -36.4588,
  -36.4859,
  -36.5137,
  -36.5419,
  -36.5703,
  -36.5986,
  -36.6266,
  -36.6544,
  -36.6824,
  -36.7105,
  -36.7389,
  -36.7672,
  -36.7951,
  -36.8223,
  -36.8493,
  -36.8759,
  -36.9026,
  -36.9294,
  -36.956,
  -36.9812,
  -37.007,
  -37.0327,
  -37.0586,
  -37.085,
  -37.1122,
  -37.1403,
  -37.1691,
  -37.1982,
  -37.2273,
  -37.2564,
  -37.2849,
  -37.3131,
  -37.3408,
  -37.3678,
  -37.3944,
  -37.4207,
  -37.4472,
  -37.4739,
  -37.5013,
  -37.5293,
  -37.5579,
  -37.5859,
  -37.6151,
  -37.6443,
  -37.6735,
  -37.7028,
  -37.7321,
  -37.7613,
  -37.7899,
  -37.8174,
  -37.8439,
  -37.8698,
  -37.8951,
  -37.9199,
  -37.9445,
  -37.9689,
  -37.9931,
  -38.0167,
  -38.0398,
  -38.0627,
  -38.0853,
  -38.1081,
  -38.1311,
  -38.1543,
  -38.178,
  -38.2008,
  -38.225,
  -38.2491,
  -38.2731,
  -38.2958,
  -38.3178,
  -38.3389,
  -38.3589,
  -38.3781,
  -38.3966,
  -38.4145,
  -38.4314,
  -38.4476,
  -38.4626,
  -38.4766,
  -38.4899,
  -38.5028,
  -38.5158,
  -38.5293,
  -38.5437,
  -38.5592,
  -38.5761,
  -38.5949,
  -38.6157,
  -38.6386,
  -38.6636,
  -38.69,
  -38.717,
  -38.7426,
  -38.7682,
  -38.7925,
  -38.8157,
  -38.8385,
  -38.8616,
  -38.8855,
  -38.9103,
  -38.9366,
  -38.9644,
  -38.9938,
  -39.0244,
  -39.0556,
  -39.0873,
  -39.119,
  -39.1505,
  -39.1818,
  -39.2127,
  -39.2431,
  -39.2727,
  -39.3017,
  -39.33,
  -39.3576,
  -39.3844,
  -39.4104,
  -39.4354,
  -39.4597,
  -39.4828,
  -39.505,
  -39.5265,
  -39.5472,
  -39.5665,
  -39.5864,
  -39.6057,
  -39.6248,
  -39.643,
  -39.6596,
  -39.6741,
  -39.6858,
  -39.6948,
  -39.702,
  -39.708,
  -39.7141,
  -39.7206,
  -39.7283,
  -39.7367,
  -39.7453,
  -39.7533,
  -39.7603,
  -39.7658,
  -39.7698,
  -39.7722,
  -39.7729,
  -39.7721,
  -39.7706,
  -39.769,
  -39.768,
  -39.7678,
  -39.7681,
  -39.7683,
  -39.7674,
  -39.7646,
  -39.7589,
  -39.7497,
  -39.7371,
  -39.7214,
  -39.7028,
  -39.6821,
  -39.6597,
  -39.6364,
  -39.6127,
  -39.5876,
  -39.5631,
  -39.5377,
  -39.5103,
  -39.4803,
  -39.4469,
  -39.41,
  -39.3694,
  -39.3245,
  -39.275,
  -39.2202,
  -39.1603,
  -39.0952,
  -39.026,
  -38.9545,
  -38.8835,
  -38.8159,
  -38.755,
  -31.0304,
  -31.0784,
  -31.1254,
  -31.1714,
  -31.2167,
  -31.2613,
  -31.3056,
  -31.3501,
  -31.3955,
  -31.442,
  -31.4894,
  -31.5373,
  -31.5839,
  -31.6304,
  -31.6758,
  -31.7201,
  -31.7637,
  -31.8073,
  -31.8513,
  -31.8961,
  -31.9421,
  -31.9892,
  -32.0368,
  -32.0846,
  -32.1321,
  -32.1793,
  -32.2251,
  -32.2716,
  -32.318,
  -32.3642,
  -32.4101,
  -32.4558,
  -32.5015,
  -32.5469,
  -32.5925,
  -32.6379,
  -32.6836,
  -32.7291,
  -32.7749,
  -32.8209,
  -32.8674,
  -32.9148,
  -32.9617,
  -33.01,
  -33.0583,
  -33.1066,
  -33.155,
  -33.2039,
  -33.2534,
  -33.3036,
  -33.3542,
  -33.4053,
  -33.457,
  -33.5093,
  -33.5623,
  -33.6159,
  -33.6698,
  -33.724,
  -33.7772,
  -33.8313,
  -33.8855,
  -33.9399,
  -33.9945,
  -34.0493,
  -34.1046,
  -34.1604,
  -34.2169,
  -34.2738,
  -34.3309,
  -34.3881,
  -34.445,
  -34.5013,
  -34.5568,
  -34.6113,
  -34.665,
  -34.7169,
  -34.7692,
  -34.8211,
  -34.8724,
  -34.9231,
  -34.9726,
  -35.0204,
  -35.0666,
  -35.1112,
  -35.1554,
  -35.1995,
  -35.244,
  -35.2893,
  -35.3353,
  -35.3819,
  -35.4282,
  -35.4743,
  -35.5187,
  -35.5637,
  -35.6079,
  -35.6511,
  -35.693,
  -35.7334,
  -35.7721,
  -35.8093,
  -35.8453,
  -35.8801,
  -35.914,
  -35.947,
  -35.9788,
  -36.0095,
  -36.0389,
  -36.0673,
  -36.095,
  -36.1228,
  -36.151,
  -36.179,
  -36.2085,
  -36.238,
  -36.267,
  -36.2954,
  -36.3233,
  -36.3509,
  -36.3785,
  -36.4062,
  -36.4342,
  -36.4626,
  -36.4915,
  -36.5207,
  -36.5497,
  -36.5783,
  -36.6065,
  -36.6344,
  -36.6625,
  -36.6907,
  -36.7188,
  -36.7456,
  -36.773,
  -36.7999,
  -36.827,
  -36.8543,
  -36.8815,
  -36.9085,
  -36.9352,
  -36.9616,
  -36.9879,
  -37.014,
  -37.0406,
  -37.0679,
  -37.0957,
  -37.1244,
  -37.1535,
  -37.1827,
  -37.212,
  -37.241,
  -37.2696,
  -37.2978,
  -37.3252,
  -37.3512,
  -37.378,
  -37.4049,
  -37.4321,
  -37.4598,
  -37.4879,
  -37.5165,
  -37.5453,
  -37.5741,
  -37.6031,
  -37.6323,
  -37.6616,
  -37.6909,
  -37.7199,
  -37.748,
  -37.7751,
  -37.8009,
  -37.8258,
  -37.85,
  -37.8739,
  -37.8976,
  -37.9211,
  -37.9443,
  -37.9661,
  -37.9883,
  -38.0102,
  -38.032,
  -38.0541,
  -38.0765,
  -38.0995,
  -38.1228,
  -38.1466,
  -38.1706,
  -38.1949,
  -38.2187,
  -38.2418,
  -38.2637,
  -38.2844,
  -38.3042,
  -38.3231,
  -38.3413,
  -38.3591,
  -38.376,
  -38.3922,
  -38.4074,
  -38.4217,
  -38.4353,
  -38.4488,
  -38.4623,
  -38.4753,
  -38.4901,
  -38.5061,
  -38.5236,
  -38.543,
  -38.5648,
  -38.5889,
  -38.6151,
  -38.6429,
  -38.671,
  -38.6984,
  -38.7248,
  -38.7498,
  -38.7737,
  -38.7971,
  -38.8208,
  -38.8454,
  -38.8712,
  -38.8979,
  -38.9262,
  -38.9562,
  -38.9873,
  -39.019,
  -39.051,
  -39.083,
  -39.1148,
  -39.1465,
  -39.1778,
  -39.2081,
  -39.2375,
  -39.2661,
  -39.2928,
  -39.3198,
  -39.346,
  -39.3713,
  -39.3957,
  -39.419,
  -39.4412,
  -39.4629,
  -39.4839,
  -39.5046,
  -39.525,
  -39.5452,
  -39.5648,
  -39.584,
  -39.602,
  -39.6183,
  -39.6321,
  -39.6432,
  -39.6516,
  -39.6578,
  -39.6632,
  -39.6687,
  -39.6749,
  -39.6825,
  -39.691,
  -39.6998,
  -39.7081,
  -39.7151,
  -39.7207,
  -39.7246,
  -39.7269,
  -39.7276,
  -39.7269,
  -39.7255,
  -39.724,
  -39.723,
  -39.7217,
  -39.7215,
  -39.7208,
  -39.7189,
  -39.7148,
  -39.708,
  -39.6979,
  -39.6843,
  -39.6676,
  -39.6484,
  -39.627,
  -39.6044,
  -39.5802,
  -39.5556,
  -39.5306,
  -39.505,
  -39.4786,
  -39.4506,
  -39.4202,
  -39.3865,
  -39.3492,
  -39.3074,
  -39.2611,
  -39.2097,
  -39.153,
  -39.091,
  -39.0246,
  -38.9546,
  -38.8833,
  -38.8131,
  -38.7477,
  -38.6909,
  -30.9584,
  -31.0063,
  -31.0533,
  -31.0993,
  -31.1444,
  -31.189,
  -31.2336,
  -31.2774,
  -31.3231,
  -31.3699,
  -31.4176,
  -31.4655,
  -31.513,
  -31.5595,
  -31.6049,
  -31.6493,
  -31.6933,
  -31.7374,
  -31.7821,
  -31.8276,
  -31.8741,
  -31.9214,
  -31.9681,
  -32.0158,
  -32.0631,
  -32.1099,
  -32.1563,
  -32.2024,
  -32.2484,
  -32.2943,
  -32.34,
  -32.3854,
  -32.4309,
  -32.4766,
  -32.5223,
  -32.5681,
  -32.6141,
  -32.6591,
  -32.7053,
  -32.7519,
  -32.7991,
  -32.8472,
  -32.896,
  -32.9451,
  -32.9943,
  -33.0434,
  -33.0928,
  -33.1425,
  -33.1929,
  -33.2439,
  -33.2955,
  -33.3473,
  -33.3996,
  -33.4514,
  -33.5047,
  -33.5586,
  -33.6128,
  -33.667,
  -33.7212,
  -33.7754,
  -33.8298,
  -33.8844,
  -33.9393,
  -33.9944,
  -34.0498,
  -34.1056,
  -34.1618,
  -34.2182,
  -34.2745,
  -34.3298,
  -34.3857,
  -34.4411,
  -34.496,
  -34.5504,
  -34.6041,
  -34.6572,
  -34.7097,
  -34.7618,
  -34.8133,
  -34.8642,
  -34.9138,
  -34.9614,
  -35.0069,
  -35.0508,
  -35.0938,
  -35.1369,
  -35.1797,
  -35.2245,
  -35.2704,
  -35.3167,
  -35.3629,
  -35.4087,
  -35.4538,
  -35.4985,
  -35.5426,
  -35.5861,
  -35.6284,
  -35.6694,
  -35.709,
  -35.7471,
  -35.7838,
  -35.8192,
  -35.8535,
  -35.8867,
  -35.9187,
  -35.9485,
  -35.9782,
  -36.0069,
  -36.0351,
  -36.0634,
  -36.0922,
  -36.1218,
  -36.1517,
  -36.1816,
  -36.211,
  -36.2399,
  -36.2684,
  -36.2969,
  -36.3255,
  -36.3541,
  -36.3829,
  -36.4121,
  -36.4418,
  -36.4715,
  -36.5001,
  -36.5293,
  -36.5578,
  -36.5858,
  -36.6137,
  -36.6415,
  -36.6693,
  -36.697,
  -36.7244,
  -36.7517,
  -36.7793,
  -36.8072,
  -36.835,
  -36.8626,
  -36.8899,
  -36.9168,
  -36.9435,
  -36.9702,
  -36.9971,
  -37.0242,
  -37.052,
  -37.0794,
  -37.1084,
  -37.1376,
  -37.1669,
  -37.1961,
  -37.2251,
  -37.2536,
  -37.2816,
  -37.3092,
  -37.3366,
  -37.364,
  -37.3916,
  -37.4195,
  -37.4477,
  -37.4761,
  -37.5047,
  -37.5334,
  -37.5621,
  -37.5912,
  -37.6204,
  -37.6496,
  -37.6781,
  -37.7057,
  -37.731,
  -37.756,
  -37.78,
  -37.8034,
  -37.8264,
  -37.8494,
  -37.8722,
  -37.8948,
  -37.9169,
  -37.9384,
  -37.9595,
  -37.9806,
  -38.0019,
  -38.0235,
  -38.0459,
  -38.0689,
  -38.0923,
  -38.1162,
  -38.1401,
  -38.1638,
  -38.1868,
  -38.2085,
  -38.2292,
  -38.2488,
  -38.2675,
  -38.2857,
  -38.3024,
  -38.3195,
  -38.3358,
  -38.3512,
  -38.366,
  -38.3802,
  -38.3943,
  -38.4084,
  -38.423,
  -38.4383,
  -38.4547,
  -38.4726,
  -38.4927,
  -38.5153,
  -38.5407,
  -38.5681,
  -38.5969,
  -38.6259,
  -38.6545,
  -38.6818,
  -38.7076,
  -38.7323,
  -38.7565,
  -38.7808,
  -38.806,
  -38.8321,
  -38.8594,
  -38.8882,
  -38.9175,
  -38.9491,
  -38.9812,
  -39.0135,
  -39.0459,
  -39.0781,
  -39.11,
  -39.1415,
  -39.1719,
  -39.201,
  -39.2292,
  -39.2564,
  -39.2827,
  -39.3082,
  -39.3326,
  -39.3559,
  -39.3784,
  -39.3998,
  -39.4208,
  -39.4416,
  -39.4622,
  -39.4828,
  -39.5033,
  -39.5233,
  -39.5425,
  -39.5603,
  -39.5762,
  -39.5894,
  -39.5999,
  -39.6077,
  -39.6134,
  -39.6182,
  -39.6232,
  -39.6292,
  -39.6357,
  -39.6443,
  -39.6532,
  -39.6616,
  -39.6688,
  -39.6743,
  -39.6782,
  -39.6804,
  -39.6811,
  -39.6805,
  -39.6791,
  -39.6776,
  -39.6767,
  -39.6762,
  -39.6755,
  -39.6739,
  -39.6706,
  -39.6652,
  -39.6572,
  -39.646,
  -39.6317,
  -39.6145,
  -39.595,
  -39.5736,
  -39.5506,
  -39.5263,
  -39.5009,
  -39.4747,
  -39.4477,
  -39.42,
  -39.3909,
  -39.3598,
  -39.3257,
  -39.2877,
  -39.2449,
  -39.1973,
  -39.1443,
  -39.0859,
  -39.0225,
  -38.9548,
  -38.8846,
  -38.8137,
  -38.7455,
  -38.6831,
  -38.6308,
  -30.8874,
  -30.9355,
  -30.9825,
  -31.0275,
  -31.0726,
  -31.1173,
  -31.162,
  -31.2073,
  -31.2534,
  -31.3005,
  -31.3484,
  -31.3963,
  -31.4439,
  -31.4904,
  -31.5358,
  -31.5804,
  -31.6249,
  -31.6688,
  -31.7143,
  -31.7606,
  -31.8076,
  -31.8551,
  -31.9029,
  -31.9505,
  -31.9976,
  -32.0441,
  -32.09,
  -32.1356,
  -32.1812,
  -32.2267,
  -32.2721,
  -32.3175,
  -32.362,
  -32.4078,
  -32.4539,
  -32.5001,
  -32.5464,
  -32.5928,
  -32.6394,
  -32.6864,
  -32.7342,
  -32.7829,
  -32.8326,
  -32.8826,
  -32.9328,
  -32.9829,
  -33.0332,
  -33.0829,
  -33.1341,
  -33.186,
  -33.2382,
  -33.2907,
  -33.3434,
  -33.3964,
  -33.4499,
  -33.504,
  -33.5583,
  -33.6125,
  -33.6667,
  -33.721,
  -33.7755,
  -33.8304,
  -33.8857,
  -33.9411,
  -33.9957,
  -34.0517,
  -34.1077,
  -34.1634,
  -34.219,
  -34.2741,
  -34.3289,
  -34.3834,
  -34.4374,
  -34.4913,
  -34.5449,
  -34.598,
  -34.6506,
  -34.7027,
  -34.7543,
  -34.8053,
  -34.8552,
  -34.9019,
  -34.9473,
  -34.9907,
  -35.0332,
  -35.0756,
  -35.1188,
  -35.1633,
  -35.2089,
  -35.2547,
  -35.3005,
  -35.3457,
  -35.39,
  -35.4342,
  -35.4781,
  -35.5215,
  -35.5641,
  -35.6055,
  -35.6458,
  -35.6837,
  -35.7212,
  -35.7573,
  -35.7921,
  -35.8256,
  -35.8581,
  -35.8894,
  -35.9196,
  -35.9489,
  -35.9777,
  -36.0066,
  -36.0361,
  -36.0662,
  -36.0967,
  -36.1267,
  -36.1563,
  -36.1854,
  -36.2144,
  -36.2435,
  -36.2719,
  -36.3013,
  -36.3308,
  -36.3604,
  -36.3907,
  -36.4212,
  -36.4515,
  -36.481,
  -36.5099,
  -36.538,
  -36.5656,
  -36.5931,
  -36.6206,
  -36.6481,
  -36.6757,
  -36.7035,
  -36.7318,
  -36.7602,
  -36.7887,
  -36.8169,
  -36.8436,
  -36.8711,
  -36.8983,
  -36.9254,
  -36.9527,
  -36.98,
  -37.0078,
  -37.036,
  -37.0647,
  -37.0938,
  -37.123,
  -37.1522,
  -37.1813,
  -37.2102,
  -37.2388,
  -37.267,
  -37.2949,
  -37.3228,
  -37.3507,
  -37.3788,
  -37.407,
  -37.4353,
  -37.4636,
  -37.4909,
  -37.5196,
  -37.5486,
  -37.5777,
  -37.6066,
  -37.6346,
  -37.6615,
  -37.687,
  -37.7111,
  -37.7342,
  -37.7569,
  -37.7794,
  -37.802,
  -37.8244,
  -37.8465,
  -37.8681,
  -37.8892,
  -37.9097,
  -37.9301,
  -37.9506,
  -37.9715,
  -37.9931,
  -38.0154,
  -38.0385,
  -38.0609,
  -38.0846,
  -38.108,
  -38.1308,
  -38.1525,
  -38.173,
  -38.1925,
  -38.2111,
  -38.2292,
  -38.2469,
  -38.2641,
  -38.2806,
  -38.2965,
  -38.3117,
  -38.3267,
  -38.3415,
  -38.3565,
  -38.3717,
  -38.3875,
  -38.4044,
  -38.4228,
  -38.4435,
  -38.4669,
  -38.4932,
  -38.5215,
  -38.5514,
  -38.5815,
  -38.6111,
  -38.6383,
  -38.6651,
  -38.6906,
  -38.7156,
  -38.7407,
  -38.7663,
  -38.7929,
  -38.8205,
  -38.8496,
  -38.8802,
  -38.912,
  -38.9444,
  -38.9771,
  -39.0097,
  -39.0422,
  -39.0742,
  -39.1056,
  -39.1361,
  -39.1653,
  -39.193,
  -39.2197,
  -39.2453,
  -39.2699,
  -39.2933,
  -39.3156,
  -39.3369,
  -39.3577,
  -39.3781,
  -39.3986,
  -39.4193,
  -39.4401,
  -39.4608,
  -39.48,
  -39.4992,
  -39.5167,
  -39.5321,
  -39.545,
  -39.555,
  -39.5625,
  -39.5679,
  -39.5725,
  -39.5772,
  -39.583,
  -39.5902,
  -39.5988,
  -39.6078,
  -39.6162,
  -39.6232,
  -39.6289,
  -39.6327,
  -39.6347,
  -39.6352,
  -39.6348,
  -39.6334,
  -39.6319,
  -39.631,
  -39.6301,
  -39.6287,
  -39.6261,
  -39.6216,
  -39.6148,
  -39.6055,
  -39.5934,
  -39.5786,
  -39.5611,
  -39.5416,
  -39.5203,
  -39.4976,
  -39.4731,
  -39.4471,
  -39.4196,
  -39.391,
  -39.3607,
  -39.3303,
  -39.2982,
  -39.2634,
  -39.2249,
  -39.1815,
  -39.1326,
  -39.0784,
  -39.0187,
  -38.9542,
  -38.8859,
  -38.8157,
  -38.7459,
  -38.6799,
  -38.6215,
  -38.5734,
  -30.8165,
  -30.8647,
  -30.9118,
  -30.9579,
  -31.0032,
  -31.0481,
  -31.0933,
  -31.139,
  -31.1855,
  -31.2329,
  -31.2808,
  -31.3288,
  -31.3754,
  -31.4221,
  -31.4677,
  -31.5128,
  -31.5579,
  -31.6035,
  -31.6499,
  -31.6969,
  -31.7443,
  -31.7921,
  -31.8398,
  -31.8873,
  -31.9342,
  -31.9805,
  -32.0261,
  -32.0702,
  -32.1152,
  -32.1603,
  -32.2054,
  -32.2507,
  -32.2964,
  -32.3426,
  -32.3891,
  -32.4359,
  -32.4827,
  -32.5294,
  -32.5763,
  -32.6235,
  -32.6719,
  -32.7212,
  -32.7706,
  -32.8218,
  -32.873,
  -32.9241,
  -32.9753,
  -33.0269,
  -33.079,
  -33.1316,
  -33.1845,
  -33.2375,
  -33.2904,
  -33.3436,
  -33.3971,
  -33.451,
  -33.5051,
  -33.5593,
  -33.6125,
  -33.6668,
  -33.7216,
  -33.7768,
  -33.8324,
  -33.8883,
  -33.9442,
  -34.0003,
  -34.056,
  -34.1114,
  -34.1665,
  -34.2204,
  -34.2739,
  -34.3273,
  -34.3804,
  -34.4335,
  -34.4866,
  -34.5385,
  -34.5909,
  -34.6427,
  -34.6947,
  -34.7458,
  -34.7955,
  -34.8435,
  -34.8892,
  -34.9327,
  -34.9752,
  -35.0176,
  -35.0607,
  -35.1048,
  -35.1498,
  -35.1951,
  -35.2401,
  -35.2842,
  -35.3279,
  -35.3706,
  -35.4139,
  -35.457,
  -35.4995,
  -35.541,
  -35.5816,
  -35.6211,
  -35.6593,
  -35.6961,
  -35.7315,
  -35.7657,
  -35.7988,
  -35.8309,
  -35.8618,
  -35.8918,
  -35.9213,
  -35.951,
  -35.9811,
  -36.0117,
  -36.0414,
  -36.0716,
  -36.1012,
  -36.1303,
  -36.1595,
  -36.1891,
  -36.219,
  -36.249,
  -36.2791,
  -36.3094,
  -36.3403,
  -36.3713,
  -36.4021,
  -36.4322,
  -36.4612,
  -36.4893,
  -36.5167,
  -36.544,
  -36.5714,
  -36.5989,
  -36.6257,
  -36.654,
  -36.683,
  -36.7122,
  -36.7412,
  -36.7698,
  -36.798,
  -36.8258,
  -36.8536,
  -36.8812,
  -36.9089,
  -36.9366,
  -36.9644,
  -36.9926,
  -37.0211,
  -37.05,
  -37.0789,
  -37.108,
  -37.1372,
  -37.1664,
  -37.1955,
  -37.2233,
  -37.2517,
  -37.2799,
  -37.3081,
  -37.3362,
  -37.3643,
  -37.3923,
  -37.4203,
  -37.4484,
  -37.4768,
  -37.5056,
  -37.5346,
  -37.563,
  -37.5906,
  -37.6169,
  -37.6416,
  -37.665,
  -37.6875,
  -37.7096,
  -37.7319,
  -37.7542,
  -37.7764,
  -37.7982,
  -37.8194,
  -37.8391,
  -37.8593,
  -37.8792,
  -37.899,
  -37.9192,
  -37.9399,
  -37.9615,
  -37.9839,
  -38.0069,
  -38.0302,
  -38.0534,
  -38.0761,
  -38.0978,
  -38.1183,
  -38.1376,
  -38.1562,
  -38.1742,
  -38.1919,
  -38.2091,
  -38.2258,
  -38.2421,
  -38.258,
  -38.2736,
  -38.2895,
  -38.3052,
  -38.3212,
  -38.3367,
  -38.3543,
  -38.3735,
  -38.3949,
  -38.4189,
  -38.4458,
  -38.4751,
  -38.5057,
  -38.5369,
  -38.5674,
  -38.5967,
  -38.6246,
  -38.6513,
  -38.6772,
  -38.7028,
  -38.7289,
  -38.7557,
  -38.7835,
  -38.8126,
  -38.8432,
  -38.8751,
  -38.9078,
  -38.9407,
  -38.9735,
  -39.006,
  -39.0382,
  -39.0695,
  -39.0998,
  -39.1288,
  -39.1563,
  -39.1825,
  -39.2062,
  -39.2299,
  -39.2522,
  -39.2733,
  -39.2938,
  -39.3138,
  -39.3338,
  -39.3543,
  -39.3751,
  -39.3961,
  -39.4171,
  -39.4374,
  -39.4564,
  -39.4735,
  -39.4885,
  -39.5009,
  -39.5107,
  -39.5182,
  -39.5236,
  -39.5282,
  -39.5328,
  -39.5385,
  -39.5457,
  -39.554,
  -39.5625,
  -39.5709,
  -39.5779,
  -39.5833,
  -39.587,
  -39.5892,
  -39.5898,
  -39.5892,
  -39.5879,
  -39.5864,
  -39.5851,
  -39.5835,
  -39.5814,
  -39.5766,
  -39.5709,
  -39.5629,
  -39.5526,
  -39.5396,
  -39.5242,
  -39.5066,
  -39.4872,
  -39.4663,
  -39.444,
  -39.4195,
  -39.3929,
  -39.3641,
  -39.3338,
  -39.3028,
  -39.2709,
  -39.2377,
  -39.2021,
  -39.1629,
  -39.1191,
  -39.0697,
  -39.0146,
  -38.9541,
  -38.889,
  -38.8204,
  -38.7506,
  -38.6824,
  -38.6191,
  -38.5645,
  -38.5207,
  -30.7478,
  -30.7961,
  -30.8433,
  -30.8896,
  -30.9352,
  -30.9806,
  -31.0263,
  -31.0725,
  -31.1184,
  -31.1659,
  -31.2139,
  -31.2619,
  -31.3096,
  -31.3565,
  -31.4025,
  -31.4482,
  -31.4939,
  -31.5404,
  -31.5875,
  -31.6351,
  -31.6829,
  -31.7306,
  -31.7773,
  -31.8249,
  -31.8718,
  -31.9177,
  -31.9629,
  -32.0075,
  -32.0519,
  -32.0965,
  -32.1414,
  -32.1868,
  -32.2327,
  -32.2796,
  -32.3269,
  -32.3744,
  -32.4217,
  -32.4678,
  -32.5149,
  -32.5626,
  -32.6115,
  -32.6617,
  -32.7129,
  -32.7648,
  -32.8169,
  -32.869,
  -32.9211,
  -32.9736,
  -33.0264,
  -33.0796,
  -33.1331,
  -33.1864,
  -33.2395,
  -33.2917,
  -33.345,
  -33.3986,
  -33.4525,
  -33.5065,
  -33.5605,
  -33.615,
  -33.67,
  -33.7256,
  -33.7816,
  -33.8379,
  -33.8942,
  -33.9503,
  -34.0057,
  -34.0606,
  -34.1146,
  -34.1681,
  -34.2196,
  -34.2718,
  -34.324,
  -34.3763,
  -34.4286,
  -34.481,
  -34.533,
  -34.585,
  -34.6362,
  -34.687,
  -34.7371,
  -34.7856,
  -34.8315,
  -34.8757,
  -34.9189,
  -34.9618,
  -35.005,
  -35.0478,
  -35.092,
  -35.1362,
  -35.18,
  -35.2232,
  -35.2661,
  -35.3091,
  -35.3523,
  -35.395,
  -35.4371,
  -35.4784,
  -35.519,
  -35.5588,
  -35.5974,
  -35.6348,
  -35.6709,
  -35.7058,
  -35.7397,
  -35.7725,
  -35.8031,
  -35.8339,
  -35.8642,
  -35.8945,
  -35.9252,
  -35.9563,
  -35.9872,
  -36.0174,
  -36.0469,
  -36.076,
  -36.1053,
  -36.1351,
  -36.1655,
  -36.196,
  -36.2265,
  -36.2575,
  -36.2889,
  -36.3205,
  -36.3518,
  -36.3812,
  -36.4104,
  -36.4384,
  -36.4658,
  -36.493,
  -36.5201,
  -36.5478,
  -36.5761,
  -36.6051,
  -36.6346,
  -36.6644,
  -36.694,
  -36.7231,
  -36.7515,
  -36.7798,
  -36.8078,
  -36.8359,
  -36.864,
  -36.8922,
  -36.9205,
  -36.9488,
  -36.9763,
  -37.0049,
  -37.0336,
  -37.0626,
  -37.0918,
  -37.1212,
  -37.1507,
  -37.1799,
  -37.2087,
  -37.2372,
  -37.2654,
  -37.2934,
  -37.3213,
  -37.349,
  -37.3765,
  -37.4042,
  -37.4322,
  -37.4607,
  -37.4894,
  -37.5175,
  -37.5448,
  -37.5704,
  -37.5947,
  -37.6164,
  -37.6386,
  -37.6606,
  -37.6827,
  -37.7048,
  -37.7267,
  -37.7483,
  -37.7693,
  -37.7897,
  -37.8096,
  -37.829,
  -37.8484,
  -37.8679,
  -37.8879,
  -37.9087,
  -37.9305,
  -37.9529,
  -37.9759,
  -37.9989,
  -38.0216,
  -38.0435,
  -38.0642,
  -38.0836,
  -38.1022,
  -38.1201,
  -38.1366,
  -38.1538,
  -38.1706,
  -38.1871,
  -38.2037,
  -38.22,
  -38.2368,
  -38.2533,
  -38.2703,
  -38.2878,
  -38.3063,
  -38.3264,
  -38.3486,
  -38.3735,
  -38.4011,
  -38.431,
  -38.4623,
  -38.4943,
  -38.5258,
  -38.5562,
  -38.5853,
  -38.6132,
  -38.6399,
  -38.6664,
  -38.6927,
  -38.7195,
  -38.7473,
  -38.7763,
  -38.8067,
  -38.8376,
  -38.8704,
  -38.9033,
  -38.9362,
  -38.9687,
  -39.0006,
  -39.0318,
  -39.062,
  -39.0908,
  -39.1179,
  -39.1436,
  -39.1677,
  -39.1903,
  -39.2114,
  -39.2315,
  -39.2512,
  -39.2706,
  -39.2906,
  -39.3111,
  -39.3321,
  -39.3533,
  -39.3743,
  -39.3945,
  -39.4132,
  -39.4298,
  -39.4444,
  -39.4566,
  -39.4664,
  -39.4739,
  -39.4797,
  -39.4845,
  -39.4893,
  -39.4951,
  -39.502,
  -39.5099,
  -39.5172,
  -39.5249,
  -39.5315,
  -39.5366,
  -39.5404,
  -39.5427,
  -39.5436,
  -39.5432,
  -39.5419,
  -39.5402,
  -39.5384,
  -39.5361,
  -39.5328,
  -39.528,
  -39.5211,
  -39.5121,
  -39.5009,
  -39.4872,
  -39.4712,
  -39.4534,
  -39.4342,
  -39.4137,
  -39.3915,
  -39.3671,
  -39.3399,
  -39.3098,
  -39.2779,
  -39.2453,
  -39.2119,
  -39.1773,
  -39.1412,
  -39.1015,
  -39.0574,
  -39.0078,
  -38.9524,
  -38.8915,
  -38.826,
  -38.7575,
  -38.6882,
  -38.6215,
  -38.5609,
  -38.5099,
  -38.4704,
  -30.6807,
  -30.7289,
  -30.7763,
  -30.8219,
  -30.868,
  -30.914,
  -30.9603,
  -31.0069,
  -31.0541,
  -31.1017,
  -31.1497,
  -31.1977,
  -31.2455,
  -31.2926,
  -31.3391,
  -31.3852,
  -31.4318,
  -31.479,
  -31.5257,
  -31.5737,
  -31.6218,
  -31.6696,
  -31.7175,
  -31.7649,
  -31.8117,
  -31.8575,
  -31.9022,
  -31.9463,
  -31.9902,
  -32.0344,
  -32.0791,
  -32.1247,
  -32.1704,
  -32.218,
  -32.2662,
  -32.3144,
  -32.3623,
  -32.41,
  -32.4577,
  -32.5061,
  -32.5555,
  -32.6064,
  -32.6583,
  -32.7107,
  -32.7635,
  -32.8163,
  -32.8691,
  -32.9223,
  -32.9748,
  -33.0286,
  -33.0824,
  -33.1361,
  -33.1894,
  -33.2426,
  -33.2957,
  -33.349,
  -33.4024,
  -33.4561,
  -33.5101,
  -33.5646,
  -33.6199,
  -33.6759,
  -33.7323,
  -33.7888,
  -33.8439,
  -33.8997,
  -33.9549,
  -34.0092,
  -34.0626,
  -34.1151,
  -34.1669,
  -34.2185,
  -34.2698,
  -34.3214,
  -34.3732,
  -34.4251,
  -34.4769,
  -34.5284,
  -34.5794,
  -34.63,
  -34.6795,
  -34.7271,
  -34.7737,
  -34.8188,
  -34.863,
  -34.9064,
  -34.9496,
  -34.9929,
  -35.0362,
  -35.0792,
  -35.1217,
  -35.1638,
  -35.206,
  -35.2486,
  -35.2914,
  -35.3339,
  -35.3756,
  -35.4167,
  -35.4572,
  -35.496,
  -35.5348,
  -35.5726,
  -35.6091,
  -35.6446,
  -35.6792,
  -35.7126,
  -35.745,
  -35.7766,
  -35.8076,
  -35.8386,
  -35.8698,
  -35.9011,
  -35.9321,
  -35.9624,
  -35.9919,
  -36.0211,
  -36.0505,
  -36.0805,
  -36.1111,
  -36.1409,
  -36.172,
  -36.2036,
  -36.2355,
  -36.2676,
  -36.2992,
  -36.3299,
  -36.3593,
  -36.3875,
  -36.4149,
  -36.442,
  -36.4693,
  -36.4972,
  -36.526,
  -36.5555,
  -36.5856,
  -36.6159,
  -36.6458,
  -36.6752,
  -36.704,
  -36.7315,
  -36.76,
  -36.7884,
  -36.8169,
  -36.8455,
  -36.8742,
  -36.9029,
  -36.9317,
  -36.9604,
  -36.9892,
  -37.0182,
  -37.0474,
  -37.0769,
  -37.1066,
  -37.136,
  -37.1651,
  -37.1937,
  -37.2218,
  -37.2495,
  -37.2769,
  -37.3041,
  -37.3311,
  -37.3571,
  -37.3846,
  -37.4127,
  -37.441,
  -37.4691,
  -37.4959,
  -37.5216,
  -37.5456,
  -37.5684,
  -37.5903,
  -37.6121,
  -37.6339,
  -37.6557,
  -37.6772,
  -37.6985,
  -37.7193,
  -37.7395,
  -37.7591,
  -37.7783,
  -37.7973,
  -37.8163,
  -37.8359,
  -37.8562,
  -37.8772,
  -37.8994,
  -37.921,
  -37.9439,
  -37.9666,
  -37.9886,
  -38.0094,
  -38.029,
  -38.0476,
  -38.0656,
  -38.0829,
  -38.1,
  -38.117,
  -38.1337,
  -38.1508,
  -38.168,
  -38.1854,
  -38.2031,
  -38.2211,
  -38.2397,
  -38.2593,
  -38.2803,
  -38.3036,
  -38.3294,
  -38.3577,
  -38.3884,
  -38.4205,
  -38.453,
  -38.4853,
  -38.5166,
  -38.5457,
  -38.5745,
  -38.6019,
  -38.629,
  -38.6555,
  -38.6824,
  -38.7102,
  -38.739,
  -38.7693,
  -38.8012,
  -38.8338,
  -38.8669,
  -38.8996,
  -38.932,
  -38.9637,
  -38.9947,
  -39.0246,
  -39.0533,
  -39.0804,
  -39.1057,
  -39.1291,
  -39.151,
  -39.1712,
  -39.1904,
  -39.2096,
  -39.2288,
  -39.2485,
  -39.269,
  -39.2899,
  -39.3109,
  -39.3315,
  -39.3513,
  -39.3684,
  -39.3847,
  -39.399,
  -39.4109,
  -39.4208,
  -39.4288,
  -39.4351,
  -39.4404,
  -39.4457,
  -39.4517,
  -39.4586,
  -39.4662,
  -39.474,
  -39.4811,
  -39.4872,
  -39.4918,
  -39.4955,
  -39.4979,
  -39.4989,
  -39.4987,
  -39.4975,
  -39.4957,
  -39.4934,
  -39.4903,
  -39.486,
  -39.48,
  -39.472,
  -39.4621,
  -39.4498,
  -39.4356,
  -39.4191,
  -39.4011,
  -39.3819,
  -39.3614,
  -39.3392,
  -39.3143,
  -39.2863,
  -39.2552,
  -39.222,
  -39.1877,
  -39.1529,
  -39.1165,
  -39.0797,
  -39.04,
  -38.9958,
  -38.9463,
  -38.8909,
  -38.8298,
  -38.764,
  -38.6954,
  -38.6266,
  -38.561,
  -38.5024,
  -38.4542,
  -38.418,
  -30.6143,
  -30.6624,
  -30.71,
  -30.757,
  -30.8036,
  -30.8502,
  -30.897,
  -30.9441,
  -30.9914,
  -31.039,
  -31.0869,
  -31.1349,
  -31.1826,
  -31.2289,
  -31.2759,
  -31.3227,
  -31.3699,
  -31.4177,
  -31.466,
  -31.5144,
  -31.5627,
  -31.6106,
  -31.6587,
  -31.706,
  -31.7527,
  -31.7982,
  -31.8427,
  -31.8864,
  -31.9289,
  -31.9729,
  -32.0176,
  -32.0637,
  -32.1109,
  -32.1594,
  -32.2085,
  -32.2576,
  -32.3063,
  -32.3546,
  -32.4031,
  -32.4522,
  -32.5025,
  -32.554,
  -32.6065,
  -32.6584,
  -32.7116,
  -32.7648,
  -32.8183,
  -32.8721,
  -32.9261,
  -32.9803,
  -33.0344,
  -33.0884,
  -33.1419,
  -33.1952,
  -33.2481,
  -33.301,
  -33.3539,
  -33.4072,
  -33.4609,
  -33.5145,
  -33.57,
  -33.6262,
  -33.6827,
  -33.7391,
  -33.7951,
  -33.8504,
  -33.9051,
  -33.9588,
  -34.0116,
  -34.0637,
  -34.1151,
  -34.1661,
  -34.217,
  -34.268,
  -34.3194,
  -34.3707,
  -34.4211,
  -34.4724,
  -34.5229,
  -34.5731,
  -34.6225,
  -34.6708,
  -34.7179,
  -34.7638,
  -34.8087,
  -34.8526,
  -34.8958,
  -34.9383,
  -34.9805,
  -35.0221,
  -35.0633,
  -35.1045,
  -35.1462,
  -35.1886,
  -35.2301,
  -35.2724,
  -35.3141,
  -35.3551,
  -35.3951,
  -35.4347,
  -35.4736,
  -35.5114,
  -35.5482,
  -35.5841,
  -35.619,
  -35.653,
  -35.6861,
  -35.7184,
  -35.7501,
  -35.7816,
  -35.8132,
  -35.8446,
  -35.8746,
  -35.9051,
  -35.9348,
  -35.9642,
  -35.9938,
  -36.024,
  -36.0547,
  -36.0858,
  -36.1175,
  -36.1495,
  -36.1819,
  -36.2143,
  -36.2462,
  -36.2772,
  -36.307,
  -36.3355,
  -36.3632,
  -36.3904,
  -36.418,
  -36.4463,
  -36.4744,
  -36.5044,
  -36.5349,
  -36.5655,
  -36.5958,
  -36.6255,
  -36.6547,
  -36.6832,
  -36.7118,
  -36.7405,
  -36.7693,
  -36.7984,
  -36.8275,
  -36.8569,
  -36.8861,
  -36.9153,
  -36.9444,
  -36.9736,
  -37.0031,
  -37.0327,
  -37.0624,
  -37.0919,
  -37.1199,
  -37.1484,
  -37.1762,
  -37.2034,
  -37.2302,
  -37.2566,
  -37.2828,
  -37.3092,
  -37.336,
  -37.3636,
  -37.3915,
  -37.4193,
  -37.4463,
  -37.472,
  -37.4962,
  -37.5192,
  -37.5412,
  -37.5627,
  -37.5841,
  -37.6055,
  -37.6269,
  -37.6478,
  -37.6682,
  -37.6881,
  -37.7065,
  -37.7256,
  -37.7445,
  -37.7633,
  -37.7825,
  -37.8023,
  -37.8231,
  -37.8447,
  -37.8669,
  -37.8897,
  -37.9124,
  -37.9345,
  -37.9555,
  -37.9752,
  -37.9939,
  -38.0117,
  -38.0289,
  -38.046,
  -38.063,
  -38.0803,
  -38.098,
  -38.116,
  -38.1342,
  -38.1528,
  -38.1718,
  -38.1916,
  -38.2115,
  -38.2339,
  -38.2583,
  -38.2853,
  -38.3147,
  -38.346,
  -38.3788,
  -38.4119,
  -38.4448,
  -38.4769,
  -38.5076,
  -38.537,
  -38.5652,
  -38.5924,
  -38.6193,
  -38.6463,
  -38.674,
  -38.7026,
  -38.7327,
  -38.7643,
  -38.797,
  -38.83,
  -38.8627,
  -38.8948,
  -38.9263,
  -38.957,
  -38.9868,
  -39.0154,
  -39.0423,
  -39.0674,
  -39.0905,
  -39.1106,
  -39.1301,
  -39.1489,
  -39.1678,
  -39.187,
  -39.2067,
  -39.227,
  -39.2476,
  -39.2681,
  -39.2881,
  -39.3071,
  -39.3246,
  -39.3404,
  -39.3541,
  -39.366,
  -39.3761,
  -39.3846,
  -39.3917,
  -39.3978,
  -39.4038,
  -39.41,
  -39.4171,
  -39.4246,
  -39.4317,
  -39.4382,
  -39.4435,
  -39.4478,
  -39.451,
  -39.4533,
  -39.4545,
  -39.4546,
  -39.4537,
  -39.4518,
  -39.4491,
  -39.4453,
  -39.44,
  -39.433,
  -39.423,
  -39.412,
  -39.3992,
  -39.3841,
  -39.3672,
  -39.349,
  -39.3296,
  -39.3088,
  -39.2861,
  -39.2607,
  -39.2317,
  -39.1995,
  -39.1651,
  -39.1297,
  -39.0941,
  -39.058,
  -39.0209,
  -38.9812,
  -38.9373,
  -38.8879,
  -38.8324,
  -38.7708,
  -38.7045,
  -38.6353,
  -38.5662,
  -38.5011,
  -38.4438,
  -38.3975,
  -38.3641,
  -30.5506,
  -30.5986,
  -30.6463,
  -30.6937,
  -30.7409,
  -30.788,
  -30.8353,
  -30.8827,
  -30.9292,
  -30.9769,
  -31.0246,
  -31.0723,
  -31.1198,
  -31.1671,
  -31.2143,
  -31.2617,
  -31.3096,
  -31.3582,
  -31.4069,
  -31.4558,
  -31.5044,
  -31.5528,
  -31.6009,
  -31.6474,
  -31.694,
  -31.7393,
  -31.7835,
  -31.8269,
  -31.8703,
  -31.9143,
  -31.9594,
  -32.0058,
  -32.0539,
  -32.1032,
  -32.1532,
  -32.2031,
  -32.2526,
  -32.3017,
  -32.3499,
  -32.3999,
  -32.451,
  -32.503,
  -32.5559,
  -32.609,
  -32.6625,
  -32.7162,
  -32.7702,
  -32.8245,
  -32.8789,
  -32.9334,
  -32.9879,
  -33.0421,
  -33.0959,
  -33.1492,
  -33.2009,
  -33.2534,
  -33.3058,
  -33.3586,
  -33.4119,
  -33.4665,
  -33.522,
  -33.5782,
  -33.6346,
  -33.6907,
  -33.7462,
  -33.801,
  -33.855,
  -33.9081,
  -33.9606,
  -34.0123,
  -34.0625,
  -34.1134,
  -34.1641,
  -34.2148,
  -34.2657,
  -34.3168,
  -34.3678,
  -34.4188,
  -34.469,
  -34.5183,
  -34.5674,
  -34.6155,
  -34.6629,
  -34.7093,
  -34.7547,
  -34.7987,
  -34.8417,
  -34.8835,
  -34.9234,
  -34.9636,
  -35.0035,
  -35.0439,
  -35.0856,
  -35.1279,
  -35.1704,
  -35.2126,
  -35.254,
  -35.2947,
  -35.3347,
  -35.3741,
  -35.4127,
  -35.4504,
  -35.4872,
  -35.5231,
  -35.5582,
  -35.5926,
  -35.6252,
  -35.6581,
  -35.6905,
  -35.7225,
  -35.7544,
  -35.7859,
  -35.8171,
  -35.8477,
  -35.8777,
  -35.9075,
  -35.9374,
  -35.9677,
  -35.9986,
  -36.0301,
  -36.0621,
  -36.0947,
  -36.1273,
  -36.16,
  -36.1921,
  -36.2233,
  -36.2526,
  -36.2817,
  -36.3099,
  -36.3376,
  -36.3655,
  -36.3941,
  -36.4236,
  -36.4539,
  -36.4846,
  -36.5155,
  -36.5459,
  -36.5758,
  -36.6053,
  -36.6341,
  -36.663,
  -36.6918,
  -36.7208,
  -36.7501,
  -36.7798,
  -36.8097,
  -36.8395,
  -36.8683,
  -36.898,
  -36.9277,
  -36.9574,
  -36.9871,
  -37.0168,
  -37.0464,
  -37.0754,
  -37.1036,
  -37.131,
  -37.1575,
  -37.1834,
  -37.2089,
  -37.2341,
  -37.2596,
  -37.2857,
  -37.3126,
  -37.3401,
  -37.3677,
  -37.3948,
  -37.4209,
  -37.4456,
  -37.469,
  -37.4902,
  -37.5117,
  -37.5328,
  -37.5537,
  -37.5746,
  -37.5951,
  -37.6152,
  -37.635,
  -37.6543,
  -37.6733,
  -37.6923,
  -37.7111,
  -37.7302,
  -37.7497,
  -37.7699,
  -37.7911,
  -37.8129,
  -37.8353,
  -37.8578,
  -37.8797,
  -37.9007,
  -37.9205,
  -37.939,
  -37.9567,
  -37.9737,
  -37.9896,
  -38.0069,
  -38.0248,
  -38.0434,
  -38.0624,
  -38.0818,
  -38.1015,
  -38.1217,
  -38.1427,
  -38.1648,
  -38.1885,
  -38.2143,
  -38.2426,
  -38.2732,
  -38.3055,
  -38.3389,
  -38.3726,
  -38.4059,
  -38.4383,
  -38.4694,
  -38.4992,
  -38.5278,
  -38.5554,
  -38.5825,
  -38.6095,
  -38.6371,
  -38.6657,
  -38.6957,
  -38.7272,
  -38.7587,
  -38.7917,
  -38.8243,
  -38.8563,
  -38.8876,
  -38.918,
  -38.9476,
  -38.9761,
  -39.003,
  -39.0279,
  -39.0508,
  -39.0717,
  -39.0911,
  -39.1097,
  -39.1284,
  -39.1476,
  -39.1673,
  -39.1872,
  -39.2072,
  -39.2267,
  -39.2458,
  -39.2639,
  -39.2806,
  -39.2957,
  -39.3091,
  -39.321,
  -39.3315,
  -39.3406,
  -39.3485,
  -39.3556,
  -39.3623,
  -39.3692,
  -39.3763,
  -39.3835,
  -39.3902,
  -39.3949,
  -39.3996,
  -39.4032,
  -39.4061,
  -39.4082,
  -39.4094,
  -39.4097,
  -39.4089,
  -39.4072,
  -39.4042,
  -39.3997,
  -39.3936,
  -39.3857,
  -39.3758,
  -39.3641,
  -39.3505,
  -39.335,
  -39.3179,
  -39.2994,
  -39.2796,
  -39.2584,
  -39.235,
  -39.2086,
  -39.1787,
  -39.1456,
  -39.1104,
  -39.0743,
  -39.0379,
  -39.0016,
  -38.9645,
  -38.9249,
  -38.8814,
  -38.832,
  -38.7759,
  -38.7136,
  -38.646,
  -38.5755,
  -38.5053,
  -38.4395,
  -38.3825,
  -38.3375,
  -38.3063,
  -30.4887,
  -30.5365,
  -30.5842,
  -30.6319,
  -30.6786,
  -30.7262,
  -30.774,
  -30.8219,
  -30.8696,
  -30.9172,
  -30.9646,
  -31.0119,
  -31.0591,
  -31.1062,
  -31.1536,
  -31.2015,
  -31.25,
  -31.299,
  -31.3474,
  -31.3969,
  -31.4461,
  -31.4951,
  -31.5434,
  -31.591,
  -31.6375,
  -31.6827,
  -31.7268,
  -31.7702,
  -31.8139,
  -31.8582,
  -31.9038,
  -31.9508,
  -31.9995,
  -32.0487,
  -32.0995,
  -32.1501,
  -32.2003,
  -32.2502,
  -32.3002,
  -32.3508,
  -32.4024,
  -32.4548,
  -32.5077,
  -32.5611,
  -32.6149,
  -32.6689,
  -32.7235,
  -32.7783,
  -32.8331,
  -32.8869,
  -32.9416,
  -32.996,
  -33.0499,
  -33.1032,
  -33.1558,
  -33.2078,
  -33.2597,
  -33.3119,
  -33.3649,
  -33.4192,
  -33.4743,
  -33.5304,
  -33.5864,
  -33.6421,
  -33.6972,
  -33.7503,
  -33.8036,
  -33.8562,
  -33.9083,
  -33.9598,
  -34.0108,
  -34.0617,
  -34.1124,
  -34.1632,
  -34.2142,
  -34.2651,
  -34.3156,
  -34.366,
  -34.4156,
  -34.4648,
  -34.513,
  -34.5609,
  -34.6073,
  -34.6537,
  -34.6992,
  -34.7432,
  -34.7855,
  -34.8266,
  -34.8662,
  -34.9055,
  -34.9446,
  -34.9848,
  -35.0261,
  -35.0685,
  -35.1109,
  -35.153,
  -35.1944,
  -35.235,
  -35.2748,
  -35.314,
  -35.3512,
  -35.3887,
  -35.4253,
  -35.4611,
  -35.4962,
  -35.5307,
  -35.5647,
  -35.5982,
  -35.6312,
  -35.6637,
  -35.6958,
  -35.7275,
  -35.7589,
  -35.7897,
  -35.8201,
  -35.8504,
  -35.8806,
  -35.9112,
  -35.9423,
  -35.9731,
  -36.0056,
  -36.0386,
  -36.0715,
  -36.1041,
  -36.1362,
  -36.1677,
  -36.1984,
  -36.2283,
  -36.2572,
  -36.2855,
  -36.3137,
  -36.3427,
  -36.3724,
  -36.4029,
  -36.4337,
  -36.4646,
  -36.4952,
  -36.5254,
  -36.5552,
  -36.5843,
  -36.6124,
  -36.6412,
  -36.6705,
  -36.7002,
  -36.7303,
  -36.7607,
  -36.7912,
  -36.8216,
  -36.852,
  -36.8822,
  -36.9123,
  -36.9422,
  -36.9719,
  -37.0014,
  -37.0303,
  -37.0582,
  -37.0851,
  -37.1109,
  -37.1357,
  -37.16,
  -37.1842,
  -37.2089,
  -37.2333,
  -37.2594,
  -37.2864,
  -37.3137,
  -37.3409,
  -37.3675,
  -37.3929,
  -37.4169,
  -37.4395,
  -37.461,
  -37.4818,
  -37.5022,
  -37.5225,
  -37.5427,
  -37.5626,
  -37.5822,
  -37.6016,
  -37.6208,
  -37.6399,
  -37.6588,
  -37.6779,
  -37.6973,
  -37.7172,
  -37.7378,
  -37.759,
  -37.7798,
  -37.8017,
  -37.8231,
  -37.8436,
  -37.863,
  -37.8813,
  -37.8986,
  -37.9155,
  -37.9325,
  -37.9502,
  -37.9689,
  -37.9887,
  -38.0091,
  -38.0299,
  -38.0508,
  -38.0723,
  -38.0945,
  -38.1179,
  -38.1429,
  -38.1701,
  -38.1998,
  -38.2317,
  -38.2651,
  -38.2993,
  -38.3334,
  -38.3671,
  -38.3996,
  -38.4309,
  -38.46,
  -38.4889,
  -38.5167,
  -38.5439,
  -38.571,
  -38.5986,
  -38.6273,
  -38.6573,
  -38.6887,
  -38.7212,
  -38.7541,
  -38.7868,
  -38.8187,
  -38.8499,
  -38.8801,
  -38.9095,
  -38.9378,
  -38.9644,
  -38.9893,
  -39.0121,
  -39.033,
  -39.0525,
  -39.0713,
  -39.0902,
  -39.1094,
  -39.1288,
  -39.1483,
  -39.1674,
  -39.1859,
  -39.2039,
  -39.221,
  -39.237,
  -39.2505,
  -39.2636,
  -39.2754,
  -39.2863,
  -39.296,
  -39.3048,
  -39.3127,
  -39.3202,
  -39.3276,
  -39.3348,
  -39.3417,
  -39.3479,
  -39.3531,
  -39.3572,
  -39.3603,
  -39.3628,
  -39.3647,
  -39.3657,
  -39.366,
  -39.3654,
  -39.3636,
  -39.3604,
  -39.3554,
  -39.3486,
  -39.3399,
  -39.3293,
  -39.3169,
  -39.3028,
  -39.287,
  -39.2698,
  -39.2512,
  -39.2314,
  -39.2096,
  -39.1855,
  -39.1582,
  -39.1275,
  -39.0937,
  -39.0578,
  -39.0213,
  -38.9846,
  -38.9482,
  -38.9103,
  -38.871,
  -38.827,
  -38.7773,
  -38.7207,
  -38.657,
  -38.5872,
  -38.5145,
  -38.4422,
  -38.3749,
  -38.317,
  -38.2723,
  -38.2429,
  -30.4271,
  -30.4746,
  -30.5224,
  -30.5704,
  -30.6184,
  -30.6666,
  -30.7149,
  -30.7632,
  -30.8112,
  -30.8589,
  -30.9061,
  -30.953,
  -30.9998,
  -31.0457,
  -31.0931,
  -31.1412,
  -31.1901,
  -31.2397,
  -31.2898,
  -31.3401,
  -31.3901,
  -31.4396,
  -31.4883,
  -31.536,
  -31.5824,
  -31.6275,
  -31.6716,
  -31.7154,
  -31.7585,
  -31.8033,
  -31.8499,
  -31.8977,
  -31.9469,
  -31.9978,
  -32.0492,
  -32.1005,
  -32.1514,
  -32.2021,
  -32.2527,
  -32.3038,
  -32.3557,
  -32.4082,
  -32.4611,
  -32.5147,
  -32.5676,
  -32.622,
  -32.677,
  -32.7322,
  -32.7873,
  -32.8424,
  -32.8971,
  -32.9516,
  -33.0055,
  -33.0588,
  -33.1112,
  -33.163,
  -33.2147,
  -33.2665,
  -33.3191,
  -33.3729,
  -33.4265,
  -33.482,
  -33.5375,
  -33.5925,
  -33.6468,
  -33.7004,
  -33.7531,
  -33.8052,
  -33.8568,
  -33.908,
  -33.9591,
  -34.0099,
  -34.0608,
  -34.1117,
  -34.1627,
  -34.2134,
  -34.2636,
  -34.3121,
  -34.3609,
  -34.4094,
  -34.4572,
  -34.5047,
  -34.5517,
  -34.5982,
  -34.6437,
  -34.6875,
  -34.7294,
  -34.7696,
  -34.8086,
  -34.8471,
  -34.8859,
  -34.926,
  -34.9673,
  -35.0094,
  -35.0507,
  -35.0926,
  -35.1339,
  -35.1744,
  -35.2142,
  -35.2532,
  -35.2913,
  -35.3286,
  -35.3651,
  -35.4007,
  -35.4357,
  -35.4703,
  -35.5045,
  -35.5384,
  -35.5719,
  -35.6049,
  -35.6374,
  -35.6694,
  -35.7008,
  -35.7309,
  -35.7618,
  -35.7924,
  -35.8231,
  -35.854,
  -35.8853,
  -35.9175,
  -35.9503,
  -35.9835,
  -36.0165,
  -36.0491,
  -36.0812,
  -36.1129,
  -36.144,
  -36.1745,
  -36.2041,
  -36.2331,
  -36.2618,
  -36.291,
  -36.3209,
  -36.3503,
  -36.381,
  -36.4118,
  -36.4425,
  -36.4728,
  -36.5027,
  -36.5324,
  -36.5617,
  -36.5912,
  -36.621,
  -36.6512,
  -36.6818,
  -36.7128,
  -36.7439,
  -36.7749,
  -36.8056,
  -36.8361,
  -36.8664,
  -36.8965,
  -36.9263,
  -36.9557,
  -36.9845,
  -37.0111,
  -37.0374,
  -37.0624,
  -37.0863,
  -37.1095,
  -37.1327,
  -37.1564,
  -37.181,
  -37.2064,
  -37.2328,
  -37.2598,
  -37.2871,
  -37.314,
  -37.34,
  -37.3647,
  -37.3878,
  -37.4095,
  -37.4302,
  -37.4503,
  -37.4701,
  -37.49,
  -37.5096,
  -37.5292,
  -37.5487,
  -37.5672,
  -37.5865,
  -37.6056,
  -37.6247,
  -37.6441,
  -37.6636,
  -37.6836,
  -37.7042,
  -37.725,
  -37.7459,
  -37.7665,
  -37.7862,
  -37.8049,
  -37.8226,
  -37.8397,
  -37.8564,
  -37.8737,
  -37.8921,
  -37.9117,
  -37.9326,
  -37.9545,
  -37.9767,
  -37.9993,
  -38.0224,
  -38.0461,
  -38.0708,
  -38.0962,
  -38.1249,
  -38.156,
  -38.1892,
  -38.2236,
  -38.2587,
  -38.2933,
  -38.3269,
  -38.3597,
  -38.3912,
  -38.4215,
  -38.4504,
  -38.4784,
  -38.5058,
  -38.5331,
  -38.5609,
  -38.5897,
  -38.6198,
  -38.6511,
  -38.6836,
  -38.7165,
  -38.7492,
  -38.7812,
  -38.8123,
  -38.8424,
  -38.8716,
  -38.8995,
  -38.9258,
  -38.9505,
  -38.9735,
  -38.9947,
  -39.0135,
  -39.0326,
  -39.0517,
  -39.0708,
  -39.0899,
  -39.1087,
  -39.127,
  -39.1446,
  -39.1617,
  -39.178,
  -39.1933,
  -39.2074,
  -39.2203,
  -39.2322,
  -39.2434,
  -39.2537,
  -39.2632,
  -39.2717,
  -39.2796,
  -39.2873,
  -39.2944,
  -39.3009,
  -39.3067,
  -39.3113,
  -39.3149,
  -39.3177,
  -39.32,
  -39.3216,
  -39.3225,
  -39.3229,
  -39.3222,
  -39.3202,
  -39.3166,
  -39.3112,
  -39.3037,
  -39.2944,
  -39.2832,
  -39.2704,
  -39.255,
  -39.2391,
  -39.222,
  -39.2034,
  -39.1834,
  -39.1614,
  -39.1367,
  -39.1087,
  -39.0774,
  -39.0432,
  -39.0072,
  -38.9705,
  -38.9339,
  -38.8975,
  -38.8606,
  -38.8213,
  -38.7775,
  -38.7271,
  -38.6691,
  -38.6031,
  -38.5306,
  -38.4545,
  -38.379,
  -38.3091,
  -38.2496,
  -38.2049,
  -38.1769,
  -30.3677,
  -30.4151,
  -30.4628,
  -30.5109,
  -30.5592,
  -30.6078,
  -30.6567,
  -30.7056,
  -30.7542,
  -30.8012,
  -30.8484,
  -30.895,
  -30.9415,
  -30.9882,
  -31.0356,
  -31.0838,
  -31.1329,
  -31.183,
  -31.2338,
  -31.2849,
  -31.3358,
  -31.386,
  -31.4351,
  -31.4817,
  -31.528,
  -31.5731,
  -31.6174,
  -31.6616,
  -31.7064,
  -31.7522,
  -31.7996,
  -31.8483,
  -31.8984,
  -31.9499,
  -32.0018,
  -32.0537,
  -32.1052,
  -32.1564,
  -32.2076,
  -32.2579,
  -32.3099,
  -32.3623,
  -32.4152,
  -32.4686,
  -32.5226,
  -32.5774,
  -32.6327,
  -32.6881,
  -32.7435,
  -32.7985,
  -32.8532,
  -32.9076,
  -32.9615,
  -33.0147,
  -33.0661,
  -33.1179,
  -33.1694,
  -33.221,
  -33.2733,
  -33.3266,
  -33.3807,
  -33.4352,
  -33.4899,
  -33.5442,
  -33.5977,
  -33.6504,
  -33.7024,
  -33.7539,
  -33.8051,
  -33.856,
  -33.9071,
  -33.9569,
  -34.0079,
  -34.059,
  -34.1102,
  -34.1607,
  -34.2104,
  -34.2592,
  -34.3071,
  -34.3545,
  -34.4019,
  -34.4491,
  -34.4961,
  -34.5425,
  -34.5876,
  -34.6312,
  -34.6727,
  -34.7123,
  -34.7498,
  -34.7879,
  -34.8268,
  -34.8668,
  -34.9081,
  -34.95,
  -34.9922,
  -35.0339,
  -35.075,
  -35.1155,
  -35.1552,
  -35.1942,
  -35.2323,
  -35.2695,
  -35.306,
  -35.3417,
  -35.3767,
  -35.4113,
  -35.4456,
  -35.4788,
  -35.5127,
  -35.5461,
  -35.5788,
  -35.611,
  -35.6426,
  -35.674,
  -35.7052,
  -35.7363,
  -35.7673,
  -35.7986,
  -35.8303,
  -35.8628,
  -35.8961,
  -35.9294,
  -35.9626,
  -35.9949,
  -36.0268,
  -36.0584,
  -36.0897,
  -36.1195,
  -36.1498,
  -36.1794,
  -36.2086,
  -36.2381,
  -36.268,
  -36.2982,
  -36.3288,
  -36.3594,
  -36.3901,
  -36.4206,
  -36.4508,
  -36.4809,
  -36.5108,
  -36.5409,
  -36.5715,
  -36.6025,
  -36.6338,
  -36.6653,
  -36.6967,
  -36.7279,
  -36.7577,
  -36.7882,
  -36.8184,
  -36.8486,
  -36.8785,
  -36.9079,
  -36.9365,
  -36.9639,
  -36.9898,
  -37.0143,
  -37.0373,
  -37.0597,
  -37.0819,
  -37.1047,
  -37.1283,
  -37.1531,
  -37.1789,
  -37.2056,
  -37.2328,
  -37.26,
  -37.2865,
  -37.3116,
  -37.3352,
  -37.3562,
  -37.377,
  -37.3969,
  -37.4165,
  -37.436,
  -37.4556,
  -37.4752,
  -37.4949,
  -37.5145,
  -37.534,
  -37.5534,
  -37.5727,
  -37.5918,
  -37.6108,
  -37.6303,
  -37.6501,
  -37.6699,
  -37.6897,
  -37.7091,
  -37.7278,
  -37.7458,
  -37.763,
  -37.7797,
  -37.7964,
  -37.8141,
  -37.8322,
  -37.853,
  -37.8751,
  -37.8983,
  -37.9221,
  -37.9464,
  -37.971,
  -37.9963,
  -38.0226,
  -38.0505,
  -38.0806,
  -38.1132,
  -38.1476,
  -38.1828,
  -38.2185,
  -38.2536,
  -38.2878,
  -38.3207,
  -38.3523,
  -38.3827,
  -38.4117,
  -38.4399,
  -38.4677,
  -38.4953,
  -38.5233,
  -38.5523,
  -38.5825,
  -38.6139,
  -38.6463,
  -38.6791,
  -38.7109,
  -38.743,
  -38.7743,
  -38.8044,
  -38.8332,
  -38.8607,
  -38.8868,
  -38.9113,
  -38.9346,
  -38.9562,
  -38.9769,
  -38.9962,
  -39.0153,
  -39.034,
  -39.0525,
  -39.0707,
  -39.0882,
  -39.1051,
  -39.1215,
  -39.1373,
  -39.1522,
  -39.166,
  -39.1788,
  -39.1907,
  -39.202,
  -39.2126,
  -39.2224,
  -39.2315,
  -39.2396,
  -39.2472,
  -39.2539,
  -39.26,
  -39.2653,
  -39.2695,
  -39.2729,
  -39.2746,
  -39.2767,
  -39.2781,
  -39.279,
  -39.2793,
  -39.2785,
  -39.2763,
  -39.2723,
  -39.2664,
  -39.2584,
  -39.2486,
  -39.2369,
  -39.2238,
  -39.2093,
  -39.1936,
  -39.1767,
  -39.1583,
  -39.1382,
  -39.1159,
  -39.0907,
  -39.0625,
  -39.0311,
  -38.997,
  -38.9613,
  -38.9247,
  -38.8881,
  -38.8517,
  -38.8148,
  -38.7751,
  -38.7308,
  -38.6796,
  -38.6198,
  -38.5512,
  -38.4752,
  -38.395,
  -38.3153,
  -38.242,
  -38.1803,
  -38.1349,
  -38.1084,
  -30.3091,
  -30.3564,
  -30.4042,
  -30.4524,
  -30.4999,
  -30.549,
  -30.5984,
  -30.6481,
  -30.6973,
  -30.7458,
  -30.7934,
  -30.8401,
  -30.8867,
  -30.9333,
  -30.9806,
  -31.0289,
  -31.0781,
  -31.1286,
  -31.18,
  -31.2308,
  -31.2826,
  -31.3332,
  -31.3826,
  -31.4304,
  -31.4766,
  -31.5217,
  -31.5663,
  -31.611,
  -31.6566,
  -31.7035,
  -31.752,
  -31.8017,
  -31.8527,
  -31.9046,
  -31.9562,
  -32.0084,
  -32.0603,
  -32.1122,
  -32.1636,
  -32.2153,
  -32.2673,
  -32.3197,
  -32.3725,
  -32.4258,
  -32.4799,
  -32.5345,
  -32.5897,
  -32.6452,
  -32.7004,
  -32.7543,
  -32.8088,
  -32.863,
  -32.9168,
  -32.9701,
  -33.0227,
  -33.0746,
  -33.1262,
  -33.1778,
  -33.2298,
  -33.2826,
  -33.3359,
  -33.3895,
  -33.443,
  -33.4962,
  -33.5488,
  -33.6008,
  -33.6511,
  -33.702,
  -33.7527,
  -33.8034,
  -33.8541,
  -33.9049,
  -33.956,
  -34.0071,
  -34.058,
  -34.1084,
  -34.1576,
  -34.2057,
  -34.2529,
  -34.2997,
  -34.3465,
  -34.3934,
  -34.4402,
  -34.4855,
  -34.5307,
  -34.5741,
  -34.6154,
  -34.6549,
  -34.6932,
  -34.7313,
  -34.7701,
  -34.8101,
  -34.8512,
  -34.893,
  -34.935,
  -34.9767,
  -35.0177,
  -35.0581,
  -35.0977,
  -35.1366,
  -35.1747,
  -35.2112,
  -35.2478,
  -35.2838,
  -35.3191,
  -35.3538,
  -35.3882,
  -35.4224,
  -35.4564,
  -35.49,
  -35.5229,
  -35.5551,
  -35.5869,
  -35.6184,
  -35.6499,
  -35.6813,
  -35.7127,
  -35.7443,
  -35.7765,
  -35.8094,
  -35.842,
  -35.8757,
  -35.9086,
  -35.9407,
  -35.9723,
  -36.0035,
  -36.0347,
  -36.0658,
  -36.0964,
  -36.1265,
  -36.1563,
  -36.186,
  -36.216,
  -36.2461,
  -36.2764,
  -36.3069,
  -36.3377,
  -36.3682,
  -36.3989,
  -36.4296,
  -36.4601,
  -36.4902,
  -36.5216,
  -36.5534,
  -36.5854,
  -36.6173,
  -36.6487,
  -36.6796,
  -36.7101,
  -36.7402,
  -36.7703,
  -36.8003,
  -36.8302,
  -36.8597,
  -36.8882,
  -36.9155,
  -36.9413,
  -36.9653,
  -36.9878,
  -37.0095,
  -37.031,
  -37.0529,
  -37.0758,
  -37.0988,
  -37.1241,
  -37.1504,
  -37.1774,
  -37.2047,
  -37.2313,
  -37.2568,
  -37.2808,
  -37.3031,
  -37.3241,
  -37.344,
  -37.3635,
  -37.3828,
  -37.4023,
  -37.422,
  -37.4417,
  -37.4616,
  -37.4812,
  -37.5006,
  -37.5199,
  -37.5389,
  -37.5577,
  -37.5766,
  -37.5956,
  -37.6145,
  -37.6321,
  -37.6504,
  -37.6681,
  -37.6853,
  -37.7021,
  -37.7186,
  -37.7356,
  -37.7538,
  -37.7737,
  -37.7955,
  -37.8187,
  -37.8431,
  -37.8683,
  -37.894,
  -37.9204,
  -37.9473,
  -37.9752,
  -38.0048,
  -38.0364,
  -38.0702,
  -38.1057,
  -38.1421,
  -38.1784,
  -38.2142,
  -38.2488,
  -38.2822,
  -38.3139,
  -38.3443,
  -38.3726,
  -38.4009,
  -38.4289,
  -38.457,
  -38.4854,
  -38.5146,
  -38.5451,
  -38.5765,
  -38.6088,
  -38.6416,
  -38.6741,
  -38.7062,
  -38.7374,
  -38.7674,
  -38.796,
  -38.8234,
  -38.8493,
  -38.874,
  -38.8976,
  -38.9202,
  -38.9409,
  -38.9608,
  -38.9794,
  -38.9977,
  -39.0156,
  -39.0332,
  -39.0503,
  -39.0668,
  -39.0828,
  -39.0982,
  -39.1129,
  -39.1266,
  -39.1393,
  -39.1502,
  -39.1615,
  -39.1722,
  -39.1822,
  -39.1913,
  -39.1995,
  -39.2067,
  -39.213,
  -39.2184,
  -39.2231,
  -39.2269,
  -39.23,
  -39.2324,
  -39.2344,
  -39.2359,
  -39.2369,
  -39.2372,
  -39.2364,
  -39.2341,
  -39.2297,
  -39.2234,
  -39.2149,
  -39.2046,
  -39.1927,
  -39.1795,
  -39.165,
  -39.1494,
  -39.1327,
  -39.1145,
  -39.0944,
  -39.0721,
  -39.047,
  -39.0188,
  -38.9876,
  -38.954,
  -38.9187,
  -38.8826,
  -38.8464,
  -38.81,
  -38.7728,
  -38.7328,
  -38.687,
  -38.6343,
  -38.572,
  -38.5,
  -38.4198,
  -38.3349,
  -38.2507,
  -38.1732,
  -38.1089,
  -38.063,
  -38.0378,
  -30.2507,
  -30.2979,
  -30.3457,
  -30.394,
  -30.4428,
  -30.4923,
  -30.5424,
  -30.5925,
  -30.6425,
  -30.6916,
  -30.7397,
  -30.7869,
  -30.8339,
  -30.8807,
  -30.9274,
  -30.9758,
  -31.0253,
  -31.076,
  -31.1277,
  -31.1801,
  -31.2322,
  -31.2833,
  -31.3329,
  -31.3809,
  -31.4273,
  -31.4725,
  -31.5175,
  -31.5628,
  -31.6094,
  -31.6565,
  -31.7061,
  -31.7569,
  -31.8086,
  -31.8611,
  -31.9138,
  -31.9665,
  -32.0189,
  -32.071,
  -32.1227,
  -32.1747,
  -32.2268,
  -32.2793,
  -32.3321,
  -32.3854,
  -32.4382,
  -32.4926,
  -32.5474,
  -32.6022,
  -32.6571,
  -32.7115,
  -32.7659,
  -32.82,
  -32.8738,
  -32.9272,
  -32.9801,
  -33.0323,
  -33.0841,
  -33.1356,
  -33.1875,
  -33.2397,
  -33.2912,
  -33.3436,
  -33.3959,
  -33.4479,
  -33.4994,
  -33.5504,
  -33.601,
  -33.6514,
  -33.7017,
  -33.752,
  -33.8026,
  -33.8532,
  -33.9041,
  -33.955,
  -34.0059,
  -34.0559,
  -34.1047,
  -34.1513,
  -34.1979,
  -34.2442,
  -34.2906,
  -34.3373,
  -34.3841,
  -34.4305,
  -34.4757,
  -34.5191,
  -34.5605,
  -34.6,
  -34.6384,
  -34.6766,
  -34.7154,
  -34.7552,
  -34.7962,
  -34.8379,
  -34.8798,
  -34.9206,
  -34.9617,
  -35.0019,
  -35.0413,
  -35.08,
  -35.1182,
  -35.156,
  -35.1931,
  -35.2295,
  -35.265,
  -35.3,
  -35.3345,
  -35.3688,
  -35.4027,
  -35.4362,
  -35.4691,
  -35.5015,
  -35.5332,
  -35.5648,
  -35.5954,
  -35.6271,
  -35.6588,
  -35.6907,
  -35.7234,
  -35.7567,
  -35.7906,
  -35.8242,
  -35.857,
  -35.8888,
  -35.9198,
  -35.9506,
  -35.9816,
  -36.0126,
  -36.0434,
  -36.0739,
  -36.104,
  -36.1341,
  -36.1642,
  -36.1943,
  -36.2237,
  -36.2542,
  -36.2848,
  -36.3158,
  -36.3467,
  -36.3779,
  -36.4091,
  -36.4409,
  -36.4732,
  -36.5059,
  -36.5384,
  -36.5704,
  -36.6016,
  -36.632,
  -36.6617,
  -36.6912,
  -36.7207,
  -36.7505,
  -36.7802,
  -36.8098,
  -36.8385,
  -36.8658,
  -36.8907,
  -36.9148,
  -36.9371,
  -36.9583,
  -36.9793,
  -37.0005,
  -37.0226,
  -37.0461,
  -37.0707,
  -37.0966,
  -37.1235,
  -37.1506,
  -37.1772,
  -37.2028,
  -37.2269,
  -37.2495,
  -37.2706,
  -37.2906,
  -37.31,
  -37.3292,
  -37.3486,
  -37.3683,
  -37.3882,
  -37.4081,
  -37.4267,
  -37.4461,
  -37.4653,
  -37.4843,
  -37.503,
  -37.5216,
  -37.54,
  -37.558,
  -37.5755,
  -37.5927,
  -37.6095,
  -37.6262,
  -37.6427,
  -37.6594,
  -37.6768,
  -37.6956,
  -37.7164,
  -37.7391,
  -37.7634,
  -37.7888,
  -37.8152,
  -37.8421,
  -37.8698,
  -37.8982,
  -37.9278,
  -37.959,
  -37.991,
  -38.026,
  -38.0624,
  -38.0995,
  -38.1369,
  -38.1733,
  -38.2086,
  -38.2425,
  -38.2747,
  -38.3054,
  -38.3348,
  -38.3635,
  -38.3918,
  -38.4203,
  -38.4493,
  -38.4789,
  -38.5095,
  -38.541,
  -38.5732,
  -38.6058,
  -38.6382,
  -38.6701,
  -38.7011,
  -38.731,
  -38.7595,
  -38.7867,
  -38.8127,
  -38.8377,
  -38.8618,
  -38.8848,
  -38.906,
  -38.9246,
  -38.9429,
  -38.9608,
  -38.9784,
  -38.9956,
  -39.0124,
  -39.0288,
  -39.0446,
  -39.0598,
  -39.0742,
  -39.0878,
  -39.1005,
  -39.1123,
  -39.1235,
  -39.1342,
  -39.1441,
  -39.1533,
  -39.1612,
  -39.1681,
  -39.1738,
  -39.1787,
  -39.1828,
  -39.1861,
  -39.1887,
  -39.1908,
  -39.1926,
  -39.1941,
  -39.1952,
  -39.1955,
  -39.1948,
  -39.1925,
  -39.1881,
  -39.1813,
  -39.1724,
  -39.1618,
  -39.1496,
  -39.1363,
  -39.1219,
  -39.1055,
  -39.0889,
  -39.0709,
  -39.0512,
  -39.0291,
  -39.0044,
  -38.9766,
  -38.946,
  -38.9131,
  -38.8785,
  -38.8431,
  -38.8073,
  -38.771,
  -38.7334,
  -38.6928,
  -38.6467,
  -38.5919,
  -38.5269,
  -38.4511,
  -38.3663,
  -38.2768,
  -38.1879,
  -38.1061,
  -38.0391,
  -37.9925,
  -37.9688,
  -30.1951,
  -30.242,
  -30.2898,
  -30.3383,
  -30.3874,
  -30.4372,
  -30.4876,
  -30.5382,
  -30.5886,
  -30.6372,
  -30.6859,
  -30.7339,
  -30.7816,
  -30.8294,
  -30.8775,
  -30.9263,
  -30.9761,
  -31.027,
  -31.079,
  -31.1316,
  -31.1839,
  -31.2353,
  -31.2851,
  -31.3332,
  -31.3789,
  -31.4246,
  -31.4701,
  -31.5162,
  -31.5638,
  -31.613,
  -31.6636,
  -31.7153,
  -31.7677,
  -31.8206,
  -31.8736,
  -31.9265,
  -31.9791,
  -32.0313,
  -32.0835,
  -32.1347,
  -32.1871,
  -32.2398,
  -32.2927,
  -32.3459,
  -32.3994,
  -32.4533,
  -32.5074,
  -32.5615,
  -32.6156,
  -32.6697,
  -32.7236,
  -32.7776,
  -32.8315,
  -32.8852,
  -32.9383,
  -32.9896,
  -33.0416,
  -33.0933,
  -33.145,
  -33.1967,
  -33.2482,
  -33.2994,
  -33.3502,
  -33.4009,
  -33.4513,
  -33.5014,
  -33.5513,
  -33.6012,
  -33.6512,
  -33.7012,
  -33.7516,
  -33.8021,
  -33.8518,
  -33.9026,
  -33.9531,
  -34.0027,
  -34.0511,
  -34.0984,
  -34.1448,
  -34.1909,
  -34.2371,
  -34.2838,
  -34.3306,
  -34.377,
  -34.4223,
  -34.4658,
  -34.5073,
  -34.547,
  -34.5856,
  -34.623,
  -34.6618,
  -34.7015,
  -34.7423,
  -34.7841,
  -34.8262,
  -34.8682,
  -34.9093,
  -34.9493,
  -34.9884,
  -35.0269,
  -35.0652,
  -35.1033,
  -35.1408,
  -35.1776,
  -35.2136,
  -35.2488,
  -35.2835,
  -35.3177,
  -35.3506,
  -35.3841,
  -35.4171,
  -35.4494,
  -35.4812,
  -35.5128,
  -35.5443,
  -35.5761,
  -35.6081,
  -35.6405,
  -35.6734,
  -35.707,
  -35.7408,
  -35.7743,
  -35.8068,
  -35.8381,
  -35.8687,
  -35.8992,
  -35.9298,
  -35.9596,
  -35.9904,
  -36.021,
  -36.0514,
  -36.0818,
  -36.1121,
  -36.1424,
  -36.1728,
  -36.2033,
  -36.2342,
  -36.2655,
  -36.2969,
  -36.3284,
  -36.3604,
  -36.3929,
  -36.4258,
  -36.4588,
  -36.4915,
  -36.5233,
  -36.5541,
  -36.5838,
  -36.6127,
  -36.6405,
  -36.6693,
  -36.6985,
  -36.728,
  -36.7574,
  -36.7864,
  -36.814,
  -36.8402,
  -36.8647,
  -36.8872,
  -36.9084,
  -36.929,
  -36.9498,
  -36.9713,
  -36.9941,
  -37.0182,
  -37.0437,
  -37.0702,
  -37.0971,
  -37.1236,
  -37.149,
  -37.1731,
  -37.1958,
  -37.2159,
  -37.2359,
  -37.2551,
  -37.2741,
  -37.2934,
  -37.3131,
  -37.3329,
  -37.3528,
  -37.3725,
  -37.3917,
  -37.4109,
  -37.43,
  -37.4488,
  -37.4674,
  -37.4853,
  -37.5027,
  -37.5194,
  -37.5356,
  -37.5517,
  -37.5678,
  -37.5841,
  -37.601,
  -37.619,
  -37.6387,
  -37.6604,
  -37.6841,
  -37.7083,
  -37.7346,
  -37.7617,
  -37.7895,
  -37.8182,
  -37.8481,
  -37.8792,
  -37.912,
  -37.9464,
  -37.9824,
  -38.0198,
  -38.0578,
  -38.0958,
  -38.1333,
  -38.1694,
  -38.2038,
  -38.2366,
  -38.2676,
  -38.2973,
  -38.3264,
  -38.3553,
  -38.3842,
  -38.4137,
  -38.4439,
  -38.4748,
  -38.5065,
  -38.5387,
  -38.5712,
  -38.6034,
  -38.6341,
  -38.6648,
  -38.6944,
  -38.7227,
  -38.7499,
  -38.7761,
  -38.8013,
  -38.8256,
  -38.8485,
  -38.8699,
  -38.8894,
  -38.9077,
  -38.9253,
  -38.9427,
  -38.9598,
  -38.9765,
  -38.9928,
  -39.0085,
  -39.0235,
  -39.0378,
  -39.0511,
  -39.0636,
  -39.0753,
  -39.0863,
  -39.0969,
  -39.1068,
  -39.1158,
  -39.1237,
  -39.1302,
  -39.1355,
  -39.14,
  -39.1436,
  -39.1463,
  -39.1484,
  -39.15,
  -39.1505,
  -39.1519,
  -39.153,
  -39.1535,
  -39.1529,
  -39.1506,
  -39.1461,
  -39.1391,
  -39.1298,
  -39.1187,
  -39.1063,
  -39.0929,
  -39.0786,
  -39.0634,
  -39.0471,
  -39.0296,
  -39.0103,
  -38.9889,
  -38.9648,
  -38.9378,
  -38.908,
  -38.8759,
  -38.8421,
  -38.8074,
  -38.7719,
  -38.7356,
  -38.6975,
  -38.6559,
  -38.6079,
  -38.5508,
  -38.4827,
  -38.4032,
  -38.3143,
  -38.2199,
  -38.1264,
  -38.0414,
  -37.972,
  -37.9245,
  -37.9019,
  -30.1417,
  -30.1885,
  -30.2362,
  -30.2847,
  -30.334,
  -30.383,
  -30.4335,
  -30.4843,
  -30.5349,
  -30.5849,
  -30.6341,
  -30.6828,
  -30.7315,
  -30.7803,
  -30.8292,
  -30.8787,
  -30.929,
  -30.9803,
  -31.0325,
  -31.0842,
  -31.1366,
  -31.188,
  -31.238,
  -31.2864,
  -31.3334,
  -31.3798,
  -31.426,
  -31.473,
  -31.5216,
  -31.5717,
  -31.6232,
  -31.6755,
  -31.7283,
  -31.7813,
  -31.8334,
  -31.8865,
  -31.9391,
  -31.9916,
  -32.0441,
  -32.0967,
  -32.1496,
  -32.2026,
  -32.2558,
  -32.309,
  -32.3621,
  -32.4154,
  -32.4687,
  -32.522,
  -32.5753,
  -32.6287,
  -32.6812,
  -32.7349,
  -32.7887,
  -32.8423,
  -32.8955,
  -32.9482,
  -33.0003,
  -33.052,
  -33.1034,
  -33.1545,
  -33.205,
  -33.2551,
  -33.3046,
  -33.3539,
  -33.4032,
  -33.4525,
  -33.5009,
  -33.5504,
  -33.6002,
  -33.6502,
  -33.7005,
  -33.751,
  -33.8017,
  -33.8522,
  -33.9024,
  -33.9519,
  -34,
  -34.047,
  -34.0933,
  -34.1395,
  -34.1858,
  -34.2323,
  -34.2792,
  -34.3256,
  -34.3698,
  -34.4134,
  -34.455,
  -34.495,
  -34.5338,
  -34.5723,
  -34.6112,
  -34.651,
  -34.6919,
  -34.7338,
  -34.7762,
  -34.8183,
  -34.8595,
  -34.8995,
  -34.9383,
  -34.9767,
  -35.015,
  -35.0532,
  -35.09,
  -35.1271,
  -35.1634,
  -35.1989,
  -35.2337,
  -35.268,
  -35.3019,
  -35.3354,
  -35.3684,
  -35.4008,
  -35.4327,
  -35.4644,
  -35.4961,
  -35.528,
  -35.5603,
  -35.5929,
  -35.626,
  -35.6595,
  -35.693,
  -35.7251,
  -35.7571,
  -35.788,
  -35.8182,
  -35.8484,
  -35.8786,
  -35.9092,
  -35.9398,
  -35.9705,
  -36.0011,
  -36.0317,
  -36.0623,
  -36.0929,
  -36.1235,
  -36.1542,
  -36.1853,
  -36.2167,
  -36.2485,
  -36.2806,
  -36.3132,
  -36.346,
  -36.378,
  -36.4109,
  -36.4434,
  -36.4749,
  -36.5051,
  -36.5342,
  -36.5625,
  -36.5905,
  -36.6186,
  -36.6471,
  -36.6761,
  -36.7053,
  -36.7342,
  -36.7624,
  -36.7892,
  -36.8141,
  -36.8372,
  -36.8587,
  -36.8794,
  -36.8999,
  -36.9209,
  -36.9432,
  -36.9658,
  -36.9908,
  -37.0168,
  -37.0433,
  -37.0695,
  -37.0946,
  -37.1186,
  -37.1412,
  -37.1622,
  -37.1821,
  -37.2011,
  -37.2198,
  -37.239,
  -37.2585,
  -37.2782,
  -37.2979,
  -37.3175,
  -37.3369,
  -37.3562,
  -37.3754,
  -37.3944,
  -37.4131,
  -37.4309,
  -37.4477,
  -37.4638,
  -37.4783,
  -37.4937,
  -37.5094,
  -37.5257,
  -37.5428,
  -37.5613,
  -37.5819,
  -37.6047,
  -37.6292,
  -37.6551,
  -37.6819,
  -37.7096,
  -37.7382,
  -37.7679,
  -37.7991,
  -37.8317,
  -37.8659,
  -37.9017,
  -37.9389,
  -37.9771,
  -38.0159,
  -38.0549,
  -38.093,
  -38.13,
  -38.1652,
  -38.1984,
  -38.23,
  -38.2603,
  -38.2888,
  -38.3183,
  -38.348,
  -38.378,
  -38.4087,
  -38.4401,
  -38.4721,
  -38.5043,
  -38.5366,
  -38.5687,
  -38.6001,
  -38.6305,
  -38.6598,
  -38.6879,
  -38.7149,
  -38.7411,
  -38.7663,
  -38.7906,
  -38.8134,
  -38.8346,
  -38.8541,
  -38.8724,
  -38.8901,
  -38.9075,
  -38.9247,
  -38.9414,
  -38.9576,
  -38.9731,
  -38.9878,
  -39.0018,
  -39.0151,
  -39.0274,
  -39.0388,
  -39.0486,
  -39.0589,
  -39.0686,
  -39.0775,
  -39.0853,
  -39.0917,
  -39.0967,
  -39.101,
  -39.1043,
  -39.1066,
  -39.1083,
  -39.1096,
  -39.1106,
  -39.1117,
  -39.1127,
  -39.1131,
  -39.1125,
  -39.1102,
  -39.1056,
  -39.0984,
  -39.0888,
  -39.0774,
  -39.0648,
  -39.0511,
  -39.0368,
  -39.0221,
  -39.0062,
  -38.9892,
  -38.9707,
  -38.9501,
  -38.9269,
  -38.9009,
  -38.872,
  -38.8407,
  -38.8078,
  -38.7736,
  -38.7384,
  -38.7018,
  -38.6629,
  -38.62,
  -38.5699,
  -38.5103,
  -38.4381,
  -38.3552,
  -38.2625,
  -38.1642,
  -38.067,
  -37.9791,
  -37.9082,
  -37.8602,
  -37.8384,
  -30.0902,
  -30.1368,
  -30.1843,
  -30.2327,
  -30.2819,
  -30.3319,
  -30.3824,
  -30.4331,
  -30.4836,
  -30.5337,
  -30.5835,
  -30.633,
  -30.6826,
  -30.7323,
  -30.7823,
  -30.8315,
  -30.8825,
  -30.9343,
  -30.9868,
  -31.0396,
  -31.0921,
  -31.1436,
  -31.1937,
  -31.2424,
  -31.29,
  -31.3369,
  -31.384,
  -31.432,
  -31.4813,
  -31.531,
  -31.5832,
  -31.6359,
  -31.6888,
  -31.7418,
  -31.7949,
  -31.848,
  -31.9009,
  -31.9536,
  -32.0064,
  -32.0594,
  -32.1128,
  -32.1662,
  -32.2197,
  -32.2728,
  -32.3257,
  -32.3772,
  -32.4297,
  -32.4822,
  -32.5348,
  -32.5876,
  -32.6405,
  -32.6936,
  -32.747,
  -32.8004,
  -32.8536,
  -32.9064,
  -32.9587,
  -33.0104,
  -33.0615,
  -33.1119,
  -33.1616,
  -33.2095,
  -33.2578,
  -33.306,
  -33.3543,
  -33.4029,
  -33.4518,
  -33.5012,
  -33.5509,
  -33.601,
  -33.6514,
  -33.702,
  -33.7526,
  -33.8031,
  -33.853,
  -33.9019,
  -33.95,
  -33.9969,
  -34.0424,
  -34.0891,
  -34.1355,
  -34.182,
  -34.2288,
  -34.275,
  -34.3204,
  -34.3639,
  -34.4058,
  -34.446,
  -34.4852,
  -34.5241,
  -34.5632,
  -34.6032,
  -34.6442,
  -34.6863,
  -34.7288,
  -34.7711,
  -34.8114,
  -34.8513,
  -34.89,
  -34.9282,
  -34.9663,
  -35.0046,
  -35.0425,
  -35.0798,
  -35.1164,
  -35.1521,
  -35.1872,
  -35.2216,
  -35.2555,
  -35.289,
  -35.322,
  -35.3545,
  -35.3867,
  -35.4186,
  -35.4506,
  -35.4817,
  -35.5143,
  -35.547,
  -35.5799,
  -35.613,
  -35.6461,
  -35.6785,
  -35.71,
  -35.7404,
  -35.7704,
  -35.8002,
  -35.8303,
  -35.8605,
  -35.8909,
  -35.9214,
  -35.9522,
  -35.9831,
  -36.014,
  -36.045,
  -36.0757,
  -36.1057,
  -36.137,
  -36.1686,
  -36.2006,
  -36.2329,
  -36.2656,
  -36.2985,
  -36.3314,
  -36.364,
  -36.3959,
  -36.4269,
  -36.4566,
  -36.4855,
  -36.5134,
  -36.5408,
  -36.5683,
  -36.5961,
  -36.6245,
  -36.6532,
  -36.682,
  -36.7103,
  -36.7376,
  -36.7622,
  -36.786,
  -36.8081,
  -36.8291,
  -36.8497,
  -36.8705,
  -36.8923,
  -36.9154,
  -36.9399,
  -36.9653,
  -36.9912,
  -37.0168,
  -37.0416,
  -37.0652,
  -37.0876,
  -37.1085,
  -37.1282,
  -37.1469,
  -37.1655,
  -37.1844,
  -37.2036,
  -37.2233,
  -37.2429,
  -37.2623,
  -37.2808,
  -37.3003,
  -37.3198,
  -37.339,
  -37.3577,
  -37.3754,
  -37.392,
  -37.4077,
  -37.4227,
  -37.4376,
  -37.4529,
  -37.469,
  -37.4861,
  -37.5054,
  -37.5271,
  -37.5506,
  -37.5759,
  -37.6024,
  -37.6296,
  -37.6577,
  -37.6871,
  -37.7178,
  -37.7502,
  -37.7844,
  -37.8202,
  -37.8574,
  -37.8957,
  -37.9339,
  -37.9735,
  -38.0131,
  -38.052,
  -38.0897,
  -38.1256,
  -38.1595,
  -38.1918,
  -38.2227,
  -38.2529,
  -38.2831,
  -38.3134,
  -38.3441,
  -38.3754,
  -38.4072,
  -38.4394,
  -38.4718,
  -38.5039,
  -38.5359,
  -38.5669,
  -38.597,
  -38.626,
  -38.6538,
  -38.6806,
  -38.7066,
  -38.7316,
  -38.7556,
  -38.7784,
  -38.7995,
  -38.819,
  -38.8374,
  -38.8543,
  -38.8719,
  -38.8892,
  -38.906,
  -38.922,
  -38.9372,
  -38.9514,
  -38.9652,
  -38.9781,
  -38.9902,
  -39.0013,
  -39.0118,
  -39.0218,
  -39.0312,
  -39.0399,
  -39.0475,
  -39.0539,
  -39.0592,
  -39.0632,
  -39.0664,
  -39.0688,
  -39.0704,
  -39.0715,
  -39.0723,
  -39.073,
  -39.0735,
  -39.0737,
  -39.0729,
  -39.0704,
  -39.0657,
  -39.0584,
  -39.0486,
  -39.0369,
  -39.0239,
  -39.0102,
  -38.996,
  -38.9813,
  -38.9659,
  -38.9487,
  -38.931,
  -38.9113,
  -38.8891,
  -38.864,
  -38.836,
  -38.8056,
  -38.7735,
  -38.7399,
  -38.7047,
  -38.6677,
  -38.6278,
  -38.5832,
  -38.5313,
  -38.4691,
  -38.3954,
  -38.3095,
  -38.2136,
  -38.1124,
  -38.0129,
  -37.923,
  -37.8509,
  -37.8028,
  -37.7815,
  -30.0429,
  -30.0892,
  -30.1364,
  -30.1845,
  -30.2335,
  -30.2832,
  -30.3335,
  -30.384,
  -30.4344,
  -30.4845,
  -30.5335,
  -30.5836,
  -30.6338,
  -30.6844,
  -30.7354,
  -30.7865,
  -30.8382,
  -30.8906,
  -30.9434,
  -30.9963,
  -31.0488,
  -31.1005,
  -31.1509,
  -31.2001,
  -31.2483,
  -31.295,
  -31.3428,
  -31.3915,
  -31.4413,
  -31.4924,
  -31.5446,
  -31.5974,
  -31.6504,
  -31.7035,
  -31.7565,
  -31.8094,
  -31.8623,
  -31.9153,
  -31.9687,
  -32.0224,
  -32.0754,
  -32.1294,
  -32.183,
  -32.2361,
  -32.2885,
  -32.3404,
  -32.3922,
  -32.444,
  -32.4959,
  -32.5481,
  -32.6005,
  -32.653,
  -32.7056,
  -32.7585,
  -32.8114,
  -32.8642,
  -32.9156,
  -32.9673,
  -33.0181,
  -33.0679,
  -33.1166,
  -33.1645,
  -33.2119,
  -33.2592,
  -33.3067,
  -33.3547,
  -33.4034,
  -33.4528,
  -33.5027,
  -33.5529,
  -33.6035,
  -33.6541,
  -33.7037,
  -33.754,
  -33.8038,
  -33.8526,
  -33.9007,
  -33.9477,
  -33.9944,
  -34.0412,
  -34.0877,
  -34.1346,
  -34.1814,
  -34.2277,
  -34.2727,
  -34.3164,
  -34.3585,
  -34.3992,
  -34.439,
  -34.4784,
  -34.5169,
  -34.5571,
  -34.5983,
  -34.6404,
  -34.683,
  -34.7252,
  -34.7664,
  -34.8063,
  -34.845,
  -34.8832,
  -34.9214,
  -34.9595,
  -34.9974,
  -35.0348,
  -35.0715,
  -35.1075,
  -35.1427,
  -35.1773,
  -35.2113,
  -35.2438,
  -35.2768,
  -35.3095,
  -35.3419,
  -35.3743,
  -35.4067,
  -35.4392,
  -35.4718,
  -35.5043,
  -35.5369,
  -35.5696,
  -35.602,
  -35.6337,
  -35.6644,
  -35.6945,
  -35.7242,
  -35.7539,
  -35.7836,
  -35.8134,
  -35.8425,
  -35.8729,
  -35.9038,
  -35.935,
  -35.9663,
  -35.9976,
  -36.0286,
  -36.0597,
  -36.091,
  -36.1224,
  -36.1544,
  -36.1868,
  -36.2194,
  -36.2521,
  -36.2846,
  -36.3166,
  -36.3479,
  -36.3785,
  -36.4081,
  -36.4368,
  -36.4647,
  -36.4919,
  -36.518,
  -36.5452,
  -36.5728,
  -36.6009,
  -36.6292,
  -36.6575,
  -36.6851,
  -36.7113,
  -36.7358,
  -36.7586,
  -36.7801,
  -36.8009,
  -36.8217,
  -36.8433,
  -36.8659,
  -36.8897,
  -36.9144,
  -36.9395,
  -36.9644,
  -36.9888,
  -37.0121,
  -37.0341,
  -37.0548,
  -37.0732,
  -37.0917,
  -37.11,
  -37.1286,
  -37.1476,
  -37.1668,
  -37.1862,
  -37.2056,
  -37.2251,
  -37.2448,
  -37.2646,
  -37.284,
  -37.3027,
  -37.3205,
  -37.3371,
  -37.3525,
  -37.3672,
  -37.3817,
  -37.3967,
  -37.4127,
  -37.4304,
  -37.4504,
  -37.4724,
  -37.4966,
  -37.5225,
  -37.5493,
  -37.5761,
  -37.6049,
  -37.635,
  -37.667,
  -37.7009,
  -37.7367,
  -37.7741,
  -37.8128,
  -37.8523,
  -37.8924,
  -37.933,
  -37.9732,
  -38.0129,
  -38.0511,
  -38.0876,
  -38.1222,
  -38.1552,
  -38.187,
  -38.218,
  -38.2487,
  -38.2796,
  -38.311,
  -38.3428,
  -38.375,
  -38.4073,
  -38.4397,
  -38.4718,
  -38.5035,
  -38.5344,
  -38.563,
  -38.5916,
  -38.6191,
  -38.6455,
  -38.6711,
  -38.6958,
  -38.7196,
  -38.7426,
  -38.7634,
  -38.7831,
  -38.8019,
  -38.8201,
  -38.8379,
  -38.8554,
  -38.872,
  -38.8877,
  -38.9024,
  -38.9163,
  -38.9296,
  -38.9422,
  -38.9539,
  -38.9647,
  -38.9748,
  -38.9844,
  -38.9935,
  -39.002,
  -39.0097,
  -39.0163,
  -39.0217,
  -39.026,
  -39.0294,
  -39.0319,
  -39.0336,
  -39.0347,
  -39.0354,
  -39.0358,
  -39.0349,
  -39.0344,
  -39.0331,
  -39.0303,
  -39.0255,
  -39.0182,
  -39.0084,
  -38.9965,
  -38.9833,
  -38.9694,
  -38.9551,
  -38.9405,
  -38.9256,
  -38.91,
  -38.8931,
  -38.8742,
  -38.8527,
  -38.8285,
  -38.8014,
  -38.7719,
  -38.7406,
  -38.7073,
  -38.6722,
  -38.6347,
  -38.5938,
  -38.5477,
  -38.4938,
  -38.4294,
  -38.3534,
  -38.2652,
  -38.1671,
  -38.064,
  -37.963,
  -37.8724,
  -37.8001,
  -37.7522,
  -37.731,
  -29.9986,
  -30.0447,
  -30.0916,
  -30.1393,
  -30.1878,
  -30.2361,
  -30.2861,
  -30.3363,
  -30.3865,
  -30.4367,
  -30.4868,
  -30.5372,
  -30.588,
  -30.6393,
  -30.691,
  -30.7431,
  -30.7955,
  -30.8482,
  -30.9013,
  -30.9544,
  -31.0061,
  -31.0579,
  -31.1086,
  -31.1583,
  -31.2072,
  -31.2556,
  -31.3042,
  -31.3535,
  -31.4037,
  -31.4551,
  -31.5072,
  -31.56,
  -31.6129,
  -31.6657,
  -31.7188,
  -31.7706,
  -31.8235,
  -31.8769,
  -31.9307,
  -31.9848,
  -32.0391,
  -32.0934,
  -32.1471,
  -32.1999,
  -32.2518,
  -32.3032,
  -32.3544,
  -32.4058,
  -32.4574,
  -32.5091,
  -32.561,
  -32.6118,
  -32.6637,
  -32.716,
  -32.7685,
  -32.821,
  -32.8732,
  -32.9247,
  -32.9751,
  -33.0243,
  -33.0723,
  -33.1194,
  -33.1662,
  -33.2129,
  -33.2598,
  -33.3074,
  -33.3559,
  -33.4042,
  -33.4543,
  -33.5048,
  -33.5555,
  -33.6062,
  -33.6569,
  -33.7073,
  -33.7571,
  -33.8061,
  -33.8541,
  -33.9015,
  -33.9484,
  -33.9953,
  -34.0422,
  -34.0892,
  -34.1362,
  -34.1823,
  -34.2264,
  -34.2701,
  -34.3124,
  -34.3536,
  -34.3936,
  -34.4335,
  -34.4734,
  -34.514,
  -34.5555,
  -34.5978,
  -34.6402,
  -34.6823,
  -34.7233,
  -34.7631,
  -34.802,
  -34.8404,
  -34.8785,
  -34.9167,
  -34.9536,
  -34.991,
  -35.0278,
  -35.064,
  -35.0995,
  -35.1342,
  -35.1683,
  -35.2019,
  -35.235,
  -35.2677,
  -35.3003,
  -35.3329,
  -35.3655,
  -35.3983,
  -35.4308,
  -35.4632,
  -35.4954,
  -35.5275,
  -35.5592,
  -35.5903,
  -35.6196,
  -35.6493,
  -35.6786,
  -35.7079,
  -35.7373,
  -35.7667,
  -35.7964,
  -35.8267,
  -35.8576,
  -35.8891,
  -35.9206,
  -35.9521,
  -35.9833,
  -36.0145,
  -36.0455,
  -36.0768,
  -36.1086,
  -36.1407,
  -36.1731,
  -36.2055,
  -36.2376,
  -36.2682,
  -36.2992,
  -36.3295,
  -36.359,
  -36.3879,
  -36.4158,
  -36.443,
  -36.4698,
  -36.4964,
  -36.5234,
  -36.5508,
  -36.5786,
  -36.6065,
  -36.6339,
  -36.6604,
  -36.6853,
  -36.7088,
  -36.7309,
  -36.7521,
  -36.7732,
  -36.7947,
  -36.8169,
  -36.8389,
  -36.8627,
  -36.8868,
  -36.9109,
  -36.9346,
  -36.9574,
  -36.9791,
  -36.9995,
  -37.0187,
  -37.0371,
  -37.0553,
  -37.0738,
  -37.0926,
  -37.1118,
  -37.1312,
  -37.1506,
  -37.1701,
  -37.1897,
  -37.2093,
  -37.2286,
  -37.2472,
  -37.2649,
  -37.2813,
  -37.2967,
  -37.3113,
  -37.3248,
  -37.3399,
  -37.3563,
  -37.3744,
  -37.3947,
  -37.4172,
  -37.4419,
  -37.4681,
  -37.4954,
  -37.5237,
  -37.5533,
  -37.5846,
  -37.6178,
  -37.6533,
  -37.6908,
  -37.7299,
  -37.7702,
  -37.8111,
  -37.8524,
  -37.8937,
  -37.9346,
  -37.9744,
  -38.013,
  -38.0498,
  -38.0851,
  -38.1187,
  -38.1516,
  -38.1833,
  -38.2138,
  -38.2455,
  -38.2773,
  -38.3095,
  -38.3419,
  -38.3743,
  -38.4066,
  -38.4387,
  -38.4701,
  -38.5007,
  -38.53,
  -38.5583,
  -38.5855,
  -38.6116,
  -38.6369,
  -38.6616,
  -38.6853,
  -38.708,
  -38.7291,
  -38.7491,
  -38.7682,
  -38.7868,
  -38.8048,
  -38.8222,
  -38.8387,
  -38.854,
  -38.8682,
  -38.8817,
  -38.8944,
  -38.9063,
  -38.9175,
  -38.9278,
  -38.9375,
  -38.9456,
  -38.9544,
  -38.9629,
  -38.9706,
  -38.9775,
  -38.9833,
  -38.9881,
  -38.9919,
  -38.9949,
  -38.997,
  -38.9984,
  -38.9992,
  -38.9993,
  -38.9989,
  -38.9979,
  -38.9959,
  -38.9927,
  -38.9877,
  -38.9803,
  -38.9705,
  -38.9587,
  -38.9454,
  -38.9313,
  -38.9168,
  -38.9023,
  -38.8874,
  -38.8721,
  -38.8558,
  -38.8375,
  -38.8167,
  -38.7933,
  -38.7673,
  -38.7386,
  -38.708,
  -38.675,
  -38.6397,
  -38.6015,
  -38.5592,
  -38.5114,
  -38.4556,
  -38.3895,
  -38.3115,
  -38.2215,
  -38.121,
  -38.0172,
  -37.9159,
  -37.8253,
  -37.7537,
  -37.7062,
  -37.6851,
  -29.9571,
  -30.0021,
  -30.0486,
  -30.0959,
  -30.144,
  -30.1929,
  -30.2424,
  -30.2924,
  -30.3422,
  -30.3922,
  -30.4424,
  -30.4929,
  -30.544,
  -30.5958,
  -30.6482,
  -30.6999,
  -30.753,
  -30.8064,
  -30.8596,
  -30.9126,
  -30.9654,
  -31.0172,
  -31.0684,
  -31.1188,
  -31.1684,
  -31.2176,
  -31.2668,
  -31.3165,
  -31.3669,
  -31.4182,
  -31.4691,
  -31.5216,
  -31.5744,
  -31.6272,
  -31.6801,
  -31.733,
  -31.7863,
  -31.8399,
  -31.894,
  -31.9485,
  -32.003,
  -32.0572,
  -32.1107,
  -32.1632,
  -32.2146,
  -32.2656,
  -32.3156,
  -32.3669,
  -32.4184,
  -32.4699,
  -32.5214,
  -32.5726,
  -32.6237,
  -32.6752,
  -32.727,
  -32.779,
  -32.8308,
  -32.8819,
  -32.9318,
  -32.9802,
  -33.0278,
  -33.0745,
  -33.12,
  -33.1664,
  -33.2131,
  -33.2604,
  -33.3087,
  -33.3581,
  -33.4082,
  -33.4588,
  -33.5097,
  -33.5606,
  -33.6115,
  -33.6621,
  -33.712,
  -33.761,
  -33.809,
  -33.8564,
  -33.9036,
  -33.9497,
  -33.997,
  -34.0444,
  -34.0914,
  -34.1377,
  -34.183,
  -34.2268,
  -34.2694,
  -34.3107,
  -34.3511,
  -34.3914,
  -34.4318,
  -34.4728,
  -34.5145,
  -34.557,
  -34.5993,
  -34.6409,
  -34.6818,
  -34.7207,
  -34.76,
  -34.7985,
  -34.8369,
  -34.8751,
  -34.9132,
  -34.9506,
  -34.9875,
  -35.0237,
  -35.0593,
  -35.0943,
  -35.1286,
  -35.1622,
  -35.1952,
  -35.228,
  -35.2607,
  -35.2934,
  -35.3262,
  -35.3589,
  -35.3903,
  -35.4223,
  -35.454,
  -35.4854,
  -35.5165,
  -35.5471,
  -35.577,
  -35.6063,
  -35.6354,
  -35.6643,
  -35.6933,
  -35.7223,
  -35.7517,
  -35.7818,
  -35.8126,
  -35.844,
  -35.8757,
  -35.9073,
  -35.9386,
  -35.9696,
  -35.9994,
  -36.0303,
  -36.0617,
  -36.0935,
  -36.1255,
  -36.1575,
  -36.1893,
  -36.2206,
  -36.2515,
  -36.2818,
  -36.3116,
  -36.3407,
  -36.3689,
  -36.3963,
  -36.4231,
  -36.4495,
  -36.4759,
  -36.5025,
  -36.5295,
  -36.5565,
  -36.5835,
  -36.6097,
  -36.6338,
  -36.6577,
  -36.6805,
  -36.7024,
  -36.7237,
  -36.7451,
  -36.7667,
  -36.7888,
  -36.8116,
  -36.8347,
  -36.8579,
  -36.8809,
  -36.9033,
  -36.9246,
  -36.9448,
  -36.9639,
  -36.9823,
  -37.0005,
  -37.019,
  -37.0378,
  -37.057,
  -37.0764,
  -37.0959,
  -37.1153,
  -37.1337,
  -37.1528,
  -37.1716,
  -37.1899,
  -37.2073,
  -37.2236,
  -37.239,
  -37.2538,
  -37.2687,
  -37.2843,
  -37.3011,
  -37.3196,
  -37.3403,
  -37.363,
  -37.3878,
  -37.4142,
  -37.4419,
  -37.4711,
  -37.5018,
  -37.5345,
  -37.5693,
  -37.6065,
  -37.646,
  -37.687,
  -37.729,
  -37.7714,
  -37.8138,
  -37.8551,
  -37.8964,
  -37.9363,
  -37.9749,
  -38.0119,
  -38.0476,
  -38.0822,
  -38.1157,
  -38.1485,
  -38.1807,
  -38.2129,
  -38.2452,
  -38.2777,
  -38.3102,
  -38.3426,
  -38.3747,
  -38.4064,
  -38.4374,
  -38.4676,
  -38.4968,
  -38.5248,
  -38.5517,
  -38.5778,
  -38.6029,
  -38.6273,
  -38.6508,
  -38.6737,
  -38.6952,
  -38.7157,
  -38.7352,
  -38.7541,
  -38.7713,
  -38.7888,
  -38.805,
  -38.82,
  -38.8337,
  -38.8464,
  -38.8584,
  -38.8696,
  -38.8801,
  -38.8898,
  -38.899,
  -38.9077,
  -38.9164,
  -38.925,
  -38.9329,
  -38.9404,
  -38.9467,
  -38.952,
  -38.9564,
  -38.96,
  -38.9626,
  -38.9644,
  -38.9653,
  -38.9653,
  -38.9644,
  -38.9627,
  -38.96,
  -38.9564,
  -38.951,
  -38.9437,
  -38.934,
  -38.9223,
  -38.9089,
  -38.8946,
  -38.8799,
  -38.8651,
  -38.8502,
  -38.835,
  -38.819,
  -38.8001,
  -38.7801,
  -38.7576,
  -38.7324,
  -38.7046,
  -38.6745,
  -38.6418,
  -38.6062,
  -38.5672,
  -38.5237,
  -38.4741,
  -38.4164,
  -38.3484,
  -38.2686,
  -38.1772,
  -38.0769,
  -37.9724,
  -37.8712,
  -37.7822,
  -37.7118,
  -37.6652,
  -37.6442,
  -29.9171,
  -29.9632,
  -30.0094,
  -30.0562,
  -30.1039,
  -30.1522,
  -30.2014,
  -30.2508,
  -30.3004,
  -30.3502,
  -30.4003,
  -30.45,
  -30.5013,
  -30.5535,
  -30.6065,
  -30.6599,
  -30.7136,
  -30.7672,
  -30.8206,
  -30.8737,
  -30.9262,
  -30.9782,
  -31.0298,
  -31.0807,
  -31.1309,
  -31.1797,
  -31.2294,
  -31.2795,
  -31.33,
  -31.3812,
  -31.4331,
  -31.4855,
  -31.5382,
  -31.5909,
  -31.6437,
  -31.6967,
  -31.7501,
  -31.804,
  -31.8582,
  -31.9125,
  -31.9667,
  -32.0196,
  -32.0727,
  -32.1247,
  -32.176,
  -32.2268,
  -32.2778,
  -32.3292,
  -32.3809,
  -32.4325,
  -32.4837,
  -32.5344,
  -32.5848,
  -32.6354,
  -32.6864,
  -32.7378,
  -32.789,
  -32.8385,
  -32.8876,
  -32.9356,
  -32.9827,
  -33.0292,
  -33.0758,
  -33.1222,
  -33.169,
  -33.2163,
  -33.2644,
  -33.3136,
  -33.3637,
  -33.4142,
  -33.4652,
  -33.5162,
  -33.5673,
  -33.6172,
  -33.6674,
  -33.7165,
  -33.7647,
  -33.8121,
  -33.8595,
  -33.9068,
  -33.9545,
  -34.0021,
  -34.0494,
  -34.0958,
  -34.1411,
  -34.1852,
  -34.2279,
  -34.2694,
  -34.3104,
  -34.3509,
  -34.3916,
  -34.4319,
  -34.4741,
  -34.5164,
  -34.5588,
  -34.6007,
  -34.6416,
  -34.6814,
  -34.7209,
  -34.7597,
  -34.7983,
  -34.8366,
  -34.8747,
  -34.9121,
  -34.9488,
  -34.9851,
  -35.0209,
  -35.0561,
  -35.0905,
  -35.1231,
  -35.1562,
  -35.189,
  -35.2217,
  -35.2544,
  -35.2871,
  -35.3195,
  -35.3514,
  -35.3828,
  -35.4139,
  -35.4447,
  -35.4754,
  -35.5056,
  -35.5351,
  -35.5641,
  -35.5928,
  -35.6214,
  -35.6501,
  -35.6788,
  -35.708,
  -35.7367,
  -35.7672,
  -35.7984,
  -35.8299,
  -35.8613,
  -35.8924,
  -35.9233,
  -35.9538,
  -35.9844,
  -36.0153,
  -36.0466,
  -36.0783,
  -36.11,
  -36.1416,
  -36.1729,
  -36.2039,
  -36.2345,
  -36.2647,
  -36.2943,
  -36.3229,
  -36.3507,
  -36.3775,
  -36.4028,
  -36.4287,
  -36.4546,
  -36.4805,
  -36.5068,
  -36.5327,
  -36.5585,
  -36.5835,
  -36.6076,
  -36.6308,
  -36.6531,
  -36.6747,
  -36.6958,
  -36.7168,
  -36.7379,
  -36.7596,
  -36.7818,
  -36.8043,
  -36.8267,
  -36.8486,
  -36.8697,
  -36.8897,
  -36.9088,
  -36.9262,
  -36.9447,
  -36.9632,
  -36.9822,
  -37.0016,
  -37.021,
  -37.0404,
  -37.0599,
  -37.0787,
  -37.0972,
  -37.1153,
  -37.133,
  -37.15,
  -37.1663,
  -37.1817,
  -37.1968,
  -37.2123,
  -37.2285,
  -37.246,
  -37.2651,
  -37.286,
  -37.3089,
  -37.3337,
  -37.3604,
  -37.3887,
  -37.4187,
  -37.4496,
  -37.484,
  -37.5203,
  -37.5596,
  -37.6009,
  -37.6437,
  -37.6873,
  -37.7313,
  -37.775,
  -37.818,
  -37.8598,
  -37.8999,
  -37.9384,
  -37.9757,
  -38.0117,
  -38.0468,
  -38.0811,
  -38.1146,
  -38.1476,
  -38.1805,
  -38.2132,
  -38.246,
  -38.2784,
  -38.3103,
  -38.342,
  -38.3731,
  -38.4037,
  -38.4336,
  -38.4626,
  -38.4906,
  -38.5167,
  -38.5428,
  -38.5679,
  -38.5922,
  -38.616,
  -38.6389,
  -38.6609,
  -38.6819,
  -38.702,
  -38.7213,
  -38.7398,
  -38.7572,
  -38.7731,
  -38.7876,
  -38.8006,
  -38.8125,
  -38.8236,
  -38.834,
  -38.8438,
  -38.8528,
  -38.8616,
  -38.8702,
  -38.8787,
  -38.8872,
  -38.8957,
  -38.9037,
  -38.9108,
  -38.9168,
  -38.9219,
  -38.9261,
  -38.9293,
  -38.9314,
  -38.9323,
  -38.932,
  -38.9307,
  -38.9275,
  -38.9242,
  -38.9199,
  -38.9142,
  -38.9069,
  -38.8974,
  -38.8859,
  -38.8724,
  -38.8579,
  -38.8428,
  -38.8276,
  -38.8126,
  -38.7974,
  -38.7815,
  -38.7643,
  -38.7452,
  -38.7235,
  -38.6993,
  -38.6722,
  -38.6425,
  -38.6097,
  -38.5737,
  -38.5337,
  -38.4887,
  -38.4375,
  -38.3779,
  -38.3081,
  -38.2267,
  -38.1337,
  -38.0326,
  -37.9283,
  -37.8283,
  -37.7404,
  -37.6713,
  -37.6258,
  -37.6048,
  -29.8809,
  -29.9266,
  -29.9726,
  -30.019,
  -30.066,
  -30.1138,
  -30.1613,
  -30.2102,
  -30.2594,
  -30.3091,
  -30.3593,
  -30.4103,
  -30.462,
  -30.5148,
  -30.5683,
  -30.6224,
  -30.6765,
  -30.7304,
  -30.7838,
  -30.8367,
  -30.8891,
  -30.9402,
  -30.9919,
  -31.0431,
  -31.0937,
  -31.144,
  -31.1941,
  -31.2445,
  -31.2953,
  -31.3466,
  -31.3984,
  -31.4507,
  -31.5033,
  -31.5559,
  -31.6086,
  -31.6616,
  -31.7141,
  -31.7679,
  -31.822,
  -31.8758,
  -31.9294,
  -31.9828,
  -32.0353,
  -32.087,
  -32.1381,
  -32.189,
  -32.2402,
  -32.2918,
  -32.3437,
  -32.3954,
  -32.4465,
  -32.4959,
  -32.5459,
  -32.5959,
  -32.6461,
  -32.6966,
  -32.747,
  -32.7966,
  -32.8451,
  -32.8926,
  -32.9394,
  -32.9862,
  -33.033,
  -33.0798,
  -33.1268,
  -33.1741,
  -33.2222,
  -33.2711,
  -33.3198,
  -33.3703,
  -33.421,
  -33.4722,
  -33.5235,
  -33.5746,
  -33.6251,
  -33.6745,
  -33.7229,
  -33.7705,
  -33.8181,
  -33.8657,
  -33.9137,
  -33.9615,
  -34.009,
  -34.0554,
  -34.1008,
  -34.1437,
  -34.1864,
  -34.2283,
  -34.2696,
  -34.3105,
  -34.3516,
  -34.3932,
  -34.4357,
  -34.4784,
  -34.5211,
  -34.5632,
  -34.6044,
  -34.6444,
  -34.6839,
  -34.7228,
  -34.7613,
  -34.7996,
  -34.8376,
  -34.874,
  -34.9109,
  -34.9472,
  -34.983,
  -35.0182,
  -35.0526,
  -35.0863,
  -35.1194,
  -35.1523,
  -35.1851,
  -35.2176,
  -35.2499,
  -35.2818,
  -35.3131,
  -35.3437,
  -35.3742,
  -35.4045,
  -35.4347,
  -35.4645,
  -35.4937,
  -35.5213,
  -35.5496,
  -35.578,
  -35.6063,
  -35.6348,
  -35.6637,
  -35.6931,
  -35.7232,
  -35.7538,
  -35.7847,
  -35.8158,
  -35.8468,
  -35.8773,
  -35.9075,
  -35.9376,
  -35.9681,
  -35.999,
  -36.0303,
  -36.0619,
  -36.0935,
  -36.1249,
  -36.1551,
  -36.1862,
  -36.2169,
  -36.2469,
  -36.2761,
  -36.3042,
  -36.3313,
  -36.3574,
  -36.3829,
  -36.4082,
  -36.4333,
  -36.4585,
  -36.4838,
  -36.5088,
  -36.5335,
  -36.5575,
  -36.5809,
  -36.6033,
  -36.6248,
  -36.6456,
  -36.6659,
  -36.6862,
  -36.7058,
  -36.7272,
  -36.749,
  -36.7709,
  -36.7926,
  -36.8135,
  -36.8334,
  -36.8525,
  -36.8711,
  -36.8897,
  -36.9085,
  -36.9277,
  -36.9472,
  -36.967,
  -36.9864,
  -37.0056,
  -37.0239,
  -37.0415,
  -37.0589,
  -37.0761,
  -37.0927,
  -37.1088,
  -37.1244,
  -37.1398,
  -37.1559,
  -37.1718,
  -37.19,
  -37.2097,
  -37.2311,
  -37.2542,
  -37.2792,
  -37.306,
  -37.3349,
  -37.3658,
  -37.3991,
  -37.4347,
  -37.4732,
  -37.514,
  -37.557,
  -37.6016,
  -37.647,
  -37.6925,
  -37.7375,
  -37.7813,
  -37.8234,
  -37.8638,
  -37.9024,
  -37.9396,
  -37.9758,
  -38.0115,
  -38.0464,
  -38.0807,
  -38.1145,
  -38.148,
  -38.1801,
  -38.213,
  -38.2452,
  -38.2768,
  -38.3078,
  -38.3383,
  -38.3682,
  -38.3976,
  -38.4264,
  -38.4546,
  -38.482,
  -38.5084,
  -38.5338,
  -38.5583,
  -38.582,
  -38.6052,
  -38.6275,
  -38.6493,
  -38.67,
  -38.6898,
  -38.7087,
  -38.7259,
  -38.7415,
  -38.7555,
  -38.7678,
  -38.7788,
  -38.7892,
  -38.7987,
  -38.8077,
  -38.8163,
  -38.8247,
  -38.8331,
  -38.8415,
  -38.8493,
  -38.8583,
  -38.8667,
  -38.8744,
  -38.8812,
  -38.887,
  -38.8918,
  -38.8954,
  -38.8976,
  -38.8984,
  -38.8978,
  -38.8961,
  -38.8931,
  -38.889,
  -38.8842,
  -38.8785,
  -38.8713,
  -38.8622,
  -38.8509,
  -38.8377,
  -38.8229,
  -38.8074,
  -38.7919,
  -38.7766,
  -38.7614,
  -38.7458,
  -38.7292,
  -38.7109,
  -38.6903,
  -38.6669,
  -38.6404,
  -38.6108,
  -38.5777,
  -38.5411,
  -38.5001,
  -38.4537,
  -38.4009,
  -38.3394,
  -38.2676,
  -38.1845,
  -38.0903,
  -37.9883,
  -37.884,
  -37.7834,
  -37.6967,
  -37.6293,
  -37.5843,
  -37.563,
  -29.8466,
  -29.892,
  -29.9366,
  -29.9825,
  -30.029,
  -30.0762,
  -30.124,
  -30.1724,
  -30.2214,
  -30.271,
  -30.3213,
  -30.3727,
  -30.4252,
  -30.4785,
  -30.5327,
  -30.5873,
  -30.6408,
  -30.6949,
  -30.7481,
  -30.8007,
  -30.853,
  -30.9051,
  -30.9569,
  -31.0082,
  -31.0592,
  -31.1099,
  -31.1605,
  -31.2112,
  -31.2621,
  -31.3134,
  -31.3652,
  -31.4165,
  -31.469,
  -31.5215,
  -31.5739,
  -31.6267,
  -31.6802,
  -31.7337,
  -31.7872,
  -31.8405,
  -31.8934,
  -31.9458,
  -31.9978,
  -32.049,
  -32.1001,
  -32.1512,
  -32.2017,
  -32.2537,
  -32.3057,
  -32.3574,
  -32.4085,
  -32.4587,
  -32.5085,
  -32.558,
  -32.6075,
  -32.6572,
  -32.7066,
  -32.7552,
  -32.803,
  -32.8503,
  -32.8973,
  -32.9444,
  -32.9908,
  -33.0381,
  -33.0856,
  -33.133,
  -33.1809,
  -33.2294,
  -33.2787,
  -33.3288,
  -33.3794,
  -33.4305,
  -33.482,
  -33.5335,
  -33.5843,
  -33.6341,
  -33.6829,
  -33.7309,
  -33.7786,
  -33.8256,
  -33.8738,
  -33.9218,
  -33.9692,
  -34.0157,
  -34.061,
  -34.1048,
  -34.1475,
  -34.1894,
  -34.2309,
  -34.2722,
  -34.3137,
  -34.3555,
  -34.3982,
  -34.4415,
  -34.4846,
  -34.5272,
  -34.5688,
  -34.6082,
  -34.6477,
  -34.6865,
  -34.7249,
  -34.7631,
  -34.8009,
  -34.8383,
  -34.8753,
  -34.9116,
  -34.9474,
  -34.9824,
  -35.0168,
  -35.0503,
  -35.0835,
  -35.1166,
  -35.1493,
  -35.1817,
  -35.2135,
  -35.2447,
  -35.2742,
  -35.3043,
  -35.3341,
  -35.364,
  -35.3937,
  -35.4229,
  -35.4516,
  -35.4798,
  -35.5078,
  -35.5357,
  -35.5636,
  -35.5918,
  -35.6202,
  -35.6492,
  -35.6788,
  -35.709,
  -35.7394,
  -35.77,
  -35.8003,
  -35.8304,
  -35.8603,
  -35.8891,
  -35.9192,
  -35.9498,
  -35.9809,
  -36.0123,
  -36.0439,
  -36.0756,
  -36.107,
  -36.1385,
  -36.1695,
  -36.2,
  -36.2295,
  -36.2579,
  -36.2851,
  -36.3112,
  -36.3365,
  -36.3614,
  -36.386,
  -36.4105,
  -36.435,
  -36.4594,
  -36.4835,
  -36.5063,
  -36.5296,
  -36.5519,
  -36.5732,
  -36.5933,
  -36.6128,
  -36.6321,
  -36.652,
  -36.6725,
  -36.694,
  -36.7158,
  -36.7372,
  -36.7581,
  -36.7781,
  -36.7973,
  -36.8161,
  -36.8349,
  -36.8539,
  -36.8734,
  -36.8933,
  -36.9133,
  -36.9329,
  -36.9517,
  -36.9695,
  -36.9855,
  -37.0022,
  -37.0187,
  -37.035,
  -37.0509,
  -37.0666,
  -37.0826,
  -37.0992,
  -37.117,
  -37.1358,
  -37.1561,
  -37.1779,
  -37.2013,
  -37.2265,
  -37.2539,
  -37.2834,
  -37.3149,
  -37.3494,
  -37.3866,
  -37.4265,
  -37.4691,
  -37.5139,
  -37.56,
  -37.6069,
  -37.6538,
  -37.6999,
  -37.7445,
  -37.7861,
  -37.8267,
  -37.8653,
  -37.9026,
  -37.939,
  -37.975,
  -38.0105,
  -38.0457,
  -38.0802,
  -38.1143,
  -38.1478,
  -38.1806,
  -38.2126,
  -38.2437,
  -38.2739,
  -38.3037,
  -38.3329,
  -38.3618,
  -38.3904,
  -38.4187,
  -38.4466,
  -38.4735,
  -38.4994,
  -38.5241,
  -38.5479,
  -38.5711,
  -38.5939,
  -38.6162,
  -38.6377,
  -38.6581,
  -38.6772,
  -38.6944,
  -38.7086,
  -38.7221,
  -38.7338,
  -38.7442,
  -38.7537,
  -38.7626,
  -38.7711,
  -38.7794,
  -38.7875,
  -38.7957,
  -38.8044,
  -38.8135,
  -38.8227,
  -38.8315,
  -38.8396,
  -38.8469,
  -38.8533,
  -38.8585,
  -38.8623,
  -38.8645,
  -38.865,
  -38.864,
  -38.8616,
  -38.858,
  -38.8535,
  -38.8484,
  -38.8425,
  -38.8358,
  -38.8273,
  -38.8164,
  -38.8032,
  -38.7884,
  -38.7726,
  -38.7568,
  -38.7413,
  -38.7263,
  -38.7111,
  -38.6951,
  -38.6776,
  -38.6568,
  -38.6341,
  -38.608,
  -38.5783,
  -38.5447,
  -38.5073,
  -38.4654,
  -38.4179,
  -38.3636,
  -38.3004,
  -38.2264,
  -38.1411,
  -38.0451,
  -37.9413,
  -37.8363,
  -37.7372,
  -37.651,
  -37.5839,
  -37.539,
  -37.5175,
  -29.813,
  -29.8579,
  -29.9031,
  -29.9485,
  -29.9944,
  -30.0409,
  -30.0882,
  -30.1362,
  -30.185,
  -30.2346,
  -30.2853,
  -30.3362,
  -30.3893,
  -30.4432,
  -30.498,
  -30.5531,
  -30.6081,
  -30.6621,
  -30.7154,
  -30.768,
  -30.8201,
  -30.8721,
  -30.9239,
  -30.9754,
  -31.0266,
  -31.0776,
  -31.1276,
  -31.1785,
  -31.2295,
  -31.2808,
  -31.3324,
  -31.3845,
  -31.4367,
  -31.4889,
  -31.5412,
  -31.5939,
  -31.6469,
  -31.7,
  -31.753,
  -31.8056,
  -31.8577,
  -31.9085,
  -31.9599,
  -32.0108,
  -32.0619,
  -32.1131,
  -32.1648,
  -32.2167,
  -32.2687,
  -32.3202,
  -32.3711,
  -32.4213,
  -32.4708,
  -32.52,
  -32.569,
  -32.6178,
  -32.6664,
  -32.7134,
  -32.7608,
  -32.808,
  -32.8554,
  -32.903,
  -32.9509,
  -32.9988,
  -33.0466,
  -33.0943,
  -33.142,
  -33.1902,
  -33.2391,
  -33.2888,
  -33.3393,
  -33.3905,
  -33.4421,
  -33.4938,
  -33.5441,
  -33.5943,
  -33.6435,
  -33.692,
  -33.74,
  -33.7881,
  -33.8365,
  -33.8848,
  -33.932,
  -33.9784,
  -34.0233,
  -34.0668,
  -34.1094,
  -34.1515,
  -34.1933,
  -34.2351,
  -34.277,
  -34.3194,
  -34.3613,
  -34.4049,
  -34.4486,
  -34.4917,
  -34.5337,
  -34.5743,
  -34.6139,
  -34.6526,
  -34.6908,
  -34.7288,
  -34.7666,
  -34.8042,
  -34.8413,
  -34.8776,
  -34.9132,
  -34.9479,
  -34.9819,
  -35.0154,
  -35.0476,
  -35.0805,
  -35.1133,
  -35.1455,
  -35.1769,
  -35.2075,
  -35.2373,
  -35.2667,
  -35.2959,
  -35.325,
  -35.354,
  -35.3826,
  -35.4106,
  -35.4383,
  -35.4659,
  -35.4934,
  -35.5209,
  -35.5486,
  -35.5765,
  -35.605,
  -35.6332,
  -35.6629,
  -35.6929,
  -35.7229,
  -35.7528,
  -35.7824,
  -35.8119,
  -35.8414,
  -35.8712,
  -35.9014,
  -35.9322,
  -35.9634,
  -35.9949,
  -36.0266,
  -36.0581,
  -36.0896,
  -36.1208,
  -36.1515,
  -36.1813,
  -36.2099,
  -36.2372,
  -36.2633,
  -36.2874,
  -36.312,
  -36.3362,
  -36.3603,
  -36.3843,
  -36.4082,
  -36.432,
  -36.4556,
  -36.4787,
  -36.5008,
  -36.5216,
  -36.5413,
  -36.56,
  -36.5787,
  -36.5978,
  -36.618,
  -36.639,
  -36.6606,
  -36.6821,
  -36.7031,
  -36.7232,
  -36.7426,
  -36.7615,
  -36.7793,
  -36.7985,
  -36.8182,
  -36.8383,
  -36.8586,
  -36.8784,
  -36.8972,
  -36.9146,
  -36.9311,
  -36.9474,
  -36.9635,
  -36.9794,
  -36.9952,
  -37.011,
  -37.0272,
  -37.0443,
  -37.0626,
  -37.0823,
  -37.1032,
  -37.1255,
  -37.1494,
  -37.1751,
  -37.2028,
  -37.2328,
  -37.2654,
  -37.3007,
  -37.3382,
  -37.3795,
  -37.4236,
  -37.4699,
  -37.5177,
  -37.5661,
  -37.6142,
  -37.6613,
  -37.7066,
  -37.7496,
  -37.7904,
  -37.829,
  -37.8663,
  -37.903,
  -37.9392,
  -37.9754,
  -38.0114,
  -38.0466,
  -38.0813,
  -38.1152,
  -38.1479,
  -38.1794,
  -38.2101,
  -38.2396,
  -38.2686,
  -38.2972,
  -38.3256,
  -38.3539,
  -38.3824,
  -38.4107,
  -38.4371,
  -38.4635,
  -38.4884,
  -38.5123,
  -38.5358,
  -38.5588,
  -38.5814,
  -38.6034,
  -38.6241,
  -38.6433,
  -38.6605,
  -38.6755,
  -38.6886,
  -38.7,
  -38.71,
  -38.719,
  -38.7275,
  -38.7356,
  -38.7437,
  -38.7519,
  -38.7603,
  -38.7691,
  -38.7782,
  -38.7875,
  -38.7964,
  -38.8048,
  -38.8124,
  -38.8191,
  -38.8245,
  -38.8283,
  -38.8304,
  -38.8305,
  -38.8289,
  -38.8259,
  -38.8217,
  -38.8168,
  -38.8105,
  -38.805,
  -38.7987,
  -38.7907,
  -38.7804,
  -38.7676,
  -38.7529,
  -38.7371,
  -38.7215,
  -38.7061,
  -38.6914,
  -38.6767,
  -38.6612,
  -38.6442,
  -38.625,
  -38.6027,
  -38.5768,
  -38.547,
  -38.5132,
  -38.4753,
  -38.4326,
  -38.3842,
  -38.3284,
  -38.2634,
  -38.1873,
  -38.0994,
  -38.0012,
  -37.8956,
  -37.789,
  -37.6883,
  -37.601,
  -37.5328,
  -37.4876,
  -37.4659,
  -29.7818,
  -29.8262,
  -29.8708,
  -29.9156,
  -29.9608,
  -30.0069,
  -30.0539,
  -30.1008,
  -30.1496,
  -30.1995,
  -30.2506,
  -30.3029,
  -30.3564,
  -30.411,
  -30.4663,
  -30.5218,
  -30.5769,
  -30.631,
  -30.6844,
  -30.7369,
  -30.7891,
  -30.8402,
  -30.8919,
  -30.9435,
  -30.9949,
  -31.046,
  -31.0972,
  -31.1483,
  -31.1994,
  -31.2504,
  -31.3019,
  -31.3536,
  -31.4055,
  -31.4576,
  -31.5097,
  -31.5619,
  -31.6135,
  -31.6661,
  -31.7184,
  -31.7702,
  -31.8216,
  -31.8727,
  -31.9235,
  -31.9743,
  -32.0253,
  -32.0767,
  -32.1284,
  -32.1801,
  -32.2317,
  -32.2828,
  -32.3332,
  -32.383,
  -32.4312,
  -32.4802,
  -32.5289,
  -32.5772,
  -32.6252,
  -32.6729,
  -32.7204,
  -32.7678,
  -32.8157,
  -32.8639,
  -32.9123,
  -32.9607,
  -33.0087,
  -33.0564,
  -33.104,
  -33.1519,
  -33.2004,
  -33.249,
  -33.2994,
  -33.3506,
  -33.4024,
  -33.4546,
  -33.5063,
  -33.5571,
  -33.607,
  -33.6559,
  -33.7044,
  -33.7526,
  -33.8008,
  -33.8488,
  -33.8959,
  -33.9419,
  -33.9864,
  -34.0297,
  -34.0713,
  -34.1136,
  -34.1559,
  -34.1983,
  -34.2406,
  -34.2833,
  -34.3267,
  -34.3706,
  -34.4146,
  -34.458,
  -34.5003,
  -34.5412,
  -34.5808,
  -34.6194,
  -34.6575,
  -34.6955,
  -34.7334,
  -34.7713,
  -34.8076,
  -34.844,
  -34.8793,
  -34.9136,
  -34.9471,
  -34.9802,
  -35.0132,
  -35.046,
  -35.0787,
  -35.1106,
  -35.1415,
  -35.1715,
  -35.2008,
  -35.2296,
  -35.2581,
  -35.2864,
  -35.3145,
  -35.3422,
  -35.3696,
  -35.3967,
  -35.4227,
  -35.4498,
  -35.4769,
  -35.5042,
  -35.5318,
  -35.5599,
  -35.5886,
  -35.6177,
  -35.647,
  -35.6766,
  -35.706,
  -35.7351,
  -35.7644,
  -35.7936,
  -35.8232,
  -35.8533,
  -35.8839,
  -35.9147,
  -35.9459,
  -35.9773,
  -36.0086,
  -36.0388,
  -36.0699,
  -36.1004,
  -36.1301,
  -36.1587,
  -36.1859,
  -36.212,
  -36.2371,
  -36.2615,
  -36.2856,
  -36.3095,
  -36.3332,
  -36.3569,
  -36.3806,
  -36.404,
  -36.4269,
  -36.4488,
  -36.4694,
  -36.4886,
  -36.507,
  -36.5252,
  -36.544,
  -36.5627,
  -36.5834,
  -36.6049,
  -36.6264,
  -36.6476,
  -36.6679,
  -36.6874,
  -36.7063,
  -36.7251,
  -36.7442,
  -36.7639,
  -36.7842,
  -36.8047,
  -36.8247,
  -36.8437,
  -36.8613,
  -36.8778,
  -36.8937,
  -36.9096,
  -36.9253,
  -36.941,
  -36.9568,
  -36.9731,
  -36.9906,
  -37.0093,
  -37.0285,
  -37.05,
  -37.0729,
  -37.0974,
  -37.1238,
  -37.1522,
  -37.1829,
  -37.2163,
  -37.2524,
  -37.2919,
  -37.3345,
  -37.38,
  -37.4278,
  -37.477,
  -37.5267,
  -37.5759,
  -37.6238,
  -37.6696,
  -37.7129,
  -37.7536,
  -37.7925,
  -37.8297,
  -37.8664,
  -37.9034,
  -37.9402,
  -37.9766,
  -38.0128,
  -38.048,
  -38.0821,
  -38.1138,
  -38.145,
  -38.1749,
  -38.204,
  -38.2322,
  -38.2601,
  -38.288,
  -38.3162,
  -38.3447,
  -38.3733,
  -38.4013,
  -38.428,
  -38.4533,
  -38.4774,
  -38.5008,
  -38.5238,
  -38.5465,
  -38.5685,
  -38.5893,
  -38.6084,
  -38.6255,
  -38.6407,
  -38.6537,
  -38.665,
  -38.6747,
  -38.6836,
  -38.6918,
  -38.7,
  -38.7084,
  -38.717,
  -38.7256,
  -38.7344,
  -38.7434,
  -38.7523,
  -38.76,
  -38.7681,
  -38.7757,
  -38.7825,
  -38.788,
  -38.7917,
  -38.7937,
  -38.7933,
  -38.7911,
  -38.7875,
  -38.7829,
  -38.7779,
  -38.7729,
  -38.7677,
  -38.762,
  -38.7546,
  -38.7448,
  -38.7324,
  -38.7181,
  -38.7029,
  -38.6876,
  -38.6729,
  -38.6587,
  -38.6443,
  -38.6292,
  -38.6124,
  -38.5935,
  -38.5715,
  -38.5458,
  -38.516,
  -38.4818,
  -38.4434,
  -38.4003,
  -38.3511,
  -38.2941,
  -38.2274,
  -38.1491,
  -38.0587,
  -37.9574,
  -37.8491,
  -37.7395,
  -37.6361,
  -37.5463,
  -37.4764,
  -37.4292,
  -37.4069,
  -29.7519,
  -29.7957,
  -29.8387,
  -29.883,
  -29.9279,
  -29.9736,
  -30.0205,
  -30.0686,
  -30.1176,
  -30.1678,
  -30.2192,
  -30.2718,
  -30.3257,
  -30.3805,
  -30.436,
  -30.4919,
  -30.547,
  -30.6003,
  -30.6537,
  -30.7062,
  -30.7585,
  -30.8105,
  -30.8623,
  -30.9139,
  -30.9654,
  -31.0166,
  -31.0678,
  -31.1189,
  -31.1699,
  -31.2208,
  -31.272,
  -31.3235,
  -31.3743,
  -31.4261,
  -31.4779,
  -31.5298,
  -31.5818,
  -31.6338,
  -31.6853,
  -31.7363,
  -31.787,
  -31.8374,
  -31.8878,
  -31.9386,
  -31.9897,
  -32.0411,
  -32.0926,
  -32.1429,
  -32.1937,
  -32.244,
  -32.2938,
  -32.3429,
  -32.3918,
  -32.4404,
  -32.4888,
  -32.537,
  -32.5849,
  -32.6327,
  -32.6805,
  -32.7286,
  -32.7771,
  -32.8258,
  -32.8745,
  -32.9221,
  -32.9703,
  -33.0179,
  -33.0654,
  -33.1132,
  -33.1617,
  -33.2111,
  -33.2616,
  -33.313,
  -33.3653,
  -33.4177,
  -33.4699,
  -33.5213,
  -33.5715,
  -33.621,
  -33.6697,
  -33.7181,
  -33.7653,
  -33.8129,
  -33.8595,
  -33.905,
  -33.9493,
  -33.9926,
  -34.0354,
  -34.078,
  -34.1207,
  -34.1636,
  -34.2065,
  -34.2495,
  -34.293,
  -34.337,
  -34.381,
  -34.4246,
  -34.467,
  -34.508,
  -34.5468,
  -34.5856,
  -34.6239,
  -34.6622,
  -34.7004,
  -34.7385,
  -34.776,
  -34.8124,
  -34.8474,
  -34.8812,
  -34.9142,
  -34.9469,
  -34.9796,
  -35.0121,
  -35.0444,
  -35.076,
  -35.1065,
  -35.1359,
  -35.1645,
  -35.1915,
  -35.2191,
  -35.2466,
  -35.2738,
  -35.3006,
  -35.3272,
  -35.3538,
  -35.3806,
  -35.4074,
  -35.4342,
  -35.4612,
  -35.4885,
  -35.5162,
  -35.5444,
  -35.5727,
  -35.6014,
  -35.6303,
  -35.6594,
  -35.6883,
  -35.7173,
  -35.7465,
  -35.7749,
  -35.8048,
  -35.8349,
  -35.8653,
  -35.8958,
  -35.9265,
  -35.9573,
  -35.9881,
  -36.0187,
  -36.0489,
  -36.0783,
  -36.1065,
  -36.1337,
  -36.1596,
  -36.1847,
  -36.2092,
  -36.2333,
  -36.2571,
  -36.2807,
  -36.3044,
  -36.3281,
  -36.3515,
  -36.3734,
  -36.3952,
  -36.4156,
  -36.4347,
  -36.453,
  -36.4709,
  -36.4896,
  -36.5091,
  -36.5296,
  -36.5508,
  -36.5725,
  -36.5937,
  -36.6142,
  -36.6338,
  -36.6528,
  -36.6715,
  -36.6903,
  -36.7097,
  -36.7299,
  -36.7505,
  -36.7707,
  -36.7898,
  -36.8077,
  -36.8246,
  -36.8399,
  -36.8558,
  -36.8715,
  -36.8871,
  -36.9029,
  -36.9192,
  -36.9368,
  -36.9558,
  -36.9763,
  -36.9983,
  -37.0217,
  -37.0469,
  -37.0741,
  -37.1033,
  -37.135,
  -37.1692,
  -37.2063,
  -37.2469,
  -37.2907,
  -37.3375,
  -37.3867,
  -37.4375,
  -37.4885,
  -37.5387,
  -37.5872,
  -37.6333,
  -37.6767,
  -37.7164,
  -37.7553,
  -37.7927,
  -37.8294,
  -37.8665,
  -37.9039,
  -37.9411,
  -37.978,
  -38.0137,
  -38.0479,
  -38.0805,
  -38.1114,
  -38.1407,
  -38.169,
  -38.1967,
  -38.2241,
  -38.2514,
  -38.2795,
  -38.308,
  -38.3368,
  -38.365,
  -38.392,
  -38.4174,
  -38.4417,
  -38.465,
  -38.4878,
  -38.5103,
  -38.5321,
  -38.5528,
  -38.5719,
  -38.5891,
  -38.6042,
  -38.6165,
  -38.6278,
  -38.6376,
  -38.6464,
  -38.6548,
  -38.6632,
  -38.6719,
  -38.6808,
  -38.6897,
  -38.6985,
  -38.7071,
  -38.7156,
  -38.7239,
  -38.7317,
  -38.7389,
  -38.7453,
  -38.7507,
  -38.7545,
  -38.7562,
  -38.7555,
  -38.7533,
  -38.7493,
  -38.7448,
  -38.7398,
  -38.735,
  -38.7303,
  -38.7249,
  -38.718,
  -38.7086,
  -38.6968,
  -38.6832,
  -38.6687,
  -38.6543,
  -38.6404,
  -38.6267,
  -38.6127,
  -38.5977,
  -38.5811,
  -38.5623,
  -38.5404,
  -38.5138,
  -38.484,
  -38.4499,
  -38.4112,
  -38.3676,
  -38.3179,
  -38.2599,
  -38.1916,
  -38.1111,
  -38.0178,
  -37.9132,
  -37.8014,
  -37.6877,
  -37.5806,
  -37.4871,
  -37.4146,
  -37.3663,
  -37.3432,
  -29.7225,
  -29.7661,
  -29.8095,
  -29.8532,
  -29.8977,
  -29.9433,
  -29.9902,
  -30.0385,
  -30.0881,
  -30.1387,
  -30.1904,
  -30.243,
  -30.296,
  -30.3509,
  -30.4065,
  -30.4622,
  -30.5173,
  -30.5715,
  -30.6249,
  -30.6775,
  -30.7297,
  -30.7817,
  -30.8335,
  -30.8852,
  -30.9367,
  -30.988,
  -31.0391,
  -31.089,
  -31.1398,
  -31.1905,
  -31.2415,
  -31.2929,
  -31.3446,
  -31.3963,
  -31.448,
  -31.4994,
  -31.5509,
  -31.6021,
  -31.6527,
  -31.7028,
  -31.7526,
  -31.8025,
  -31.8517,
  -31.9025,
  -31.9536,
  -32.0052,
  -32.0565,
  -32.1071,
  -32.157,
  -32.2062,
  -32.2549,
  -32.3033,
  -32.3516,
  -32.4,
  -32.4482,
  -32.4965,
  -32.5448,
  -32.5932,
  -32.6407,
  -32.6894,
  -32.7385,
  -32.7876,
  -32.8364,
  -32.885,
  -32.9331,
  -32.9807,
  -33.0281,
  -33.0758,
  -33.1242,
  -33.1737,
  -33.2245,
  -33.2763,
  -33.329,
  -33.3819,
  -33.4345,
  -33.4854,
  -33.5361,
  -33.5859,
  -33.635,
  -33.6834,
  -33.7313,
  -33.7786,
  -33.8248,
  -33.8698,
  -33.914,
  -33.9571,
  -34.0001,
  -34.0434,
  -34.0867,
  -34.1299,
  -34.1731,
  -34.2164,
  -34.259,
  -34.3029,
  -34.3468,
  -34.3901,
  -34.4325,
  -34.4736,
  -34.5135,
  -34.5527,
  -34.5913,
  -34.6299,
  -34.6686,
  -34.707,
  -34.7447,
  -34.7808,
  -34.8156,
  -34.849,
  -34.8818,
  -34.914,
  -34.9462,
  -34.9773,
  -35.009,
  -35.0401,
  -35.0701,
  -35.099,
  -35.1269,
  -35.154,
  -35.1807,
  -35.2072,
  -35.2334,
  -35.2596,
  -35.2856,
  -35.3119,
  -35.3384,
  -35.365,
  -35.3917,
  -35.4185,
  -35.4458,
  -35.4731,
  -35.5007,
  -35.5274,
  -35.5552,
  -35.5836,
  -35.6122,
  -35.6409,
  -35.6699,
  -35.699,
  -35.7284,
  -35.758,
  -35.7875,
  -35.8172,
  -35.8467,
  -35.8765,
  -35.9065,
  -35.9366,
  -35.9667,
  -35.9963,
  -36.0253,
  -36.0532,
  -36.08,
  -36.1058,
  -36.1309,
  -36.1543,
  -36.1785,
  -36.2024,
  -36.2261,
  -36.2499,
  -36.2737,
  -36.2972,
  -36.3201,
  -36.3419,
  -36.3625,
  -36.3818,
  -36.4002,
  -36.4183,
  -36.4367,
  -36.4563,
  -36.4766,
  -36.4977,
  -36.519,
  -36.5402,
  -36.5608,
  -36.5806,
  -36.5995,
  -36.618,
  -36.6355,
  -36.6547,
  -36.6744,
  -36.6947,
  -36.7149,
  -36.7344,
  -36.7529,
  -36.7705,
  -36.7873,
  -36.8036,
  -36.8194,
  -36.835,
  -36.8507,
  -36.8672,
  -36.8847,
  -36.9037,
  -36.9244,
  -36.9466,
  -36.9706,
  -36.9966,
  -37.0249,
  -37.0552,
  -37.088,
  -37.1234,
  -37.1618,
  -37.2035,
  -37.2475,
  -37.2956,
  -37.3462,
  -37.3982,
  -37.4504,
  -37.5015,
  -37.5504,
  -37.5966,
  -37.6399,
  -37.6806,
  -37.7191,
  -37.7567,
  -37.7939,
  -37.8313,
  -37.8692,
  -37.9072,
  -37.9445,
  -37.9805,
  -38.0149,
  -38.0472,
  -38.0775,
  -38.1061,
  -38.1334,
  -38.1603,
  -38.1874,
  -38.2147,
  -38.2428,
  -38.2713,
  -38.3001,
  -38.3284,
  -38.3544,
  -38.38,
  -38.4041,
  -38.4273,
  -38.4499,
  -38.4719,
  -38.4933,
  -38.5137,
  -38.5326,
  -38.55,
  -38.5656,
  -38.5791,
  -38.5906,
  -38.6006,
  -38.6096,
  -38.6182,
  -38.6268,
  -38.6358,
  -38.6447,
  -38.6537,
  -38.6624,
  -38.6705,
  -38.6784,
  -38.686,
  -38.6935,
  -38.7003,
  -38.7064,
  -38.7115,
  -38.7151,
  -38.7166,
  -38.7162,
  -38.7139,
  -38.7101,
  -38.7059,
  -38.7014,
  -38.697,
  -38.6926,
  -38.6866,
  -38.6799,
  -38.6709,
  -38.6597,
  -38.6469,
  -38.6334,
  -38.6199,
  -38.6068,
  -38.5938,
  -38.5802,
  -38.5653,
  -38.5487,
  -38.5298,
  -38.508,
  -38.4825,
  -38.4527,
  -38.4186,
  -38.3799,
  -38.3363,
  -38.2862,
  -38.2273,
  -38.1576,
  -38.075,
  -37.9792,
  -37.8711,
  -37.755,
  -37.6367,
  -37.5253,
  -37.427,
  -37.3506,
  -37.2999,
  -37.2761,
  -29.6952,
  -29.7388,
  -29.7822,
  -29.8256,
  -29.8697,
  -29.9151,
  -29.9621,
  -30.0096,
  -30.0595,
  -30.1105,
  -30.1623,
  -30.215,
  -30.2688,
  -30.3236,
  -30.379,
  -30.4345,
  -30.4894,
  -30.5434,
  -30.5966,
  -30.6492,
  -30.7013,
  -30.7533,
  -30.8041,
  -30.8558,
  -30.9073,
  -30.9586,
  -31.0096,
  -31.0603,
  -31.1109,
  -31.1614,
  -31.2122,
  -31.2635,
  -31.3151,
  -31.3668,
  -31.4183,
  -31.4693,
  -31.5202,
  -31.5695,
  -31.6192,
  -31.6684,
  -31.7176,
  -31.767,
  -31.8171,
  -31.8679,
  -31.9191,
  -31.9705,
  -32.0213,
  -32.0713,
  -32.1203,
  -32.1686,
  -32.2164,
  -32.264,
  -32.3119,
  -32.3589,
  -32.4072,
  -32.4557,
  -32.5044,
  -32.5535,
  -32.6029,
  -32.6525,
  -32.7019,
  -32.7511,
  -32.7999,
  -32.8482,
  -32.8963,
  -32.9439,
  -32.9914,
  -33.0391,
  -33.0876,
  -33.1361,
  -33.187,
  -33.2391,
  -33.2922,
  -33.3455,
  -33.3985,
  -33.4508,
  -33.5019,
  -33.5521,
  -33.6014,
  -33.6499,
  -33.6976,
  -33.7445,
  -33.7903,
  -33.835,
  -33.8792,
  -33.9227,
  -33.9663,
  -34.0089,
  -34.0526,
  -34.096,
  -34.1393,
  -34.1825,
  -34.226,
  -34.2698,
  -34.3134,
  -34.3565,
  -34.3987,
  -34.4398,
  -34.4801,
  -34.5196,
  -34.5588,
  -34.5978,
  -34.6367,
  -34.6752,
  -34.7127,
  -34.7476,
  -34.782,
  -34.8152,
  -34.8477,
  -34.8795,
  -34.9115,
  -34.9431,
  -34.9744,
  -35.0051,
  -35.0345,
  -35.0628,
  -35.0899,
  -35.1163,
  -35.1421,
  -35.1677,
  -35.1931,
  -35.2185,
  -35.2442,
  -35.2703,
  -35.2966,
  -35.3221,
  -35.3487,
  -35.3754,
  -35.4025,
  -35.4295,
  -35.4564,
  -35.4838,
  -35.5109,
  -35.5383,
  -35.5666,
  -35.5952,
  -35.6242,
  -35.6534,
  -35.6825,
  -35.7117,
  -35.7406,
  -35.7692,
  -35.7978,
  -35.8266,
  -35.8556,
  -35.8849,
  -35.9134,
  -35.9424,
  -35.9708,
  -35.9983,
  -36.0248,
  -36.0504,
  -36.0753,
  -36.0999,
  -36.1242,
  -36.1483,
  -36.1722,
  -36.1962,
  -36.2201,
  -36.2437,
  -36.2666,
  -36.2885,
  -36.3091,
  -36.3287,
  -36.3473,
  -36.3659,
  -36.3844,
  -36.4039,
  -36.4228,
  -36.4436,
  -36.4647,
  -36.4858,
  -36.5063,
  -36.5261,
  -36.5451,
  -36.5636,
  -36.582,
  -36.6008,
  -36.6201,
  -36.6398,
  -36.66,
  -36.6799,
  -36.6987,
  -36.7172,
  -36.7349,
  -36.7518,
  -36.7679,
  -36.7834,
  -36.7991,
  -36.8155,
  -36.8329,
  -36.8521,
  -36.8728,
  -36.8955,
  -36.9189,
  -36.946,
  -36.9755,
  -37.0072,
  -37.0414,
  -37.0784,
  -37.1183,
  -37.1614,
  -37.2078,
  -37.2571,
  -37.3088,
  -37.3617,
  -37.4146,
  -37.4662,
  -37.5153,
  -37.5614,
  -37.6045,
  -37.645,
  -37.6835,
  -37.7211,
  -37.7587,
  -37.7968,
  -37.8353,
  -37.8738,
  -37.9114,
  -37.9475,
  -37.9817,
  -38.0135,
  -38.0422,
  -38.0699,
  -38.0965,
  -38.1226,
  -38.1492,
  -38.1763,
  -38.2046,
  -38.2333,
  -38.2621,
  -38.2902,
  -38.317,
  -38.3424,
  -38.3665,
  -38.3896,
  -38.4119,
  -38.4337,
  -38.4547,
  -38.4748,
  -38.4937,
  -38.5112,
  -38.5271,
  -38.5409,
  -38.5528,
  -38.563,
  -38.5721,
  -38.5808,
  -38.5895,
  -38.5985,
  -38.6073,
  -38.6162,
  -38.6244,
  -38.6325,
  -38.6397,
  -38.6469,
  -38.6524,
  -38.6586,
  -38.6642,
  -38.6691,
  -38.6725,
  -38.6743,
  -38.6741,
  -38.6724,
  -38.6694,
  -38.6658,
  -38.6619,
  -38.658,
  -38.6539,
  -38.6489,
  -38.6424,
  -38.6338,
  -38.6234,
  -38.6115,
  -38.5988,
  -38.5862,
  -38.5739,
  -38.5615,
  -38.5484,
  -38.5338,
  -38.5173,
  -38.4983,
  -38.4763,
  -38.4507,
  -38.421,
  -38.3869,
  -38.3484,
  -38.3048,
  -38.2544,
  -38.1951,
  -38.1242,
  -38.0397,
  -37.9409,
  -37.8295,
  -37.7093,
  -37.5865,
  -37.4696,
  -37.3663,
  -37.2849,
  -37.231,
  -37.2059,
  -29.6693,
  -29.7132,
  -29.7565,
  -29.799,
  -29.843,
  -29.8883,
  -29.9352,
  -29.9837,
  -30.0337,
  -30.0845,
  -30.1363,
  -30.189,
  -30.2426,
  -30.2971,
  -30.3523,
  -30.4075,
  -30.4622,
  -30.515,
  -30.568,
  -30.6204,
  -30.6723,
  -30.7242,
  -30.776,
  -30.8277,
  -30.8792,
  -30.9304,
  -30.9813,
  -31.0318,
  -31.082,
  -31.1323,
  -31.1829,
  -31.2341,
  -31.2846,
  -31.3361,
  -31.3874,
  -31.4381,
  -31.4882,
  -31.5377,
  -31.5866,
  -31.6351,
  -31.6837,
  -31.7328,
  -31.7827,
  -31.8334,
  -31.8846,
  -31.9356,
  -31.9859,
  -32.0352,
  -32.0826,
  -32.1302,
  -32.1775,
  -32.2248,
  -32.2723,
  -32.3202,
  -32.3686,
  -32.4173,
  -32.4666,
  -32.5164,
  -32.5665,
  -32.6166,
  -32.6664,
  -32.7156,
  -32.7643,
  -32.8125,
  -32.8594,
  -32.907,
  -32.9546,
  -33.0023,
  -33.0507,
  -33.1001,
  -33.1511,
  -33.2034,
  -33.2567,
  -33.3103,
  -33.3635,
  -33.4159,
  -33.4673,
  -33.5177,
  -33.5672,
  -33.6159,
  -33.6635,
  -33.7092,
  -33.7548,
  -33.7996,
  -33.844,
  -33.8881,
  -33.9323,
  -33.9764,
  -34.0203,
  -34.0637,
  -34.1068,
  -34.1498,
  -34.193,
  -34.2365,
  -34.2798,
  -34.3227,
  -34.3648,
  -34.4062,
  -34.4469,
  -34.4859,
  -34.5254,
  -34.5647,
  -34.6036,
  -34.6417,
  -34.6787,
  -34.7142,
  -34.7483,
  -34.7812,
  -34.8135,
  -34.8453,
  -34.8771,
  -34.9084,
  -34.9394,
  -34.9696,
  -34.9986,
  -35.0264,
  -35.0528,
  -35.0783,
  -35.1024,
  -35.1273,
  -35.1522,
  -35.1773,
  -35.2028,
  -35.2287,
  -35.2548,
  -35.2811,
  -35.3074,
  -35.3338,
  -35.3607,
  -35.3875,
  -35.4139,
  -35.4404,
  -35.4671,
  -35.4939,
  -35.5218,
  -35.5503,
  -35.5791,
  -35.6083,
  -35.6371,
  -35.6648,
  -35.693,
  -35.7207,
  -35.7482,
  -35.7758,
  -35.804,
  -35.8326,
  -35.8614,
  -35.8898,
  -35.9177,
  -35.9447,
  -35.9708,
  -35.9963,
  -36.0211,
  -36.0457,
  -36.0701,
  -36.0944,
  -36.1186,
  -36.1427,
  -36.1667,
  -36.1903,
  -36.2132,
  -36.234,
  -36.2548,
  -36.2744,
  -36.2934,
  -36.312,
  -36.3306,
  -36.3499,
  -36.3698,
  -36.3903,
  -36.4111,
  -36.432,
  -36.4525,
  -36.4724,
  -36.4916,
  -36.5103,
  -36.5287,
  -36.5472,
  -36.5661,
  -36.5855,
  -36.6054,
  -36.6254,
  -36.645,
  -36.6643,
  -36.6827,
  -36.6991,
  -36.7154,
  -36.7314,
  -36.7471,
  -36.7634,
  -36.781,
  -36.8001,
  -36.8207,
  -36.8436,
  -36.8691,
  -36.8974,
  -36.9281,
  -36.9616,
  -36.9978,
  -37.0366,
  -37.0782,
  -37.1229,
  -37.1705,
  -37.221,
  -37.2734,
  -37.3268,
  -37.38,
  -37.4316,
  -37.4805,
  -37.5264,
  -37.5693,
  -37.6096,
  -37.6482,
  -37.6852,
  -37.7232,
  -37.7619,
  -37.8009,
  -37.8397,
  -37.8774,
  -37.9133,
  -37.947,
  -37.9783,
  -38.0071,
  -38.034,
  -38.0597,
  -38.0851,
  -38.1113,
  -38.1385,
  -38.1669,
  -38.1956,
  -38.2243,
  -38.2521,
  -38.2787,
  -38.3038,
  -38.3278,
  -38.3508,
  -38.3731,
  -38.3947,
  -38.4156,
  -38.4356,
  -38.4546,
  -38.4723,
  -38.4883,
  -38.5024,
  -38.5144,
  -38.5238,
  -38.5329,
  -38.5416,
  -38.55,
  -38.5588,
  -38.5674,
  -38.5757,
  -38.5837,
  -38.5914,
  -38.5982,
  -38.6044,
  -38.6104,
  -38.6159,
  -38.6211,
  -38.6257,
  -38.6291,
  -38.6313,
  -38.6318,
  -38.6311,
  -38.6291,
  -38.6264,
  -38.6233,
  -38.6197,
  -38.6157,
  -38.6106,
  -38.6041,
  -38.5959,
  -38.5861,
  -38.5749,
  -38.5631,
  -38.5514,
  -38.5398,
  -38.5281,
  -38.5157,
  -38.5016,
  -38.4853,
  -38.4663,
  -38.4441,
  -38.4183,
  -38.3886,
  -38.3536,
  -38.3152,
  -38.2718,
  -38.2214,
  -38.1615,
  -38.0894,
  -38.0033,
  -37.902,
  -37.7877,
  -37.663,
  -37.5361,
  -37.4134,
  -37.3043,
  -37.2179,
  -37.1605,
  -37.1342,
  -29.6433,
  -29.6876,
  -29.7315,
  -29.7753,
  -29.8194,
  -29.8647,
  -29.9114,
  -29.9598,
  -30.0093,
  -30.06,
  -30.1114,
  -30.1638,
  -30.2171,
  -30.2703,
  -30.3252,
  -30.3802,
  -30.4346,
  -30.4883,
  -30.5412,
  -30.5933,
  -30.6452,
  -30.6969,
  -30.7484,
  -30.8001,
  -30.8515,
  -30.9026,
  -30.9533,
  -31.0025,
  -31.0524,
  -31.1023,
  -31.1527,
  -31.2036,
  -31.2548,
  -31.3061,
  -31.3569,
  -31.4072,
  -31.4568,
  -31.5057,
  -31.5541,
  -31.6021,
  -31.6503,
  -31.6991,
  -31.7488,
  -31.7982,
  -31.849,
  -31.8996,
  -31.9493,
  -31.9981,
  -32.0461,
  -32.0934,
  -32.1407,
  -32.188,
  -32.2357,
  -32.2837,
  -32.3322,
  -32.3812,
  -32.4308,
  -32.481,
  -32.5316,
  -32.5811,
  -32.631,
  -32.6803,
  -32.7289,
  -32.7769,
  -32.8247,
  -32.8723,
  -32.9199,
  -32.9676,
  -33.016,
  -33.0653,
  -33.1161,
  -33.1684,
  -33.2216,
  -33.2751,
  -33.3283,
  -33.3806,
  -33.4311,
  -33.4817,
  -33.5312,
  -33.5799,
  -33.6277,
  -33.6745,
  -33.7201,
  -33.7654,
  -33.8102,
  -33.855,
  -33.8998,
  -33.9444,
  -33.9884,
  -34.0318,
  -34.0746,
  -34.1172,
  -34.16,
  -34.2021,
  -34.2452,
  -34.288,
  -34.3304,
  -34.372,
  -34.4131,
  -34.4535,
  -34.4933,
  -34.5324,
  -34.5709,
  -34.6084,
  -34.6447,
  -34.6796,
  -34.7133,
  -34.7461,
  -34.7784,
  -34.8104,
  -34.842,
  -34.8732,
  -34.9029,
  -34.9327,
  -34.9613,
  -34.9885,
  -35.0145,
  -35.0394,
  -35.064,
  -35.0883,
  -35.1129,
  -35.1379,
  -35.1632,
  -35.1891,
  -35.215,
  -35.2409,
  -35.2668,
  -35.2928,
  -35.3191,
  -35.3455,
  -35.3716,
  -35.3974,
  -35.4224,
  -35.4488,
  -35.4764,
  -35.5047,
  -35.5336,
  -35.5627,
  -35.5914,
  -35.6196,
  -35.6469,
  -35.6738,
  -35.7003,
  -35.7271,
  -35.7544,
  -35.7822,
  -35.8103,
  -35.8382,
  -35.8655,
  -35.8921,
  -35.9179,
  -35.9431,
  -35.9678,
  -35.9924,
  -36.0159,
  -36.0403,
  -36.0647,
  -36.089,
  -36.113,
  -36.1366,
  -36.1594,
  -36.1813,
  -36.202,
  -36.2215,
  -36.2404,
  -36.259,
  -36.2777,
  -36.2968,
  -36.3166,
  -36.337,
  -36.3577,
  -36.3783,
  -36.3988,
  -36.4188,
  -36.4382,
  -36.4571,
  -36.4756,
  -36.4931,
  -36.5118,
  -36.531,
  -36.5507,
  -36.5708,
  -36.5909,
  -36.6107,
  -36.6297,
  -36.6478,
  -36.6646,
  -36.6806,
  -36.6965,
  -36.7129,
  -36.7305,
  -36.7496,
  -36.7707,
  -36.7941,
  -36.8204,
  -36.8498,
  -36.8823,
  -36.9177,
  -36.9558,
  -36.9967,
  -37.0403,
  -37.0867,
  -37.1356,
  -37.1869,
  -37.2389,
  -37.2926,
  -37.3456,
  -37.3968,
  -37.4453,
  -37.4908,
  -37.5334,
  -37.5737,
  -37.6125,
  -37.6509,
  -37.6895,
  -37.7286,
  -37.7679,
  -37.8067,
  -37.8443,
  -37.8797,
  -37.9128,
  -37.9433,
  -37.9713,
  -37.9973,
  -38.0223,
  -38.0472,
  -38.0731,
  -38.1002,
  -38.1284,
  -38.1572,
  -38.1856,
  -38.213,
  -38.2392,
  -38.2642,
  -38.287,
  -38.31,
  -38.3323,
  -38.3539,
  -38.3749,
  -38.3951,
  -38.4143,
  -38.4323,
  -38.4481,
  -38.4624,
  -38.4746,
  -38.4849,
  -38.4939,
  -38.5023,
  -38.5104,
  -38.5187,
  -38.527,
  -38.5351,
  -38.5427,
  -38.5497,
  -38.556,
  -38.5616,
  -38.5666,
  -38.5715,
  -38.5762,
  -38.5804,
  -38.5841,
  -38.5867,
  -38.5883,
  -38.5886,
  -38.5879,
  -38.5863,
  -38.5838,
  -38.5806,
  -38.5764,
  -38.5712,
  -38.5646,
  -38.5555,
  -38.5461,
  -38.5357,
  -38.5246,
  -38.5135,
  -38.5027,
  -38.4919,
  -38.4803,
  -38.4669,
  -38.4511,
  -38.4323,
  -38.4102,
  -38.3842,
  -38.3543,
  -38.3203,
  -38.2822,
  -38.2387,
  -38.1882,
  -38.1279,
  -38.055,
  -37.9674,
  -37.8642,
  -37.747,
  -37.6193,
  -37.4877,
  -37.36,
  -37.2458,
  -37.1548,
  -37.0934,
  -37.0651,
  -29.6189,
  -29.664,
  -29.7086,
  -29.7531,
  -29.7978,
  -29.8433,
  -29.89,
  -29.9379,
  -29.9859,
  -30.0361,
  -30.087,
  -30.1389,
  -30.1918,
  -30.2456,
  -30.3001,
  -30.3545,
  -30.4089,
  -30.4625,
  -30.5152,
  -30.5673,
  -30.619,
  -30.6705,
  -30.7219,
  -30.7722,
  -30.8233,
  -30.8741,
  -30.9245,
  -30.9744,
  -31.024,
  -31.0736,
  -31.1236,
  -31.1741,
  -31.225,
  -31.2758,
  -31.3262,
  -31.3761,
  -31.4254,
  -31.474,
  -31.521,
  -31.5688,
  -31.6167,
  -31.6652,
  -31.7146,
  -31.7646,
  -31.815,
  -31.865,
  -31.9142,
  -31.9627,
  -32.0106,
  -32.058,
  -32.1054,
  -32.1531,
  -32.201,
  -32.2494,
  -32.2971,
  -32.3464,
  -32.3962,
  -32.4466,
  -32.4972,
  -32.5479,
  -32.598,
  -32.6473,
  -32.6958,
  -32.7437,
  -32.7913,
  -32.8389,
  -32.8865,
  -32.9343,
  -32.9825,
  -33.0317,
  -33.0813,
  -33.1331,
  -33.186,
  -33.2391,
  -33.2919,
  -33.3439,
  -33.3952,
  -33.4455,
  -33.4952,
  -33.5441,
  -33.5921,
  -33.6392,
  -33.6854,
  -33.7311,
  -33.7766,
  -33.822,
  -33.8673,
  -33.9123,
  -33.9555,
  -33.9989,
  -34.0415,
  -34.0837,
  -34.1261,
  -34.1688,
  -34.2117,
  -34.2546,
  -34.2972,
  -34.3393,
  -34.3809,
  -34.4217,
  -34.4614,
  -34.5003,
  -34.5381,
  -34.5748,
  -34.6101,
  -34.6443,
  -34.6766,
  -34.7094,
  -34.7417,
  -34.7737,
  -34.8055,
  -34.8366,
  -34.8671,
  -34.8966,
  -34.9249,
  -34.9518,
  -34.9774,
  -35.002,
  -35.0261,
  -35.0502,
  -35.0746,
  -35.0994,
  -35.1247,
  -35.1503,
  -35.1759,
  -35.2014,
  -35.2257,
  -35.2511,
  -35.2767,
  -35.3025,
  -35.3281,
  -35.3535,
  -35.3791,
  -35.4053,
  -35.4325,
  -35.4607,
  -35.4896,
  -35.5185,
  -35.5468,
  -35.5745,
  -35.6014,
  -35.6275,
  -35.6533,
  -35.6794,
  -35.7059,
  -35.7331,
  -35.7605,
  -35.7868,
  -35.8136,
  -35.8398,
  -35.8653,
  -35.8903,
  -35.9149,
  -35.9394,
  -35.9638,
  -35.9882,
  -36.0127,
  -36.0371,
  -36.0613,
  -36.085,
  -36.1078,
  -36.1295,
  -36.1501,
  -36.1693,
  -36.188,
  -36.2064,
  -36.225,
  -36.2442,
  -36.264,
  -36.2834,
  -36.304,
  -36.3246,
  -36.3449,
  -36.3649,
  -36.3844,
  -36.4035,
  -36.4221,
  -36.4406,
  -36.4591,
  -36.4782,
  -36.4979,
  -36.518,
  -36.5384,
  -36.5587,
  -36.5783,
  -36.5968,
  -36.6141,
  -36.6305,
  -36.6466,
  -36.6632,
  -36.6809,
  -36.7002,
  -36.7217,
  -36.7458,
  -36.773,
  -36.8027,
  -36.8367,
  -36.874,
  -36.9143,
  -36.9574,
  -37.003,
  -37.0511,
  -37.1014,
  -37.1536,
  -37.2071,
  -37.2608,
  -37.3136,
  -37.3643,
  -37.412,
  -37.4569,
  -37.4992,
  -37.5395,
  -37.5785,
  -37.6174,
  -37.6563,
  -37.6956,
  -37.735,
  -37.7737,
  -37.8108,
  -37.8457,
  -37.878,
  -37.9077,
  -37.9349,
  -37.9604,
  -37.9837,
  -38.0082,
  -38.0337,
  -38.0605,
  -38.0884,
  -38.1169,
  -38.1449,
  -38.172,
  -38.1979,
  -38.2226,
  -38.2464,
  -38.2694,
  -38.2918,
  -38.3136,
  -38.3349,
  -38.3554,
  -38.3748,
  -38.3929,
  -38.4089,
  -38.423,
  -38.4349,
  -38.4448,
  -38.4537,
  -38.4619,
  -38.4698,
  -38.4778,
  -38.4857,
  -38.4935,
  -38.5009,
  -38.5074,
  -38.5128,
  -38.5175,
  -38.5216,
  -38.5257,
  -38.5287,
  -38.5326,
  -38.5365,
  -38.5396,
  -38.5421,
  -38.5437,
  -38.5443,
  -38.5436,
  -38.5418,
  -38.5388,
  -38.5347,
  -38.5292,
  -38.5222,
  -38.514,
  -38.5048,
  -38.4947,
  -38.4844,
  -38.4741,
  -38.4642,
  -38.4543,
  -38.4436,
  -38.4311,
  -38.416,
  -38.3977,
  -38.3757,
  -38.3498,
  -38.3198,
  -38.2858,
  -38.2476,
  -38.2041,
  -38.1534,
  -38.0928,
  -38.0193,
  -37.9309,
  -37.8264,
  -37.7072,
  -37.5769,
  -37.4418,
  -37.3101,
  -37.1917,
  -37.0961,
  -37.0311,
  -36.9999,
  -29.5951,
  -29.641,
  -29.6867,
  -29.732,
  -29.7767,
  -29.8227,
  -29.8695,
  -29.917,
  -29.9654,
  -30.0148,
  -30.0652,
  -30.1167,
  -30.1691,
  -30.2223,
  -30.2762,
  -30.3302,
  -30.3842,
  -30.4376,
  -30.4894,
  -30.5415,
  -30.593,
  -30.6442,
  -30.6951,
  -30.7459,
  -30.7965,
  -30.8469,
  -30.8971,
  -30.9468,
  -30.9962,
  -31.0455,
  -31.095,
  -31.1449,
  -31.1951,
  -31.2443,
  -31.2942,
  -31.3439,
  -31.393,
  -31.4416,
  -31.4897,
  -31.5374,
  -31.5852,
  -31.6334,
  -31.6823,
  -31.7318,
  -31.7815,
  -31.831,
  -31.8798,
  -31.928,
  -31.9761,
  -32.023,
  -32.071,
  -32.1192,
  -32.1677,
  -32.2164,
  -32.2654,
  -32.3148,
  -32.3646,
  -32.4149,
  -32.4655,
  -32.516,
  -32.5661,
  -32.6155,
  -32.6639,
  -32.7117,
  -32.7592,
  -32.8057,
  -32.8534,
  -32.9013,
  -32.9496,
  -32.9987,
  -33.0487,
  -33.1001,
  -33.1522,
  -33.2045,
  -33.2565,
  -33.3081,
  -33.3589,
  -33.4091,
  -33.4589,
  -33.5081,
  -33.5564,
  -33.604,
  -33.6497,
  -33.696,
  -33.7421,
  -33.7879,
  -33.8337,
  -33.879,
  -33.9234,
  -33.9669,
  -34.0094,
  -34.0514,
  -34.0936,
  -34.136,
  -34.1787,
  -34.2216,
  -34.2646,
  -34.3072,
  -34.3492,
  -34.3902,
  -34.429,
  -34.4674,
  -34.5043,
  -34.54,
  -34.5745,
  -34.6081,
  -34.6411,
  -34.6736,
  -34.7059,
  -34.7381,
  -34.7699,
  -34.8011,
  -34.8315,
  -34.8608,
  -34.8888,
  -34.9155,
  -34.941,
  -34.9656,
  -34.9894,
  -35.0122,
  -35.0365,
  -35.061,
  -35.0861,
  -35.1113,
  -35.1364,
  -35.1612,
  -35.186,
  -35.2107,
  -35.2356,
  -35.2607,
  -35.2859,
  -35.311,
  -35.3363,
  -35.3622,
  -35.3891,
  -35.4171,
  -35.4458,
  -35.4745,
  -35.5026,
  -35.5299,
  -35.5552,
  -35.5809,
  -35.6062,
  -35.6316,
  -35.6576,
  -35.6841,
  -35.7109,
  -35.7377,
  -35.7641,
  -35.7899,
  -35.8151,
  -35.8398,
  -35.8643,
  -35.8886,
  -35.9128,
  -35.9372,
  -35.9618,
  -35.9864,
  -36.0108,
  -36.0345,
  -36.0574,
  -36.079,
  -36.0981,
  -36.1171,
  -36.1354,
  -36.1537,
  -36.1723,
  -36.1916,
  -36.2115,
  -36.232,
  -36.2526,
  -36.2731,
  -36.2933,
  -36.3131,
  -36.3326,
  -36.3516,
  -36.3703,
  -36.3889,
  -36.4075,
  -36.4264,
  -36.4458,
  -36.4659,
  -36.4865,
  -36.5072,
  -36.5273,
  -36.5463,
  -36.563,
  -36.5799,
  -36.5963,
  -36.6133,
  -36.6313,
  -36.6511,
  -36.673,
  -36.6978,
  -36.726,
  -36.7579,
  -36.7935,
  -36.8325,
  -36.8748,
  -36.92,
  -36.9677,
  -37.0176,
  -37.0693,
  -37.1224,
  -37.1764,
  -37.2303,
  -37.2828,
  -37.3331,
  -37.38,
  -37.4243,
  -37.4662,
  -37.5063,
  -37.5455,
  -37.5846,
  -37.6227,
  -37.6621,
  -37.7015,
  -37.7397,
  -37.7762,
  -37.8104,
  -37.842,
  -37.8709,
  -37.8974,
  -37.9222,
  -37.9461,
  -37.9703,
  -37.9952,
  -38.0215,
  -38.049,
  -38.0769,
  -38.1045,
  -38.1312,
  -38.1568,
  -38.1814,
  -38.2052,
  -38.2284,
  -38.2511,
  -38.2732,
  -38.2948,
  -38.3157,
  -38.3353,
  -38.3534,
  -38.3692,
  -38.3828,
  -38.3941,
  -38.4039,
  -38.4116,
  -38.4198,
  -38.4276,
  -38.4353,
  -38.4428,
  -38.4502,
  -38.4571,
  -38.463,
  -38.4678,
  -38.4716,
  -38.475,
  -38.4782,
  -38.4816,
  -38.4855,
  -38.4891,
  -38.4926,
  -38.4959,
  -38.4985,
  -38.5,
  -38.5002,
  -38.499,
  -38.4963,
  -38.492,
  -38.4861,
  -38.4788,
  -38.4704,
  -38.4612,
  -38.4515,
  -38.4417,
  -38.4321,
  -38.4231,
  -38.4142,
  -38.4046,
  -38.3932,
  -38.3789,
  -38.3612,
  -38.3396,
  -38.314,
  -38.2841,
  -38.25,
  -38.2116,
  -38.1669,
  -38.1159,
  -38.0551,
  -37.9814,
  -37.8928,
  -37.7879,
  -37.668,
  -37.5362,
  -37.399,
  -37.2645,
  -37.1426,
  -37.0431,
  -36.9744,
  -36.9403,
  -29.5716,
  -29.618,
  -29.6646,
  -29.7111,
  -29.7578,
  -29.8045,
  -29.8513,
  -29.8986,
  -29.9464,
  -29.9952,
  -30.0453,
  -30.0963,
  -30.1484,
  -30.2,
  -30.253,
  -30.3064,
  -30.3598,
  -30.413,
  -30.4657,
  -30.5178,
  -30.5693,
  -30.6202,
  -30.6706,
  -30.7207,
  -30.7707,
  -30.8207,
  -30.8705,
  -30.92,
  -30.9681,
  -31.017,
  -31.066,
  -31.1152,
  -31.1645,
  -31.214,
  -31.2635,
  -31.3128,
  -31.362,
  -31.4109,
  -31.4593,
  -31.5071,
  -31.5547,
  -31.6026,
  -31.651,
  -31.6999,
  -31.7478,
  -31.7968,
  -31.8453,
  -31.8936,
  -31.9421,
  -31.9905,
  -32.0392,
  -32.0881,
  -32.137,
  -32.1861,
  -32.2353,
  -32.2846,
  -32.3344,
  -32.3845,
  -32.4349,
  -32.4853,
  -32.5343,
  -32.5835,
  -32.6319,
  -32.6796,
  -32.7269,
  -32.7744,
  -32.8222,
  -32.8703,
  -32.9188,
  -32.9678,
  -33.0176,
  -33.0682,
  -33.1194,
  -33.1709,
  -33.2221,
  -33.2731,
  -33.3224,
  -33.3725,
  -33.4223,
  -33.4716,
  -33.5204,
  -33.5685,
  -33.6158,
  -33.6626,
  -33.7089,
  -33.7552,
  -33.8011,
  -33.8464,
  -33.8909,
  -33.9345,
  -33.9771,
  -34.0193,
  -34.0613,
  -34.1037,
  -34.1454,
  -34.1884,
  -34.2317,
  -34.2748,
  -34.3172,
  -34.3584,
  -34.3981,
  -34.436,
  -34.4721,
  -34.5068,
  -34.5406,
  -34.5736,
  -34.6062,
  -34.6386,
  -34.6708,
  -34.7029,
  -34.7348,
  -34.7659,
  -34.7963,
  -34.8244,
  -34.8524,
  -34.8792,
  -34.9049,
  -34.9295,
  -34.9532,
  -34.977,
  -35.0006,
  -35.0247,
  -35.0493,
  -35.0738,
  -35.0982,
  -35.1224,
  -35.1464,
  -35.1705,
  -35.1947,
  -35.2192,
  -35.2439,
  -35.2688,
  -35.2939,
  -35.3186,
  -35.3452,
  -35.373,
  -35.4014,
  -35.4299,
  -35.4577,
  -35.4845,
  -35.5104,
  -35.5357,
  -35.5606,
  -35.5855,
  -35.611,
  -35.6369,
  -35.6631,
  -35.6894,
  -35.7153,
  -35.7407,
  -35.7656,
  -35.7901,
  -35.8143,
  -35.8385,
  -35.8627,
  -35.8861,
  -35.9107,
  -35.9354,
  -35.96,
  -35.9839,
  -36.0068,
  -36.0281,
  -36.048,
  -36.0666,
  -36.0848,
  -36.103,
  -36.1217,
  -36.1412,
  -36.1614,
  -36.1821,
  -36.2028,
  -36.2232,
  -36.2432,
  -36.2629,
  -36.2821,
  -36.3011,
  -36.3198,
  -36.3382,
  -36.3557,
  -36.3743,
  -36.3936,
  -36.4136,
  -36.4343,
  -36.4553,
  -36.4756,
  -36.4951,
  -36.5134,
  -36.5306,
  -36.5476,
  -36.5651,
  -36.5837,
  -36.604,
  -36.6267,
  -36.6523,
  -36.6816,
  -36.7147,
  -36.7517,
  -36.7922,
  -36.8361,
  -36.8832,
  -36.9328,
  -36.9844,
  -37.0375,
  -37.0917,
  -37.1463,
  -37.1994,
  -37.2519,
  -37.3018,
  -37.3483,
  -37.3922,
  -37.4333,
  -37.4731,
  -37.5122,
  -37.5512,
  -37.5904,
  -37.6298,
  -37.6688,
  -37.7067,
  -37.7426,
  -37.7761,
  -37.807,
  -37.8352,
  -37.8612,
  -37.8854,
  -37.9088,
  -37.9325,
  -37.9568,
  -37.9826,
  -38.0093,
  -38.0366,
  -38.0635,
  -38.0898,
  -38.1152,
  -38.1398,
  -38.1637,
  -38.1862,
  -38.2093,
  -38.232,
  -38.2541,
  -38.2751,
  -38.2947,
  -38.3126,
  -38.3279,
  -38.3408,
  -38.3517,
  -38.3613,
  -38.37,
  -38.3783,
  -38.3861,
  -38.3936,
  -38.4008,
  -38.4076,
  -38.4139,
  -38.4191,
  -38.4232,
  -38.4262,
  -38.429,
  -38.4315,
  -38.4345,
  -38.438,
  -38.4416,
  -38.4453,
  -38.4491,
  -38.4522,
  -38.4543,
  -38.4551,
  -38.4542,
  -38.4518,
  -38.4474,
  -38.4413,
  -38.4336,
  -38.425,
  -38.4157,
  -38.4052,
  -38.396,
  -38.3871,
  -38.3789,
  -38.3709,
  -38.3623,
  -38.3519,
  -38.3386,
  -38.3217,
  -38.3007,
  -38.2755,
  -38.2457,
  -38.2116,
  -38.1731,
  -38.1291,
  -38.0778,
  -38.0167,
  -37.9435,
  -37.8554,
  -37.7513,
  -37.6315,
  -37.4999,
  -37.3618,
  -37.2259,
  -37.1019,
  -36.9995,
  -36.9271,
  -36.8903,
  -29.5506,
  -29.5975,
  -29.6448,
  -29.6921,
  -29.7394,
  -29.7866,
  -29.8335,
  -29.8806,
  -29.9282,
  -29.9758,
  -30.0256,
  -30.0765,
  -30.1281,
  -30.1802,
  -30.2325,
  -30.285,
  -30.3378,
  -30.3906,
  -30.4431,
  -30.4951,
  -30.5465,
  -30.5972,
  -30.6472,
  -30.6958,
  -30.7452,
  -30.7945,
  -30.8438,
  -30.8928,
  -30.9414,
  -30.9897,
  -31.038,
  -31.0865,
  -31.1352,
  -31.184,
  -31.233,
  -31.2825,
  -31.332,
  -31.381,
  -31.4296,
  -31.4765,
  -31.524,
  -31.5716,
  -31.6195,
  -31.6676,
  -31.716,
  -31.7644,
  -31.8129,
  -31.8615,
  -31.9104,
  -31.9594,
  -32.0086,
  -32.058,
  -32.1072,
  -32.1566,
  -32.2049,
  -32.2544,
  -32.3041,
  -32.3541,
  -32.4042,
  -32.4542,
  -32.5038,
  -32.5528,
  -32.6009,
  -32.6486,
  -32.696,
  -32.7436,
  -32.7916,
  -32.8399,
  -32.8886,
  -32.9377,
  -32.9873,
  -33.0363,
  -33.0869,
  -33.1377,
  -33.1885,
  -33.2389,
  -33.2892,
  -33.3391,
  -33.3888,
  -33.4382,
  -33.4871,
  -33.5354,
  -33.5832,
  -33.6302,
  -33.6767,
  -33.7229,
  -33.7688,
  -33.8139,
  -33.8572,
  -33.9007,
  -33.9435,
  -33.9859,
  -34.0282,
  -34.0707,
  -34.1137,
  -34.157,
  -34.2006,
  -34.2441,
  -34.2868,
  -34.3281,
  -34.3677,
  -34.4053,
  -34.4408,
  -34.4749,
  -34.508,
  -34.5404,
  -34.5726,
  -34.6036,
  -34.6356,
  -34.6676,
  -34.6993,
  -34.7304,
  -34.7606,
  -34.7897,
  -34.8177,
  -34.8446,
  -34.8703,
  -34.8949,
  -34.9189,
  -34.9423,
  -34.9654,
  -34.9889,
  -35.0127,
  -35.0365,
  -35.0602,
  -35.0837,
  -35.1072,
  -35.1297,
  -35.1534,
  -35.1774,
  -35.2016,
  -35.2262,
  -35.2512,
  -35.2767,
  -35.3032,
  -35.3307,
  -35.3589,
  -35.387,
  -35.4144,
  -35.4407,
  -35.4661,
  -35.4908,
  -35.5153,
  -35.5397,
  -35.5645,
  -35.5898,
  -35.6153,
  -35.641,
  -35.6655,
  -35.6906,
  -35.7153,
  -35.7398,
  -35.764,
  -35.788,
  -35.8124,
  -35.8369,
  -35.8615,
  -35.8861,
  -35.9106,
  -35.9345,
  -35.9573,
  -35.9785,
  -35.9981,
  -36.0166,
  -36.0347,
  -36.0531,
  -36.0721,
  -36.092,
  -36.1125,
  -36.1334,
  -36.1542,
  -36.1736,
  -36.1934,
  -36.2128,
  -36.2319,
  -36.2506,
  -36.2693,
  -36.2877,
  -36.3058,
  -36.3241,
  -36.3431,
  -36.363,
  -36.3837,
  -36.4049,
  -36.4255,
  -36.4453,
  -36.4639,
  -36.4817,
  -36.4992,
  -36.5174,
  -36.5367,
  -36.5578,
  -36.5815,
  -36.6082,
  -36.6387,
  -36.6731,
  -36.7104,
  -36.7523,
  -36.7978,
  -36.8463,
  -36.8974,
  -36.9506,
  -37.0049,
  -37.0599,
  -37.115,
  -37.1695,
  -37.2221,
  -37.2717,
  -37.318,
  -37.3613,
  -37.4019,
  -37.4412,
  -37.48,
  -37.5188,
  -37.558,
  -37.5973,
  -37.6361,
  -37.6735,
  -37.709,
  -37.742,
  -37.7723,
  -37.7999,
  -37.8252,
  -37.8489,
  -37.872,
  -37.8939,
  -37.9177,
  -37.9427,
  -37.9685,
  -37.9949,
  -38.0213,
  -38.0471,
  -38.0723,
  -38.0969,
  -38.1212,
  -38.1452,
  -38.1688,
  -38.192,
  -38.2144,
  -38.2355,
  -38.2549,
  -38.2721,
  -38.2869,
  -38.2993,
  -38.3097,
  -38.3191,
  -38.3279,
  -38.3364,
  -38.3441,
  -38.3513,
  -38.3581,
  -38.3645,
  -38.3698,
  -38.3743,
  -38.3777,
  -38.3802,
  -38.3822,
  -38.3844,
  -38.387,
  -38.3902,
  -38.3926,
  -38.3965,
  -38.4005,
  -38.4041,
  -38.4066,
  -38.4077,
  -38.4071,
  -38.4046,
  -38.4002,
  -38.394,
  -38.3862,
  -38.3773,
  -38.368,
  -38.3587,
  -38.3497,
  -38.3414,
  -38.3337,
  -38.3264,
  -38.3185,
  -38.309,
  -38.2967,
  -38.2807,
  -38.2605,
  -38.2357,
  -38.2063,
  -38.1725,
  -38.1339,
  -38.0898,
  -38.0386,
  -37.9778,
  -37.9053,
  -37.8183,
  -37.7156,
  -37.5975,
  -37.4674,
  -37.3304,
  -37.1946,
  -37.0698,
  -36.9657,
  -36.8909,
  -36.8514,
  -29.5313,
  -29.5783,
  -29.6258,
  -29.6736,
  -29.7202,
  -29.7676,
  -29.8146,
  -29.8617,
  -29.9094,
  -29.9581,
  -30.008,
  -30.0588,
  -30.1101,
  -30.1617,
  -30.2133,
  -30.265,
  -30.317,
  -30.3693,
  -30.4215,
  -30.4723,
  -30.5237,
  -30.5743,
  -30.6241,
  -30.6732,
  -30.722,
  -30.7708,
  -30.8191,
  -30.8673,
  -30.9152,
  -30.9627,
  -31.0101,
  -31.0579,
  -31.1061,
  -31.1546,
  -31.2026,
  -31.2522,
  -31.3017,
  -31.351,
  -31.3997,
  -31.4475,
  -31.4948,
  -31.5419,
  -31.5892,
  -31.6368,
  -31.6846,
  -31.7329,
  -31.7814,
  -31.8304,
  -31.8798,
  -31.9283,
  -31.9779,
  -32.0274,
  -32.0769,
  -32.1264,
  -32.1761,
  -32.2256,
  -32.2753,
  -32.3251,
  -32.3748,
  -32.4243,
  -32.4733,
  -32.5217,
  -32.5695,
  -32.6173,
  -32.6649,
  -32.7128,
  -32.7601,
  -32.8086,
  -32.8577,
  -32.9069,
  -32.9565,
  -33.0063,
  -33.0565,
  -33.1069,
  -33.1574,
  -33.2077,
  -33.258,
  -33.3079,
  -33.3576,
  -33.4068,
  -33.4557,
  -33.5041,
  -33.5519,
  -33.5983,
  -33.6449,
  -33.6908,
  -33.7361,
  -33.7807,
  -33.8247,
  -33.868,
  -33.911,
  -33.9537,
  -33.9964,
  -34.0394,
  -34.0828,
  -34.1266,
  -34.1705,
  -34.2142,
  -34.2571,
  -34.2985,
  -34.338,
  -34.3744,
  -34.4098,
  -34.4434,
  -34.4759,
  -34.5078,
  -34.5393,
  -34.5708,
  -34.6025,
  -34.6341,
  -34.6655,
  -34.6964,
  -34.7264,
  -34.7554,
  -34.7834,
  -34.8104,
  -34.8363,
  -34.8612,
  -34.885,
  -34.908,
  -34.9296,
  -34.9524,
  -34.9752,
  -34.9982,
  -35.0212,
  -35.0442,
  -35.0672,
  -35.0903,
  -35.1135,
  -35.137,
  -35.1608,
  -35.1852,
  -35.2099,
  -35.2356,
  -35.262,
  -35.2892,
  -35.317,
  -35.3447,
  -35.3714,
  -35.3972,
  -35.422,
  -35.4452,
  -35.4689,
  -35.4927,
  -35.5167,
  -35.541,
  -35.5658,
  -35.5909,
  -35.616,
  -35.641,
  -35.6656,
  -35.6902,
  -35.7145,
  -35.7388,
  -35.7632,
  -35.7878,
  -35.8126,
  -35.8372,
  -35.8615,
  -35.8853,
  -35.9077,
  -35.9286,
  -35.9481,
  -35.9657,
  -35.984,
  -36.0027,
  -36.0221,
  -36.0424,
  -36.0633,
  -36.0844,
  -36.1053,
  -36.1256,
  -36.1454,
  -36.1647,
  -36.1836,
  -36.2022,
  -36.2206,
  -36.2388,
  -36.2566,
  -36.2746,
  -36.2934,
  -36.3132,
  -36.3339,
  -36.3551,
  -36.376,
  -36.3961,
  -36.4151,
  -36.4335,
  -36.4507,
  -36.4696,
  -36.4897,
  -36.5118,
  -36.5365,
  -36.5646,
  -36.5963,
  -36.632,
  -36.6715,
  -36.7147,
  -36.7616,
  -36.8114,
  -36.8638,
  -36.9179,
  -36.9732,
  -37.029,
  -37.0846,
  -37.1392,
  -37.1918,
  -37.2413,
  -37.2875,
  -37.3301,
  -37.3704,
  -37.4092,
  -37.4477,
  -37.4864,
  -37.5255,
  -37.5646,
  -37.6021,
  -37.6393,
  -37.6744,
  -37.707,
  -37.7369,
  -37.764,
  -37.7888,
  -37.812,
  -37.8346,
  -37.8571,
  -37.8801,
  -37.9042,
  -37.9292,
  -37.9546,
  -37.9802,
  -38.0055,
  -38.0305,
  -38.0552,
  -38.0799,
  -38.1044,
  -38.1287,
  -38.1524,
  -38.1748,
  -38.1955,
  -38.2144,
  -38.2311,
  -38.2453,
  -38.2572,
  -38.2674,
  -38.2768,
  -38.2857,
  -38.2941,
  -38.301,
  -38.3078,
  -38.3143,
  -38.3199,
  -38.3244,
  -38.328,
  -38.3308,
  -38.3328,
  -38.3344,
  -38.3364,
  -38.3388,
  -38.3418,
  -38.3453,
  -38.349,
  -38.353,
  -38.3566,
  -38.3593,
  -38.3605,
  -38.3598,
  -38.3575,
  -38.353,
  -38.3468,
  -38.3391,
  -38.3302,
  -38.3209,
  -38.3117,
  -38.3029,
  -38.2948,
  -38.2873,
  -38.2802,
  -38.2726,
  -38.2637,
  -38.2521,
  -38.237,
  -38.2177,
  -38.1937,
  -38.165,
  -38.1317,
  -38.0934,
  -38.0496,
  -37.9987,
  -37.9386,
  -37.8659,
  -37.7805,
  -37.6801,
  -37.5648,
  -37.4372,
  -37.3029,
  -37.169,
  -37.045,
  -36.9405,
  -36.8641,
  -36.8213,
  -29.5125,
  -29.5596,
  -29.607,
  -29.6546,
  -29.7022,
  -29.7494,
  -29.7964,
  -29.8436,
  -29.8915,
  -29.9405,
  -29.9905,
  -30.0413,
  -30.0925,
  -30.1436,
  -30.1937,
  -30.2449,
  -30.2964,
  -30.348,
  -30.3998,
  -30.4513,
  -30.5024,
  -30.5529,
  -30.6026,
  -30.6516,
  -30.6999,
  -30.7478,
  -30.7953,
  -30.8424,
  -30.8891,
  -30.9347,
  -30.9814,
  -31.0286,
  -31.0765,
  -31.1251,
  -31.1744,
  -31.2241,
  -31.2738,
  -31.3231,
  -31.3716,
  -31.4192,
  -31.4661,
  -31.5127,
  -31.5595,
  -31.6066,
  -31.6532,
  -31.7012,
  -31.7498,
  -31.799,
  -31.8486,
  -31.8984,
  -31.9482,
  -31.9979,
  -32.0476,
  -32.0974,
  -32.1473,
  -32.197,
  -32.2467,
  -32.2962,
  -32.3454,
  -32.3941,
  -32.4413,
  -32.4891,
  -32.5368,
  -32.5845,
  -32.6325,
  -32.6809,
  -32.7296,
  -32.7787,
  -32.828,
  -32.8773,
  -32.9269,
  -32.9765,
  -33.0265,
  -33.0768,
  -33.1273,
  -33.1778,
  -33.228,
  -33.277,
  -33.3266,
  -33.3758,
  -33.4246,
  -33.473,
  -33.521,
  -33.5683,
  -33.6149,
  -33.6607,
  -33.7055,
  -33.7496,
  -33.7931,
  -33.8362,
  -33.8791,
  -33.922,
  -33.9652,
  -34.0088,
  -34.0528,
  -34.096,
  -34.1402,
  -34.1841,
  -34.2271,
  -34.2686,
  -34.3082,
  -34.3455,
  -34.3807,
  -34.414,
  -34.4461,
  -34.4774,
  -34.5083,
  -34.5392,
  -34.5703,
  -34.6015,
  -34.6325,
  -34.6629,
  -34.6926,
  -34.7213,
  -34.7481,
  -34.7751,
  -34.801,
  -34.8259,
  -34.8495,
  -34.8723,
  -34.8945,
  -34.9165,
  -34.9386,
  -34.9609,
  -34.9833,
  -35.0059,
  -35.0285,
  -35.0512,
  -35.074,
  -35.0972,
  -35.1207,
  -35.1449,
  -35.1697,
  -35.1953,
  -35.2207,
  -35.2478,
  -35.2752,
  -35.3022,
  -35.3283,
  -35.3533,
  -35.3773,
  -35.4004,
  -35.4232,
  -35.4458,
  -35.4687,
  -35.4921,
  -35.5161,
  -35.5406,
  -35.5656,
  -35.5906,
  -35.6155,
  -35.6404,
  -35.6651,
  -35.6898,
  -35.7145,
  -35.7394,
  -35.7632,
  -35.7877,
  -35.8117,
  -35.835,
  -35.857,
  -35.8776,
  -35.897,
  -35.9158,
  -35.9344,
  -35.9536,
  -35.9734,
  -35.994,
  -36.0151,
  -36.0364,
  -36.0573,
  -36.0778,
  -36.0975,
  -36.1168,
  -36.1356,
  -36.1542,
  -36.1725,
  -36.1904,
  -36.2081,
  -36.226,
  -36.2437,
  -36.2634,
  -36.2841,
  -36.3053,
  -36.3263,
  -36.3466,
  -36.3661,
  -36.3849,
  -36.4038,
  -36.4234,
  -36.4444,
  -36.4675,
  -36.4936,
  -36.523,
  -36.5561,
  -36.5933,
  -36.6342,
  -36.6787,
  -36.7267,
  -36.7776,
  -36.8309,
  -36.8859,
  -36.9417,
  -36.9978,
  -37.0534,
  -37.1078,
  -37.159,
  -37.2082,
  -37.254,
  -37.2966,
  -37.3368,
  -37.3756,
  -37.4141,
  -37.4529,
  -37.492,
  -37.5311,
  -37.5694,
  -37.6063,
  -37.6411,
  -37.6734,
  -37.7028,
  -37.7295,
  -37.7538,
  -37.7765,
  -37.7985,
  -37.8203,
  -37.8427,
  -37.8659,
  -37.8899,
  -37.9144,
  -37.9393,
  -37.9641,
  -37.9889,
  -38.0139,
  -38.0389,
  -38.0639,
  -38.0885,
  -38.1113,
  -38.1335,
  -38.1539,
  -38.1723,
  -38.1885,
  -38.2024,
  -38.2141,
  -38.2243,
  -38.2336,
  -38.2424,
  -38.2506,
  -38.2582,
  -38.2648,
  -38.2705,
  -38.2753,
  -38.2792,
  -38.2821,
  -38.2843,
  -38.286,
  -38.2876,
  -38.2895,
  -38.292,
  -38.2949,
  -38.2984,
  -38.3021,
  -38.3058,
  -38.3092,
  -38.3118,
  -38.3129,
  -38.3123,
  -38.31,
  -38.3057,
  -38.2997,
  -38.2921,
  -38.2833,
  -38.2739,
  -38.2646,
  -38.2558,
  -38.2466,
  -38.2391,
  -38.2319,
  -38.2244,
  -38.2156,
  -38.2047,
  -38.1904,
  -38.1719,
  -38.1489,
  -38.1211,
  -38.0886,
  -38.0511,
  -38.0079,
  -37.9576,
  -37.8985,
  -37.8283,
  -37.745,
  -37.6474,
  -37.5358,
  -37.4123,
  -37.2819,
  -37.1515,
  -37.0299,
  -36.9263,
  -36.849,
  -36.8036,
  -29.4961,
  -29.543,
  -29.5902,
  -29.6374,
  -29.6844,
  -29.7313,
  -29.7782,
  -29.8256,
  -29.8739,
  -29.9232,
  -29.9724,
  -30.0232,
  -30.0741,
  -30.125,
  -30.1757,
  -30.2266,
  -30.2776,
  -30.3287,
  -30.3799,
  -30.4309,
  -30.4818,
  -30.5322,
  -30.582,
  -30.631,
  -30.6777,
  -30.7248,
  -30.771,
  -30.8168,
  -30.8623,
  -30.9077,
  -30.9537,
  -31.0006,
  -31.0486,
  -31.0977,
  -31.1475,
  -31.1976,
  -31.2474,
  -31.2965,
  -31.3446,
  -31.3907,
  -31.4369,
  -31.4829,
  -31.5291,
  -31.5759,
  -31.6232,
  -31.6713,
  -31.7201,
  -31.7695,
  -31.819,
  -31.8688,
  -31.9186,
  -31.9683,
  -32.0181,
  -32.0681,
  -32.1182,
  -32.1671,
  -32.2168,
  -32.266,
  -32.3146,
  -32.3625,
  -32.41,
  -32.4572,
  -32.5047,
  -32.5527,
  -32.6012,
  -32.65,
  -32.6991,
  -32.7484,
  -32.7979,
  -32.8474,
  -32.8968,
  -32.9463,
  -32.9952,
  -33.0456,
  -33.0965,
  -33.1474,
  -33.1978,
  -33.2479,
  -33.2975,
  -33.3467,
  -33.3955,
  -33.4439,
  -33.4919,
  -33.5394,
  -33.586,
  -33.6317,
  -33.6763,
  -33.7199,
  -33.7628,
  -33.8045,
  -33.8472,
  -33.8903,
  -33.9339,
  -33.978,
  -34.0224,
  -34.067,
  -34.1115,
  -34.1555,
  -34.1985,
  -34.2401,
  -34.2798,
  -34.3172,
  -34.3525,
  -34.3856,
  -34.4173,
  -34.448,
  -34.4782,
  -34.5085,
  -34.538,
  -34.5686,
  -34.599,
  -34.629,
  -34.6581,
  -34.6864,
  -34.7138,
  -34.7404,
  -34.7662,
  -34.7909,
  -34.8144,
  -34.837,
  -34.8588,
  -34.8804,
  -34.902,
  -34.9236,
  -34.9456,
  -34.9677,
  -34.9899,
  -35.0123,
  -35.0339,
  -35.0567,
  -35.08,
  -35.1039,
  -35.1287,
  -35.1543,
  -35.1807,
  -35.2076,
  -35.2344,
  -35.2609,
  -35.2863,
  -35.3104,
  -35.3334,
  -35.3555,
  -35.3769,
  -35.3982,
  -35.4198,
  -35.442,
  -35.4651,
  -35.4892,
  -35.5141,
  -35.5384,
  -35.5638,
  -35.5892,
  -35.6144,
  -35.6396,
  -35.6648,
  -35.6901,
  -35.715,
  -35.7393,
  -35.7628,
  -35.7853,
  -35.8067,
  -35.827,
  -35.8465,
  -35.8654,
  -35.8845,
  -35.904,
  -35.9243,
  -35.9451,
  -35.9663,
  -35.9876,
  -36.0086,
  -36.0292,
  -36.0483,
  -36.0677,
  -36.0867,
  -36.1054,
  -36.1236,
  -36.1415,
  -36.1591,
  -36.1771,
  -36.1956,
  -36.2156,
  -36.2364,
  -36.2576,
  -36.2786,
  -36.2991,
  -36.3189,
  -36.3383,
  -36.3577,
  -36.378,
  -36.3998,
  -36.4239,
  -36.4511,
  -36.4819,
  -36.5166,
  -36.5551,
  -36.5976,
  -36.6434,
  -36.6915,
  -36.7433,
  -36.7973,
  -36.8527,
  -36.9088,
  -36.9648,
  -37.0201,
  -37.0739,
  -37.1254,
  -37.1739,
  -37.2195,
  -37.2623,
  -37.3027,
  -37.342,
  -37.3811,
  -37.4203,
  -37.4597,
  -37.4987,
  -37.5368,
  -37.5734,
  -37.6079,
  -37.6397,
  -37.6689,
  -37.6952,
  -37.7191,
  -37.7414,
  -37.7628,
  -37.7842,
  -37.8059,
  -37.8272,
  -37.8502,
  -37.8738,
  -37.8979,
  -37.9222,
  -37.9469,
  -37.9719,
  -37.9971,
  -38.0223,
  -38.047,
  -38.0704,
  -38.0922,
  -38.1121,
  -38.1298,
  -38.1459,
  -38.1598,
  -38.1717,
  -38.182,
  -38.1912,
  -38.1998,
  -38.2077,
  -38.215,
  -38.2211,
  -38.2263,
  -38.2305,
  -38.2335,
  -38.236,
  -38.2379,
  -38.2395,
  -38.2412,
  -38.2432,
  -38.2457,
  -38.2488,
  -38.2522,
  -38.2556,
  -38.2581,
  -38.2611,
  -38.2633,
  -38.2643,
  -38.2638,
  -38.2616,
  -38.2577,
  -38.2519,
  -38.2446,
  -38.2359,
  -38.2265,
  -38.2171,
  -38.208,
  -38.1996,
  -38.1918,
  -38.1843,
  -38.1765,
  -38.1678,
  -38.1571,
  -38.1433,
  -38.1256,
  -38.1037,
  -38.0771,
  -38.0457,
  -38.0093,
  -37.9671,
  -37.918,
  -37.8602,
  -37.7918,
  -37.711,
  -37.6169,
  -37.5095,
  -37.391,
  -37.2657,
  -37.1402,
  -37.0226,
  -36.9211,
  -36.8437,
  -36.7964,
  -29.4805,
  -29.5274,
  -29.5744,
  -29.621,
  -29.6673,
  -29.7127,
  -29.7594,
  -29.807,
  -29.8556,
  -29.9053,
  -29.9557,
  -30.0065,
  -30.0573,
  -30.108,
  -30.1585,
  -30.2091,
  -30.2597,
  -30.3103,
  -30.3609,
  -30.4114,
  -30.4608,
  -30.5111,
  -30.5608,
  -30.6094,
  -30.6569,
  -30.7027,
  -30.7478,
  -30.7922,
  -30.8364,
  -30.8808,
  -30.9263,
  -30.9732,
  -31.0217,
  -31.0716,
  -31.1222,
  -31.1719,
  -31.2216,
  -31.2703,
  -31.3179,
  -31.3641,
  -31.4095,
  -31.4547,
  -31.5004,
  -31.5467,
  -31.5939,
  -31.642,
  -31.691,
  -31.7402,
  -31.7898,
  -31.8394,
  -31.888,
  -31.9377,
  -31.9875,
  -32.0376,
  -32.0877,
  -32.1377,
  -32.1874,
  -32.2364,
  -32.2846,
  -32.3319,
  -32.3787,
  -32.4256,
  -32.473,
  -32.5213,
  -32.5702,
  -32.6194,
  -32.6689,
  -32.7174,
  -32.7669,
  -32.8162,
  -32.8653,
  -32.9146,
  -32.9643,
  -33.015,
  -33.0661,
  -33.1174,
  -33.1685,
  -33.2189,
  -33.2687,
  -33.318,
  -33.3669,
  -33.4154,
  -33.4636,
  -33.5112,
  -33.5572,
  -33.6029,
  -33.6474,
  -33.6907,
  -33.7333,
  -33.7755,
  -33.818,
  -33.8611,
  -33.9048,
  -33.9492,
  -33.9939,
  -34.0387,
  -34.0832,
  -34.1272,
  -34.1702,
  -34.2117,
  -34.2514,
  -34.289,
  -34.3233,
  -34.3564,
  -34.3878,
  -34.4181,
  -34.4478,
  -34.4775,
  -34.5076,
  -34.5376,
  -34.5675,
  -34.5969,
  -34.6254,
  -34.6531,
  -34.68,
  -34.7059,
  -34.7312,
  -34.7552,
  -34.7786,
  -34.8012,
  -34.8229,
  -34.8432,
  -34.8644,
  -34.8857,
  -34.9072,
  -34.9289,
  -34.9508,
  -34.9728,
  -34.9948,
  -35.0173,
  -35.0403,
  -35.0641,
  -35.0889,
  -35.1145,
  -35.1407,
  -35.1673,
  -35.1936,
  -35.2194,
  -35.244,
  -35.2672,
  -35.2892,
  -35.3101,
  -35.3292,
  -35.349,
  -35.3691,
  -35.39,
  -35.4123,
  -35.436,
  -35.4609,
  -35.4865,
  -35.5125,
  -35.5386,
  -35.5644,
  -35.5901,
  -35.6159,
  -35.6415,
  -35.6665,
  -35.6905,
  -35.7135,
  -35.7353,
  -35.7561,
  -35.7761,
  -35.7954,
  -35.8145,
  -35.8329,
  -35.8528,
  -35.8734,
  -35.8944,
  -35.9157,
  -35.9371,
  -35.9582,
  -35.9788,
  -35.9992,
  -36.0191,
  -36.0385,
  -36.0573,
  -36.0756,
  -36.0937,
  -36.1116,
  -36.1298,
  -36.1489,
  -36.169,
  -36.1899,
  -36.2112,
  -36.2323,
  -36.2528,
  -36.2728,
  -36.2925,
  -36.3125,
  -36.3323,
  -36.3547,
  -36.3797,
  -36.408,
  -36.4402,
  -36.4763,
  -36.5164,
  -36.5602,
  -36.6074,
  -36.6576,
  -36.7102,
  -36.7646,
  -36.8201,
  -36.8761,
  -36.9317,
  -36.9862,
  -37.039,
  -37.0898,
  -37.1378,
  -37.1832,
  -37.2262,
  -37.2672,
  -37.3076,
  -37.3477,
  -37.3877,
  -37.4275,
  -37.4667,
  -37.5046,
  -37.5398,
  -37.5739,
  -37.6055,
  -37.6342,
  -37.66,
  -37.6836,
  -37.7055,
  -37.7264,
  -37.7472,
  -37.7683,
  -37.7897,
  -37.8118,
  -37.8344,
  -37.8578,
  -37.8816,
  -37.9061,
  -37.9311,
  -37.9563,
  -37.9813,
  -38.0056,
  -38.0285,
  -38.0495,
  -38.0688,
  -38.0866,
  -38.1024,
  -38.1166,
  -38.1289,
  -38.1395,
  -38.1488,
  -38.1571,
  -38.1646,
  -38.1713,
  -38.1771,
  -38.1806,
  -38.184,
  -38.1867,
  -38.1887,
  -38.1904,
  -38.1922,
  -38.1942,
  -38.1964,
  -38.1991,
  -38.2022,
  -38.2055,
  -38.2087,
  -38.2118,
  -38.2143,
  -38.2161,
  -38.2169,
  -38.2164,
  -38.2144,
  -38.211,
  -38.2057,
  -38.1986,
  -38.1902,
  -38.1808,
  -38.1713,
  -38.162,
  -38.1533,
  -38.1453,
  -38.1374,
  -38.1293,
  -38.1203,
  -38.1096,
  -38.0962,
  -38.0793,
  -38.0583,
  -38.033,
  -38.0029,
  -37.9678,
  -37.927,
  -37.8793,
  -37.8233,
  -37.7571,
  -37.6794,
  -37.5881,
  -37.4856,
  -37.3729,
  -37.2539,
  -37.1343,
  -37.0216,
  -36.9234,
  -36.8469,
  -36.7979,
  -29.4654,
  -29.5113,
  -29.5578,
  -29.6039,
  -29.6498,
  -29.6958,
  -29.7424,
  -29.7901,
  -29.839,
  -29.889,
  -29.9396,
  -29.9905,
  -30.0413,
  -30.092,
  -30.1424,
  -30.1916,
  -30.2418,
  -30.2919,
  -30.3418,
  -30.3916,
  -30.4416,
  -30.4915,
  -30.5408,
  -30.5889,
  -30.6354,
  -30.6803,
  -30.7241,
  -30.7673,
  -30.8104,
  -30.8542,
  -30.8985,
  -30.9457,
  -30.995,
  -31.0457,
  -31.0971,
  -31.1482,
  -31.198,
  -31.2464,
  -31.293,
  -31.3384,
  -31.3829,
  -31.4273,
  -31.4723,
  -31.5183,
  -31.5654,
  -31.6125,
  -31.6614,
  -31.7106,
  -31.76,
  -31.8094,
  -31.8588,
  -31.9084,
  -31.9582,
  -32.0081,
  -32.0582,
  -32.1081,
  -32.1577,
  -32.2066,
  -32.2545,
  -32.3016,
  -32.3482,
  -32.3939,
  -32.4413,
  -32.4897,
  -32.5389,
  -32.5884,
  -32.638,
  -32.6876,
  -32.7369,
  -32.7858,
  -32.8346,
  -32.8835,
  -32.9331,
  -32.9838,
  -33.0353,
  -33.087,
  -33.1385,
  -33.1894,
  -33.2386,
  -33.2882,
  -33.3375,
  -33.3863,
  -33.4349,
  -33.4829,
  -33.5301,
  -33.5761,
  -33.6207,
  -33.664,
  -33.7064,
  -33.7483,
  -33.7905,
  -33.8334,
  -33.8772,
  -33.9215,
  -33.9663,
  -34.011,
  -34.0544,
  -34.0982,
  -34.1409,
  -34.1822,
  -34.2218,
  -34.2594,
  -34.2948,
  -34.328,
  -34.3594,
  -34.3894,
  -34.4189,
  -34.4483,
  -34.478,
  -34.5077,
  -34.5371,
  -34.566,
  -34.594,
  -34.621,
  -34.6471,
  -34.6714,
  -34.6957,
  -34.7192,
  -34.7419,
  -34.7641,
  -34.7857,
  -34.8071,
  -34.8282,
  -34.8493,
  -34.8704,
  -34.8916,
  -34.913,
  -34.9344,
  -34.956,
  -34.9779,
  -35.0006,
  -35.0242,
  -35.0489,
  -35.0744,
  -35.1003,
  -35.1254,
  -35.151,
  -35.176,
  -35.1998,
  -35.2223,
  -35.2434,
  -35.2633,
  -35.2821,
  -35.3006,
  -35.3193,
  -35.3391,
  -35.3604,
  -35.3836,
  -35.4085,
  -35.4343,
  -35.4606,
  -35.4871,
  -35.5136,
  -35.54,
  -35.5663,
  -35.5921,
  -35.6171,
  -35.6398,
  -35.6623,
  -35.6835,
  -35.7038,
  -35.7235,
  -35.7427,
  -35.762,
  -35.7816,
  -35.8018,
  -35.8226,
  -35.8438,
  -35.8652,
  -35.8867,
  -35.908,
  -35.9291,
  -35.9497,
  -35.97,
  -35.9898,
  -36.009,
  -36.0275,
  -36.0458,
  -36.0642,
  -36.0831,
  -36.1029,
  -36.1225,
  -36.1437,
  -36.1651,
  -36.1861,
  -36.2066,
  -36.2267,
  -36.2466,
  -36.2669,
  -36.2882,
  -36.3112,
  -36.337,
  -36.3662,
  -36.3995,
  -36.437,
  -36.4786,
  -36.5238,
  -36.5723,
  -36.6234,
  -36.6767,
  -36.7314,
  -36.7869,
  -36.8424,
  -36.8973,
  -36.951,
  -37.0028,
  -37.0526,
  -37.1002,
  -37.1446,
  -37.1882,
  -37.2304,
  -37.2719,
  -37.3131,
  -37.3541,
  -37.3945,
  -37.4339,
  -37.4719,
  -37.5079,
  -37.5416,
  -37.5727,
  -37.6009,
  -37.6263,
  -37.6494,
  -37.6709,
  -37.6914,
  -37.7115,
  -37.7317,
  -37.7523,
  -37.7734,
  -37.7953,
  -37.8179,
  -37.8414,
  -37.8656,
  -37.8904,
  -37.9154,
  -37.94,
  -37.9635,
  -37.9856,
  -38.006,
  -38.0239,
  -38.0415,
  -38.0576,
  -38.0722,
  -38.0849,
  -38.0958,
  -38.1051,
  -38.1131,
  -38.1203,
  -38.1265,
  -38.1315,
  -38.1355,
  -38.1383,
  -38.1404,
  -38.1422,
  -38.144,
  -38.146,
  -38.1483,
  -38.1508,
  -38.1537,
  -38.1568,
  -38.16,
  -38.163,
  -38.1656,
  -38.1677,
  -38.1691,
  -38.1696,
  -38.169,
  -38.1673,
  -38.1643,
  -38.1595,
  -38.153,
  -38.1449,
  -38.1358,
  -38.1263,
  -38.117,
  -38.1083,
  -38.1,
  -38.091,
  -38.0825,
  -38.0732,
  -38.0622,
  -38.049,
  -38.0326,
  -38.0125,
  -37.9883,
  -37.9597,
  -37.9261,
  -37.8869,
  -37.841,
  -37.7871,
  -37.7236,
  -37.6493,
  -37.5635,
  -37.4666,
  -37.3604,
  -37.2484,
  -37.1357,
  -37.0289,
  -36.9347,
  -36.8596,
  -36.8087,
  -29.4492,
  -29.4961,
  -29.5424,
  -29.5882,
  -29.6338,
  -29.6797,
  -29.7263,
  -29.7742,
  -29.8233,
  -29.8734,
  -29.9232,
  -29.9743,
  -30.0252,
  -30.0759,
  -30.1262,
  -30.1762,
  -30.2259,
  -30.2753,
  -30.3245,
  -30.3738,
  -30.4232,
  -30.4724,
  -30.521,
  -30.5681,
  -30.6136,
  -30.6564,
  -30.699,
  -30.7411,
  -30.7835,
  -30.827,
  -30.8724,
  -30.9202,
  -30.9703,
  -31.0221,
  -31.0743,
  -31.1257,
  -31.1754,
  -31.2232,
  -31.2691,
  -31.3135,
  -31.3561,
  -31.3998,
  -31.4441,
  -31.4897,
  -31.5366,
  -31.5848,
  -31.6337,
  -31.6829,
  -31.7321,
  -31.7813,
  -31.8306,
  -31.88,
  -31.9295,
  -31.9791,
  -32.0288,
  -32.0784,
  -32.1269,
  -32.1759,
  -32.2239,
  -32.2711,
  -32.3177,
  -32.3644,
  -32.4119,
  -32.4603,
  -32.5095,
  -32.5591,
  -32.6087,
  -32.6583,
  -32.7072,
  -32.7557,
  -32.8038,
  -32.8523,
  -32.9018,
  -32.9515,
  -33.0031,
  -33.0552,
  -33.107,
  -33.1583,
  -33.209,
  -33.2592,
  -33.3089,
  -33.3584,
  -33.4074,
  -33.4559,
  -33.5035,
  -33.5499,
  -33.5949,
  -33.6384,
  -33.6809,
  -33.7227,
  -33.7636,
  -33.8064,
  -33.8499,
  -33.8942,
  -33.9388,
  -33.9833,
  -34.0274,
  -34.0708,
  -34.113,
  -34.1539,
  -34.1932,
  -34.2307,
  -34.2662,
  -34.2996,
  -34.331,
  -34.3611,
  -34.3905,
  -34.4198,
  -34.4492,
  -34.4778,
  -34.5069,
  -34.5354,
  -34.5629,
  -34.5894,
  -34.6147,
  -34.6389,
  -34.662,
  -34.6845,
  -34.7065,
  -34.7284,
  -34.7499,
  -34.7715,
  -34.7927,
  -34.8138,
  -34.8346,
  -34.8553,
  -34.8761,
  -34.8967,
  -34.9175,
  -34.9377,
  -34.9599,
  -34.9832,
  -35.0076,
  -35.0328,
  -35.0582,
  -35.0834,
  -35.1083,
  -35.1323,
  -35.1554,
  -35.1772,
  -35.1976,
  -35.2168,
  -35.2348,
  -35.2522,
  -35.27,
  -35.2887,
  -35.3092,
  -35.3318,
  -35.3562,
  -35.382,
  -35.4074,
  -35.4341,
  -35.4611,
  -35.4879,
  -35.5144,
  -35.5404,
  -35.5653,
  -35.5887,
  -35.6108,
  -35.6318,
  -35.6518,
  -35.6712,
  -35.6905,
  -35.7099,
  -35.7298,
  -35.7503,
  -35.7712,
  -35.7925,
  -35.8141,
  -35.8358,
  -35.8574,
  -35.8788,
  -35.8999,
  -35.9196,
  -35.9398,
  -35.9593,
  -35.9782,
  -35.9968,
  -36.0158,
  -36.0357,
  -36.0564,
  -36.0778,
  -36.0993,
  -36.1207,
  -36.1417,
  -36.1621,
  -36.1823,
  -36.2024,
  -36.2229,
  -36.2446,
  -36.2682,
  -36.2947,
  -36.3248,
  -36.3591,
  -36.3977,
  -36.4406,
  -36.4871,
  -36.5367,
  -36.5889,
  -36.6418,
  -36.6968,
  -36.7521,
  -36.8071,
  -36.8612,
  -36.9138,
  -36.9647,
  -37.0138,
  -37.0611,
  -37.1067,
  -37.151,
  -37.1943,
  -37.2369,
  -37.2792,
  -37.3211,
  -37.3621,
  -37.402,
  -37.4402,
  -37.4761,
  -37.5095,
  -37.54,
  -37.5677,
  -37.5926,
  -37.6152,
  -37.6364,
  -37.6564,
  -37.6759,
  -37.6953,
  -37.715,
  -37.7342,
  -37.7554,
  -37.7775,
  -37.8006,
  -37.8246,
  -37.8491,
  -37.8736,
  -37.8973,
  -37.9199,
  -37.9412,
  -37.9608,
  -37.9794,
  -37.997,
  -38.0134,
  -38.0284,
  -38.0414,
  -38.0525,
  -38.0618,
  -38.0697,
  -38.0765,
  -38.0823,
  -38.0868,
  -38.0902,
  -38.0925,
  -38.0942,
  -38.0959,
  -38.0976,
  -38.0998,
  -38.1022,
  -38.1049,
  -38.1079,
  -38.1109,
  -38.1139,
  -38.1167,
  -38.1192,
  -38.1209,
  -38.121,
  -38.1213,
  -38.1207,
  -38.1192,
  -38.1165,
  -38.1123,
  -38.1064,
  -38.0989,
  -38.0902,
  -38.0809,
  -38.0719,
  -38.0635,
  -38.0553,
  -38.0472,
  -38.0385,
  -38.0289,
  -38.0175,
  -38.0043,
  -37.9881,
  -37.9685,
  -37.9453,
  -37.9181,
  -37.8862,
  -37.849,
  -37.8052,
  -37.7538,
  -37.6935,
  -37.6232,
  -37.5424,
  -37.4515,
  -37.3523,
  -37.248,
  -37.1429,
  -37.0424,
  -36.9531,
  -36.88,
  -36.8277,
  -29.434,
  -29.4805,
  -29.5267,
  -29.5723,
  -29.6178,
  -29.6638,
  -29.7097,
  -29.7579,
  -29.8072,
  -29.8576,
  -29.9086,
  -29.9598,
  -30.0109,
  -30.0616,
  -30.1117,
  -30.1613,
  -30.2105,
  -30.2594,
  -30.3081,
  -30.3568,
  -30.4045,
  -30.4528,
  -30.5003,
  -30.5461,
  -30.5903,
  -30.633,
  -30.6746,
  -30.7161,
  -30.7581,
  -30.8016,
  -30.8473,
  -30.8956,
  -30.9464,
  -30.9987,
  -31.0514,
  -31.102,
  -31.1516,
  -31.1989,
  -31.2442,
  -31.288,
  -31.3309,
  -31.3739,
  -31.4178,
  -31.4629,
  -31.5096,
  -31.5577,
  -31.6065,
  -31.6557,
  -31.705,
  -31.7542,
  -31.8035,
  -31.8517,
  -31.9009,
  -31.9501,
  -31.9993,
  -32.0486,
  -32.0979,
  -32.1468,
  -32.1949,
  -32.2423,
  -32.2891,
  -32.3359,
  -32.3834,
  -32.4317,
  -32.4807,
  -32.5302,
  -32.5799,
  -32.628,
  -32.6768,
  -32.7246,
  -32.7726,
  -32.8206,
  -32.8699,
  -32.9205,
  -32.9721,
  -33.0243,
  -33.0764,
  -33.1281,
  -33.1794,
  -33.2303,
  -33.2806,
  -33.3306,
  -33.3802,
  -33.4292,
  -33.4772,
  -33.523,
  -33.5683,
  -33.6122,
  -33.6549,
  -33.6971,
  -33.739,
  -33.7816,
  -33.825,
  -33.8691,
  -33.9136,
  -33.9578,
  -34.0015,
  -34.0444,
  -34.0861,
  -34.1265,
  -34.1654,
  -34.2027,
  -34.2383,
  -34.2708,
  -34.3025,
  -34.3327,
  -34.3623,
  -34.3916,
  -34.421,
  -34.4503,
  -34.4792,
  -34.5073,
  -34.5344,
  -34.5603,
  -34.5849,
  -34.6083,
  -34.6304,
  -34.652,
  -34.6734,
  -34.6947,
  -34.7161,
  -34.7373,
  -34.7574,
  -34.7782,
  -34.7987,
  -34.8188,
  -34.8388,
  -34.8585,
  -34.8784,
  -34.8989,
  -34.9204,
  -34.943,
  -34.9668,
  -34.9913,
  -35.0159,
  -35.0404,
  -35.0643,
  -35.0875,
  -35.1098,
  -35.1311,
  -35.1512,
  -35.1698,
  -35.1874,
  -35.2034,
  -35.2204,
  -35.2383,
  -35.2579,
  -35.2796,
  -35.3033,
  -35.3285,
  -35.3546,
  -35.3811,
  -35.4079,
  -35.435,
  -35.4618,
  -35.4878,
  -35.5126,
  -35.536,
  -35.558,
  -35.579,
  -35.599,
  -35.6186,
  -35.6381,
  -35.6577,
  -35.6779,
  -35.6985,
  -35.7187,
  -35.7401,
  -35.762,
  -35.7841,
  -35.8061,
  -35.8278,
  -35.8493,
  -35.8705,
  -35.8912,
  -35.9111,
  -35.9304,
  -35.9495,
  -35.9692,
  -35.9898,
  -36.0112,
  -36.0331,
  -36.055,
  -36.0763,
  -36.0972,
  -36.1176,
  -36.1378,
  -36.1581,
  -36.1791,
  -36.2012,
  -36.2244,
  -36.2516,
  -36.2827,
  -36.318,
  -36.3575,
  -36.4013,
  -36.4489,
  -36.4995,
  -36.5526,
  -36.6073,
  -36.6626,
  -36.718,
  -36.7726,
  -36.8261,
  -36.8781,
  -36.9284,
  -36.9771,
  -37.0243,
  -37.0701,
  -37.1149,
  -37.1588,
  -37.2021,
  -37.2451,
  -37.2874,
  -37.3289,
  -37.3692,
  -37.4076,
  -37.4438,
  -37.4771,
  -37.5064,
  -37.5336,
  -37.5583,
  -37.5807,
  -37.6016,
  -37.6212,
  -37.6399,
  -37.6586,
  -37.6775,
  -37.697,
  -37.7175,
  -37.7393,
  -37.7621,
  -37.7857,
  -37.8097,
  -37.8334,
  -37.8563,
  -37.878,
  -37.8984,
  -37.9175,
  -37.9357,
  -37.9529,
  -37.9691,
  -37.9841,
  -37.9973,
  -38.0085,
  -38.0179,
  -38.0257,
  -38.0323,
  -38.0376,
  -38.0417,
  -38.0446,
  -38.0464,
  -38.0467,
  -38.048,
  -38.0496,
  -38.0517,
  -38.0543,
  -38.0571,
  -38.0601,
  -38.0632,
  -38.0665,
  -38.0691,
  -38.0714,
  -38.0729,
  -38.0738,
  -38.0739,
  -38.0732,
  -38.0717,
  -38.0695,
  -38.0659,
  -38.0609,
  -38.0544,
  -38.0465,
  -38.0381,
  -38.0294,
  -38.0211,
  -38.0129,
  -38.0046,
  -37.9956,
  -37.9856,
  -37.9739,
  -37.9604,
  -37.9444,
  -37.9252,
  -37.9029,
  -37.877,
  -37.8468,
  -37.8114,
  -37.7699,
  -37.7212,
  -37.6644,
  -37.5984,
  -37.523,
  -37.4385,
  -37.3467,
  -37.2492,
  -37.1518,
  -37.0583,
  -36.974,
  -36.9032,
  -36.8508,
  -29.4193,
  -29.4644,
  -29.5102,
  -29.5558,
  -29.6015,
  -29.6478,
  -29.695,
  -29.7435,
  -29.793,
  -29.8435,
  -29.8945,
  -29.9458,
  -29.9968,
  -30.0474,
  -30.0973,
  -30.1466,
  -30.1945,
  -30.243,
  -30.2912,
  -30.3393,
  -30.3872,
  -30.4344,
  -30.4805,
  -30.525,
  -30.568,
  -30.6096,
  -30.6505,
  -30.6915,
  -30.7334,
  -30.777,
  -30.8231,
  -30.8709,
  -30.9222,
  -30.975,
  -31.0279,
  -31.0795,
  -31.129,
  -31.176,
  -31.2208,
  -31.2641,
  -31.3067,
  -31.3492,
  -31.3927,
  -31.4375,
  -31.4839,
  -31.5319,
  -31.5798,
  -31.629,
  -31.6785,
  -31.7279,
  -31.7772,
  -31.8262,
  -31.875,
  -31.9236,
  -31.9722,
  -32.0209,
  -32.0698,
  -32.1187,
  -32.1669,
  -32.2145,
  -32.2615,
  -32.3085,
  -32.3549,
  -32.403,
  -32.4518,
  -32.501,
  -32.5503,
  -32.5993,
  -32.6476,
  -32.6954,
  -32.743,
  -32.791,
  -32.8401,
  -32.8903,
  -32.9419,
  -32.9941,
  -33.0464,
  -33.0985,
  -33.1503,
  -33.2007,
  -33.2517,
  -33.3024,
  -33.3525,
  -33.4019,
  -33.4502,
  -33.4973,
  -33.543,
  -33.5873,
  -33.6306,
  -33.6732,
  -33.7156,
  -33.7584,
  -33.8018,
  -33.8458,
  -33.89,
  -33.9339,
  -33.9772,
  -34.0185,
  -34.0596,
  -34.0995,
  -34.138,
  -34.1752,
  -34.2107,
  -34.2444,
  -34.2763,
  -34.3069,
  -34.3367,
  -34.3661,
  -34.3954,
  -34.4245,
  -34.453,
  -34.4807,
  -34.5074,
  -34.5327,
  -34.5567,
  -34.5794,
  -34.5999,
  -34.6208,
  -34.6414,
  -34.6621,
  -34.6829,
  -34.7037,
  -34.7244,
  -34.7447,
  -34.7646,
  -34.7841,
  -34.8032,
  -34.8222,
  -34.8412,
  -34.8608,
  -34.8813,
  -34.9031,
  -34.9259,
  -34.9494,
  -34.9729,
  -34.9963,
  -35.0183,
  -35.0407,
  -35.0624,
  -35.0832,
  -35.103,
  -35.1216,
  -35.139,
  -35.1558,
  -35.1724,
  -35.1898,
  -35.2087,
  -35.2294,
  -35.252,
  -35.2762,
  -35.3015,
  -35.3275,
  -35.3541,
  -35.381,
  -35.4077,
  -35.4338,
  -35.4586,
  -35.482,
  -35.5033,
  -35.5245,
  -35.5449,
  -35.5648,
  -35.5846,
  -35.6047,
  -35.6251,
  -35.6459,
  -35.6671,
  -35.6888,
  -35.711,
  -35.7334,
  -35.7559,
  -35.7781,
  -35.8001,
  -35.8217,
  -35.8428,
  -35.8631,
  -35.8828,
  -35.9025,
  -35.9227,
  -35.9439,
  -35.9659,
  -35.9882,
  -36.0092,
  -36.0306,
  -36.0514,
  -36.0718,
  -36.0923,
  -36.113,
  -36.1345,
  -36.1572,
  -36.1821,
  -36.2101,
  -36.2417,
  -36.2777,
  -36.3184,
  -36.3631,
  -36.4117,
  -36.4635,
  -36.5174,
  -36.5727,
  -36.6284,
  -36.6839,
  -36.7385,
  -36.7917,
  -36.8434,
  -36.8933,
  -36.9417,
  -36.9888,
  -37.0347,
  -37.0787,
  -37.1228,
  -37.1665,
  -37.2096,
  -37.2521,
  -37.2938,
  -37.3343,
  -37.373,
  -37.4094,
  -37.4429,
  -37.4733,
  -37.5005,
  -37.5251,
  -37.5475,
  -37.5682,
  -37.5874,
  -37.6057,
  -37.6237,
  -37.6418,
  -37.6607,
  -37.6808,
  -37.7022,
  -37.7247,
  -37.7479,
  -37.7713,
  -37.7942,
  -37.8162,
  -37.837,
  -37.8566,
  -37.875,
  -37.8925,
  -37.9092,
  -37.9239,
  -37.9385,
  -37.9515,
  -37.9627,
  -37.9722,
  -37.98,
  -37.9865,
  -37.9915,
  -37.9952,
  -37.9976,
  -37.9989,
  -37.9997,
  -38.0006,
  -38.002,
  -38.004,
  -38.0066,
  -38.0095,
  -38.0127,
  -38.0159,
  -38.019,
  -38.0218,
  -38.0241,
  -38.0256,
  -38.0264,
  -38.0263,
  -38.0255,
  -38.0241,
  -38.0222,
  -38.0195,
  -38.0155,
  -38.01,
  -38.0033,
  -37.9957,
  -37.9878,
  -37.9798,
  -37.9716,
  -37.9631,
  -37.9537,
  -37.9431,
  -37.9301,
  -37.9163,
  -37.9002,
  -37.8817,
  -37.8603,
  -37.8356,
  -37.8069,
  -37.7734,
  -37.7342,
  -37.6885,
  -37.6352,
  -37.5738,
  -37.5038,
  -37.4258,
  -37.3412,
  -37.2525,
  -37.1629,
  -37.0763,
  -36.9969,
  -36.929,
  -36.8767,
  -29.4042,
  -29.4499,
  -29.4955,
  -29.5411,
  -29.5871,
  -29.6337,
  -29.6813,
  -29.7299,
  -29.7794,
  -29.8297,
  -29.8806,
  -29.9307,
  -29.9816,
  -30.032,
  -30.0817,
  -30.1308,
  -30.1795,
  -30.2276,
  -30.2756,
  -30.3232,
  -30.37,
  -30.4159,
  -30.4605,
  -30.5036,
  -30.5455,
  -30.5863,
  -30.6259,
  -30.6668,
  -30.7088,
  -30.7527,
  -30.7991,
  -30.8483,
  -30.8999,
  -30.9528,
  -31.0058,
  -31.0575,
  -31.1066,
  -31.1535,
  -31.1981,
  -31.2412,
  -31.2835,
  -31.325,
  -31.3682,
  -31.4128,
  -31.4591,
  -31.507,
  -31.5559,
  -31.6053,
  -31.655,
  -31.7047,
  -31.7541,
  -31.803,
  -31.8513,
  -31.8991,
  -31.9469,
  -31.9948,
  -32.0432,
  -32.0907,
  -32.139,
  -32.1868,
  -32.2341,
  -32.2813,
  -32.3287,
  -32.3765,
  -32.4248,
  -32.4736,
  -32.5227,
  -32.5716,
  -32.6199,
  -32.6676,
  -32.7155,
  -32.7632,
  -32.8118,
  -32.8617,
  -32.9119,
  -32.9639,
  -33.0164,
  -33.0689,
  -33.1211,
  -33.1732,
  -33.2248,
  -33.2759,
  -33.3265,
  -33.3762,
  -33.4247,
  -33.472,
  -33.518,
  -33.5629,
  -33.607,
  -33.6505,
  -33.6936,
  -33.7358,
  -33.7794,
  -33.8233,
  -33.8673,
  -33.9109,
  -33.9536,
  -33.9953,
  -34.0358,
  -34.0753,
  -34.1135,
  -34.1505,
  -34.1859,
  -34.2197,
  -34.2519,
  -34.2828,
  -34.3128,
  -34.3423,
  -34.3715,
  -34.4003,
  -34.4274,
  -34.4546,
  -34.4807,
  -34.5056,
  -34.529,
  -34.5512,
  -34.5722,
  -34.5925,
  -34.6124,
  -34.6324,
  -34.6525,
  -34.6726,
  -34.6927,
  -34.7124,
  -34.7318,
  -34.7505,
  -34.7688,
  -34.7867,
  -34.8047,
  -34.8233,
  -34.8419,
  -34.8624,
  -34.8841,
  -34.9062,
  -34.9285,
  -34.9509,
  -34.9729,
  -34.9945,
  -35.0156,
  -35.036,
  -35.0554,
  -35.0738,
  -35.0914,
  -35.1082,
  -35.1248,
  -35.1419,
  -35.1602,
  -35.1802,
  -35.2017,
  -35.2247,
  -35.2488,
  -35.2729,
  -35.2989,
  -35.3255,
  -35.3522,
  -35.3781,
  -35.403,
  -35.4267,
  -35.4493,
  -35.4709,
  -35.4918,
  -35.5123,
  -35.5326,
  -35.5529,
  -35.5736,
  -35.5945,
  -35.6159,
  -35.6377,
  -35.6601,
  -35.683,
  -35.7059,
  -35.7287,
  -35.7512,
  -35.7732,
  -35.7937,
  -35.8145,
  -35.8346,
  -35.8547,
  -35.8754,
  -35.8971,
  -35.9196,
  -35.9421,
  -35.964,
  -35.9854,
  -36.0062,
  -36.0268,
  -36.0477,
  -36.069,
  -36.0913,
  -36.1149,
  -36.1407,
  -36.1693,
  -36.2018,
  -36.2384,
  -36.28,
  -36.3257,
  -36.3755,
  -36.4282,
  -36.483,
  -36.5388,
  -36.594,
  -36.6498,
  -36.7045,
  -36.7578,
  -36.8095,
  -36.8592,
  -36.9072,
  -36.954,
  -36.9998,
  -37.0446,
  -37.0886,
  -37.1321,
  -37.1749,
  -37.2172,
  -37.2588,
  -37.2993,
  -37.3383,
  -37.375,
  -37.4088,
  -37.4395,
  -37.467,
  -37.4918,
  -37.5143,
  -37.535,
  -37.5539,
  -37.5718,
  -37.5893,
  -37.607,
  -37.6253,
  -37.6451,
  -37.6653,
  -37.6875,
  -37.7102,
  -37.733,
  -37.7551,
  -37.7762,
  -37.7961,
  -37.8149,
  -37.8326,
  -37.8492,
  -37.8651,
  -37.88,
  -37.8937,
  -37.9062,
  -37.9172,
  -37.9266,
  -37.9345,
  -37.9408,
  -37.9455,
  -37.9489,
  -37.951,
  -37.9519,
  -37.9525,
  -37.953,
  -37.954,
  -37.9557,
  -37.9582,
  -37.9611,
  -37.9644,
  -37.9677,
  -37.971,
  -37.974,
  -37.9765,
  -37.9782,
  -37.979,
  -37.9788,
  -37.9768,
  -37.9754,
  -37.9737,
  -37.9717,
  -37.9687,
  -37.9645,
  -37.959,
  -37.9526,
  -37.9455,
  -37.938,
  -37.93,
  -37.9213,
  -37.9115,
  -37.9005,
  -37.888,
  -37.874,
  -37.8579,
  -37.8398,
  -37.8193,
  -37.7958,
  -37.7686,
  -37.7369,
  -37.6999,
  -37.657,
  -37.6074,
  -37.5503,
  -37.4858,
  -37.414,
  -37.3364,
  -37.2551,
  -37.1729,
  -37.0928,
  -37.0188,
  -36.9541,
  -36.9024,
  -29.3921,
  -29.4372,
  -29.4826,
  -29.5283,
  -29.5745,
  -29.6214,
  -29.669,
  -29.7165,
  -29.7657,
  -29.8154,
  -29.8657,
  -29.9163,
  -29.9668,
  -30.0169,
  -30.0664,
  -30.1153,
  -30.1637,
  -30.2117,
  -30.2592,
  -30.3062,
  -30.3521,
  -30.3958,
  -30.4391,
  -30.4812,
  -30.5223,
  -30.5628,
  -30.6033,
  -30.6444,
  -30.6868,
  -30.7311,
  -30.7778,
  -30.8272,
  -30.8788,
  -30.9317,
  -30.9846,
  -31.0361,
  -31.0843,
  -31.1309,
  -31.1753,
  -31.2182,
  -31.2606,
  -31.3031,
  -31.3463,
  -31.391,
  -31.4374,
  -31.4853,
  -31.5343,
  -31.5841,
  -31.634,
  -31.6839,
  -31.7333,
  -31.7819,
  -31.8286,
  -31.8755,
  -31.9223,
  -31.9694,
  -32.0169,
  -32.0649,
  -32.1131,
  -32.161,
  -32.2086,
  -32.2561,
  -32.3035,
  -32.351,
  -32.3988,
  -32.4472,
  -32.4959,
  -32.5446,
  -32.5921,
  -32.6402,
  -32.6882,
  -32.7361,
  -32.7845,
  -32.834,
  -32.8847,
  -32.9365,
  -32.9889,
  -33.0418,
  -33.0945,
  -33.1469,
  -33.199,
  -33.2505,
  -33.3013,
  -33.3512,
  -33.4,
  -33.4476,
  -33.4931,
  -33.5387,
  -33.5836,
  -33.6281,
  -33.6721,
  -33.716,
  -33.7599,
  -33.8038,
  -33.8476,
  -33.8907,
  -33.933,
  -33.9742,
  -34.0142,
  -34.0532,
  -34.0911,
  -34.1278,
  -34.1632,
  -34.1971,
  -34.2284,
  -34.2596,
  -34.2898,
  -34.3194,
  -34.3483,
  -34.3766,
  -34.4042,
  -34.4308,
  -34.4563,
  -34.4807,
  -34.5038,
  -34.5256,
  -34.5463,
  -34.5661,
  -34.5854,
  -34.6044,
  -34.6235,
  -34.6427,
  -34.6618,
  -34.6798,
  -34.6984,
  -34.7165,
  -34.734,
  -34.7512,
  -34.7685,
  -34.7862,
  -34.8046,
  -34.8238,
  -34.8438,
  -34.8643,
  -34.8851,
  -34.906,
  -34.927,
  -34.9476,
  -34.9681,
  -34.988,
  -35.0073,
  -35.0257,
  -35.0433,
  -35.0602,
  -35.0759,
  -35.0929,
  -35.111,
  -35.1303,
  -35.1509,
  -35.1727,
  -35.1957,
  -35.2198,
  -35.2451,
  -35.2712,
  -35.2975,
  -35.3233,
  -35.3484,
  -35.3722,
  -35.3952,
  -35.4173,
  -35.4387,
  -35.4597,
  -35.4804,
  -35.5011,
  -35.5218,
  -35.5429,
  -35.5644,
  -35.5855,
  -35.6083,
  -35.6317,
  -35.6552,
  -35.6785,
  -35.7016,
  -35.7241,
  -35.746,
  -35.7671,
  -35.7878,
  -35.8082,
  -35.8292,
  -35.8512,
  -35.8739,
  -35.8965,
  -35.9187,
  -35.9402,
  -35.9613,
  -35.9824,
  -36.0039,
  -36.0261,
  -36.0491,
  -36.0737,
  -36.1002,
  -36.1297,
  -36.1618,
  -36.1993,
  -36.2414,
  -36.2881,
  -36.3386,
  -36.3922,
  -36.4478,
  -36.5045,
  -36.5613,
  -36.6176,
  -36.6727,
  -36.7262,
  -36.7777,
  -36.8273,
  -36.8749,
  -36.921,
  -36.9663,
  -37.0107,
  -37.0544,
  -37.0974,
  -37.1399,
  -37.1819,
  -37.2231,
  -37.2636,
  -37.3026,
  -37.3395,
  -37.3738,
  -37.405,
  -37.4322,
  -37.4575,
  -37.4804,
  -37.5012,
  -37.5202,
  -37.538,
  -37.555,
  -37.5721,
  -37.5901,
  -37.6093,
  -37.63,
  -37.6518,
  -37.6741,
  -37.6962,
  -37.7176,
  -37.7379,
  -37.757,
  -37.7747,
  -37.7914,
  -37.8069,
  -37.8217,
  -37.8355,
  -37.8485,
  -37.8604,
  -37.8711,
  -37.8805,
  -37.8884,
  -37.8948,
  -37.8993,
  -37.9026,
  -37.9042,
  -37.905,
  -37.9051,
  -37.9055,
  -37.9052,
  -37.9067,
  -37.9089,
  -37.9119,
  -37.9153,
  -37.9189,
  -37.9224,
  -37.9258,
  -37.9284,
  -37.9302,
  -37.9308,
  -37.9303,
  -37.9292,
  -37.9278,
  -37.9263,
  -37.9248,
  -37.9229,
  -37.92,
  -37.9159,
  -37.9106,
  -37.9044,
  -37.8975,
  -37.8897,
  -37.8808,
  -37.8706,
  -37.8592,
  -37.8463,
  -37.8319,
  -37.816,
  -37.7984,
  -37.7788,
  -37.7565,
  -37.7308,
  -37.7008,
  -37.6661,
  -37.626,
  -37.5798,
  -37.5269,
  -37.4674,
  -37.4016,
  -37.3304,
  -37.2558,
  -37.1802,
  -37.1052,
  -37.0363,
  -36.9748,
  -36.9242,
  -29.3815,
  -29.4262,
  -29.4704,
  -29.5162,
  -29.5626,
  -29.6096,
  -29.6572,
  -29.7052,
  -29.7535,
  -29.8023,
  -29.8517,
  -29.9013,
  -29.951,
  -30.0006,
  -30.0498,
  -30.0986,
  -30.1469,
  -30.1935,
  -30.2406,
  -30.2868,
  -30.3319,
  -30.3757,
  -30.418,
  -30.4595,
  -30.5003,
  -30.541,
  -30.582,
  -30.6237,
  -30.6668,
  -30.7117,
  -30.7587,
  -30.8071,
  -30.8585,
  -30.911,
  -30.9633,
  -31.0145,
  -31.0635,
  -31.11,
  -31.1544,
  -31.1976,
  -31.24,
  -31.2826,
  -31.3261,
  -31.371,
  -31.4175,
  -31.4657,
  -31.515,
  -31.5639,
  -31.6142,
  -31.6641,
  -31.7134,
  -31.7617,
  -31.8087,
  -31.8547,
  -31.9004,
  -31.9463,
  -31.9928,
  -32.0402,
  -32.088,
  -32.136,
  -32.184,
  -32.2318,
  -32.2792,
  -32.3256,
  -32.3731,
  -32.4209,
  -32.4692,
  -32.5178,
  -32.5665,
  -32.615,
  -32.6633,
  -32.7116,
  -32.7599,
  -32.8091,
  -32.8592,
  -32.9106,
  -32.9632,
  -33.0161,
  -33.0691,
  -33.122,
  -33.1735,
  -33.2252,
  -33.2763,
  -33.3265,
  -33.3756,
  -33.4235,
  -33.4705,
  -33.5169,
  -33.5627,
  -33.6082,
  -33.6532,
  -33.6977,
  -33.742,
  -33.786,
  -33.8296,
  -33.8724,
  -33.9143,
  -33.9551,
  -33.9938,
  -34.0324,
  -34.07,
  -34.1065,
  -34.1418,
  -34.1757,
  -34.2082,
  -34.2395,
  -34.2699,
  -34.2994,
  -34.328,
  -34.3557,
  -34.3825,
  -34.4084,
  -34.4334,
  -34.4571,
  -34.4798,
  -34.5015,
  -34.5218,
  -34.5401,
  -34.559,
  -34.5771,
  -34.5949,
  -34.6127,
  -34.6307,
  -34.6486,
  -34.6664,
  -34.6838,
  -34.7006,
  -34.7173,
  -34.734,
  -34.7508,
  -34.7681,
  -34.7859,
  -34.8041,
  -34.8227,
  -34.8417,
  -34.8612,
  -34.8808,
  -34.8997,
  -34.9194,
  -34.9389,
  -34.9579,
  -34.9762,
  -34.9936,
  -35.0105,
  -35.0274,
  -35.0444,
  -35.0623,
  -35.0811,
  -35.101,
  -35.1219,
  -35.1438,
  -35.167,
  -35.1915,
  -35.2171,
  -35.243,
  -35.2687,
  -35.2936,
  -35.3178,
  -35.3411,
  -35.3626,
  -35.3847,
  -35.4061,
  -35.4271,
  -35.4479,
  -35.4687,
  -35.4899,
  -35.5115,
  -35.534,
  -35.5574,
  -35.5814,
  -35.6055,
  -35.6295,
  -35.6532,
  -35.6762,
  -35.6985,
  -35.72,
  -35.7409,
  -35.7617,
  -35.7828,
  -35.805,
  -35.8279,
  -35.8507,
  -35.8733,
  -35.8954,
  -35.916,
  -35.9378,
  -35.96,
  -35.983,
  -36.0072,
  -36.0326,
  -36.0601,
  -36.0904,
  -36.1243,
  -36.1626,
  -36.2055,
  -36.253,
  -36.3044,
  -36.3586,
  -36.4148,
  -36.472,
  -36.5293,
  -36.5861,
  -36.6417,
  -36.6953,
  -36.7467,
  -36.7959,
  -36.8429,
  -36.8884,
  -36.9329,
  -36.9767,
  -37.02,
  -37.0617,
  -37.1039,
  -37.1452,
  -37.186,
  -37.2262,
  -37.2651,
  -37.3023,
  -37.3369,
  -37.3687,
  -37.3978,
  -37.4241,
  -37.4476,
  -37.4689,
  -37.4882,
  -37.5059,
  -37.5227,
  -37.5393,
  -37.5566,
  -37.5752,
  -37.5952,
  -37.6163,
  -37.6381,
  -37.6598,
  -37.6805,
  -37.7001,
  -37.7182,
  -37.735,
  -37.7505,
  -37.7649,
  -37.7784,
  -37.7911,
  -37.8021,
  -37.8134,
  -37.8238,
  -37.8331,
  -37.841,
  -37.8473,
  -37.8518,
  -37.8548,
  -37.8563,
  -37.8567,
  -37.8568,
  -37.8569,
  -37.8577,
  -37.8592,
  -37.8615,
  -37.8646,
  -37.8682,
  -37.8721,
  -37.8759,
  -37.8794,
  -37.882,
  -37.8836,
  -37.8839,
  -37.8831,
  -37.8816,
  -37.8801,
  -37.8789,
  -37.8779,
  -37.877,
  -37.8752,
  -37.8723,
  -37.8684,
  -37.863,
  -37.8567,
  -37.8493,
  -37.8404,
  -37.83,
  -37.8181,
  -37.8049,
  -37.7903,
  -37.7735,
  -37.7565,
  -37.7377,
  -37.7167,
  -37.6923,
  -37.664,
  -37.6313,
  -37.5938,
  -37.5509,
  -37.5021,
  -37.4472,
  -37.3866,
  -37.321,
  -37.252,
  -37.1823,
  -37.1141,
  -37.0496,
  -36.9914,
  -36.9419,
  -29.3712,
  -29.4156,
  -29.4607,
  -29.5066,
  -29.5532,
  -29.6003,
  -29.6476,
  -29.6949,
  -29.7422,
  -29.7896,
  -29.8374,
  -29.8858,
  -29.9333,
  -29.9822,
  -30.0311,
  -30.0796,
  -30.1276,
  -30.1749,
  -30.2214,
  -30.2669,
  -30.3113,
  -30.3544,
  -30.3963,
  -30.4376,
  -30.4786,
  -30.52,
  -30.562,
  -30.6038,
  -30.6478,
  -30.6935,
  -30.7411,
  -30.7904,
  -30.8414,
  -30.8933,
  -30.9452,
  -30.9957,
  -31.0444,
  -31.0907,
  -31.135,
  -31.1781,
  -31.2207,
  -31.2637,
  -31.3065,
  -31.3516,
  -31.3984,
  -31.4468,
  -31.4963,
  -31.5467,
  -31.5971,
  -31.6472,
  -31.6964,
  -31.7441,
  -31.7904,
  -31.8354,
  -31.8799,
  -31.9244,
  -31.9698,
  -32.0163,
  -32.0627,
  -32.1107,
  -32.159,
  -32.2072,
  -32.2549,
  -32.3023,
  -32.3495,
  -32.3969,
  -32.4446,
  -32.493,
  -32.5419,
  -32.5907,
  -32.6395,
  -32.688,
  -32.7367,
  -32.7857,
  -32.8356,
  -32.8857,
  -32.9378,
  -32.9908,
  -33.0441,
  -33.0973,
  -33.1501,
  -33.2023,
  -33.2538,
  -33.3041,
  -33.3537,
  -33.4021,
  -33.4498,
  -33.4968,
  -33.5435,
  -33.5898,
  -33.6356,
  -33.6808,
  -33.7244,
  -33.7685,
  -33.8117,
  -33.8544,
  -33.8962,
  -33.9368,
  -33.9763,
  -34.0148,
  -34.0522,
  -34.0886,
  -34.1238,
  -34.1577,
  -34.1904,
  -34.2218,
  -34.2522,
  -34.2816,
  -34.3095,
  -34.3364,
  -34.3623,
  -34.3864,
  -34.4106,
  -34.4339,
  -34.4561,
  -34.4773,
  -34.4976,
  -34.5167,
  -34.5345,
  -34.5515,
  -34.5682,
  -34.5846,
  -34.6011,
  -34.6177,
  -34.6343,
  -34.6509,
  -34.6672,
  -34.6835,
  -34.6997,
  -34.716,
  -34.7322,
  -34.7475,
  -34.7639,
  -34.7805,
  -34.7975,
  -34.8152,
  -34.8334,
  -34.8523,
  -34.8714,
  -34.8902,
  -34.9088,
  -34.9267,
  -34.944,
  -34.961,
  -34.9779,
  -34.9951,
  -35.0129,
  -35.0311,
  -35.0503,
  -35.0704,
  -35.0917,
  -35.1141,
  -35.137,
  -35.1619,
  -35.1874,
  -35.2128,
  -35.2377,
  -35.2619,
  -35.2857,
  -35.3087,
  -35.3311,
  -35.3529,
  -35.3741,
  -35.395,
  -35.4159,
  -35.4372,
  -35.4592,
  -35.4821,
  -35.5061,
  -35.5306,
  -35.5554,
  -35.5801,
  -35.6043,
  -35.6279,
  -35.6506,
  -35.6722,
  -35.6924,
  -35.7133,
  -35.7348,
  -35.7571,
  -35.7802,
  -35.8036,
  -35.8268,
  -35.8497,
  -35.8723,
  -35.895,
  -35.9182,
  -35.9422,
  -35.9672,
  -35.9937,
  -36.0222,
  -36.0534,
  -36.0883,
  -36.1273,
  -36.1711,
  -36.2193,
  -36.2713,
  -36.3261,
  -36.3827,
  -36.4402,
  -36.4979,
  -36.555,
  -36.6099,
  -36.6637,
  -36.7149,
  -36.7634,
  -36.8096,
  -36.8541,
  -36.8978,
  -36.941,
  -36.9839,
  -37.0262,
  -37.0678,
  -37.1088,
  -37.1493,
  -37.1893,
  -37.2281,
  -37.2653,
  -37.3002,
  -37.3328,
  -37.3626,
  -37.3901,
  -37.4147,
  -37.4369,
  -37.4566,
  -37.4744,
  -37.4908,
  -37.5071,
  -37.5237,
  -37.5413,
  -37.5605,
  -37.5809,
  -37.601,
  -37.622,
  -37.6423,
  -37.6611,
  -37.6784,
  -37.6942,
  -37.7086,
  -37.7218,
  -37.734,
  -37.7456,
  -37.7565,
  -37.7672,
  -37.7772,
  -37.7864,
  -37.7943,
  -37.8006,
  -37.8051,
  -37.8079,
  -37.8092,
  -37.8095,
  -37.8094,
  -37.8098,
  -37.8107,
  -37.8126,
  -37.8153,
  -37.8186,
  -37.8225,
  -37.8267,
  -37.8306,
  -37.8341,
  -37.8364,
  -37.8374,
  -37.837,
  -37.8356,
  -37.8337,
  -37.8321,
  -37.83,
  -37.8296,
  -37.8293,
  -37.8287,
  -37.8271,
  -37.8241,
  -37.8197,
  -37.8142,
  -37.8073,
  -37.7987,
  -37.7884,
  -37.7763,
  -37.7629,
  -37.7483,
  -37.7327,
  -37.7161,
  -37.6981,
  -37.6779,
  -37.6549,
  -37.6281,
  -37.5973,
  -37.5623,
  -37.5225,
  -37.4775,
  -37.4269,
  -37.3709,
  -37.3103,
  -37.2465,
  -37.1816,
  -37.1178,
  -37.0574,
  -37.0021,
  -36.9541,
  -29.363,
  -29.4072,
  -29.4522,
  -29.4981,
  -29.5449,
  -29.5921,
  -29.6392,
  -29.6858,
  -29.7307,
  -29.7765,
  -29.8225,
  -29.8691,
  -29.9163,
  -29.9642,
  -30.0124,
  -30.0605,
  -30.1082,
  -30.1551,
  -30.2011,
  -30.2459,
  -30.2897,
  -30.3324,
  -30.3734,
  -30.4149,
  -30.4566,
  -30.499,
  -30.5421,
  -30.5863,
  -30.6318,
  -30.6786,
  -30.7267,
  -30.7762,
  -30.8267,
  -30.8779,
  -30.9289,
  -30.9788,
  -31.0268,
  -31.0717,
  -31.1159,
  -31.1589,
  -31.2018,
  -31.245,
  -31.2892,
  -31.3347,
  -31.3817,
  -31.4302,
  -31.48,
  -31.5305,
  -31.5812,
  -31.6313,
  -31.6803,
  -31.7276,
  -31.7731,
  -31.8162,
  -31.8594,
  -31.9027,
  -31.9469,
  -31.9924,
  -32.0393,
  -32.0873,
  -32.1358,
  -32.1843,
  -32.2324,
  -32.28,
  -32.3271,
  -32.3742,
  -32.4216,
  -32.4698,
  -32.5183,
  -32.5664,
  -32.6154,
  -32.6643,
  -32.7132,
  -32.7624,
  -32.8124,
  -32.8632,
  -32.9152,
  -32.9679,
  -33.0212,
  -33.0746,
  -33.1278,
  -33.1804,
  -33.2323,
  -33.2832,
  -33.3333,
  -33.3825,
  -33.4307,
  -33.4775,
  -33.5248,
  -33.5717,
  -33.6182,
  -33.6639,
  -33.7087,
  -33.7527,
  -33.796,
  -33.8385,
  -33.8803,
  -33.9211,
  -33.9608,
  -33.9993,
  -34.0366,
  -34.0729,
  -34.1082,
  -34.1422,
  -34.1751,
  -34.2057,
  -34.2361,
  -34.2649,
  -34.2921,
  -34.318,
  -34.3426,
  -34.3666,
  -34.39,
  -34.4126,
  -34.4345,
  -34.4552,
  -34.475,
  -34.4937,
  -34.5107,
  -34.5268,
  -34.5422,
  -34.5572,
  -34.572,
  -34.5869,
  -34.6011,
  -34.6166,
  -34.6324,
  -34.6485,
  -34.6644,
  -34.68,
  -34.6953,
  -34.7101,
  -34.7246,
  -34.7392,
  -34.7541,
  -34.7698,
  -34.7865,
  -34.804,
  -34.8223,
  -34.8406,
  -34.8588,
  -34.8764,
  -34.8936,
  -34.9106,
  -34.9275,
  -34.9437,
  -34.9612,
  -34.9791,
  -34.9974,
  -35.0168,
  -35.0375,
  -35.0595,
  -35.0828,
  -35.1073,
  -35.1324,
  -35.1575,
  -35.1823,
  -35.2067,
  -35.2307,
  -35.2541,
  -35.2768,
  -35.2988,
  -35.3201,
  -35.3411,
  -35.3621,
  -35.3835,
  -35.406,
  -35.4294,
  -35.4529,
  -35.4781,
  -35.5036,
  -35.5289,
  -35.5536,
  -35.5775,
  -35.6004,
  -35.6223,
  -35.6436,
  -35.6649,
  -35.6867,
  -35.7095,
  -35.7331,
  -35.7572,
  -35.7814,
  -35.8053,
  -35.8291,
  -35.8529,
  -35.877,
  -35.9019,
  -35.928,
  -35.9555,
  -35.9851,
  -36.0174,
  -36.0533,
  -36.0923,
  -36.137,
  -36.1858,
  -36.2384,
  -36.2934,
  -36.3502,
  -36.4078,
  -36.4658,
  -36.5233,
  -36.5791,
  -36.6328,
  -36.6837,
  -36.7315,
  -36.7767,
  -36.8202,
  -36.8629,
  -36.9054,
  -36.9478,
  -36.9898,
  -37.0312,
  -37.072,
  -37.1122,
  -37.1519,
  -37.1906,
  -37.2275,
  -37.2629,
  -37.2959,
  -37.3269,
  -37.3554,
  -37.3801,
  -37.4031,
  -37.4234,
  -37.4415,
  -37.4579,
  -37.4737,
  -37.4897,
  -37.5064,
  -37.5246,
  -37.5441,
  -37.5644,
  -37.5848,
  -37.6043,
  -37.6225,
  -37.639,
  -37.6538,
  -37.6671,
  -37.6792,
  -37.6903,
  -37.7008,
  -37.7109,
  -37.7208,
  -37.7305,
  -37.7395,
  -37.7473,
  -37.7535,
  -37.7579,
  -37.7605,
  -37.7617,
  -37.7621,
  -37.7623,
  -37.763,
  -37.7646,
  -37.7671,
  -37.7694,
  -37.7732,
  -37.7774,
  -37.7817,
  -37.7852,
  -37.7884,
  -37.7901,
  -37.7902,
  -37.7887,
  -37.7865,
  -37.7843,
  -37.7825,
  -37.7814,
  -37.7813,
  -37.7814,
  -37.7816,
  -37.7809,
  -37.7792,
  -37.7759,
  -37.7714,
  -37.7652,
  -37.7573,
  -37.7474,
  -37.7356,
  -37.7223,
  -37.7079,
  -37.6925,
  -37.6763,
  -37.6587,
  -37.6391,
  -37.6169,
  -37.5916,
  -37.5626,
  -37.5301,
  -37.4933,
  -37.4518,
  -37.4051,
  -37.3533,
  -37.297,
  -37.2377,
  -37.177,
  -37.1172,
  -37.0599,
  -37.007,
  -36.9591,
  -29.3552,
  -29.3992,
  -29.4441,
  -29.4891,
  -29.5359,
  -29.5831,
  -29.63,
  -29.6757,
  -29.7207,
  -29.7651,
  -29.8093,
  -29.8543,
  -29.9001,
  -29.9467,
  -29.9939,
  -30.0415,
  -30.0886,
  -30.1342,
  -30.1798,
  -30.2241,
  -30.2675,
  -30.3103,
  -30.3525,
  -30.3945,
  -30.437,
  -30.4803,
  -30.5248,
  -30.5705,
  -30.6174,
  -30.6654,
  -30.7141,
  -30.7638,
  -30.813,
  -30.8635,
  -30.9136,
  -30.9626,
  -31.0098,
  -31.0552,
  -31.0991,
  -31.1423,
  -31.1853,
  -31.2287,
  -31.2732,
  -31.319,
  -31.3662,
  -31.4148,
  -31.4647,
  -31.5153,
  -31.565,
  -31.6149,
  -31.6637,
  -31.7106,
  -31.7556,
  -31.7988,
  -31.8411,
  -31.8833,
  -31.9264,
  -31.9709,
  -32.0172,
  -32.0649,
  -32.1135,
  -32.1622,
  -32.2106,
  -32.2584,
  -32.3047,
  -32.3517,
  -32.3988,
  -32.4465,
  -32.495,
  -32.5444,
  -32.5935,
  -32.6426,
  -32.6918,
  -32.7414,
  -32.7916,
  -32.8423,
  -32.894,
  -32.9464,
  -32.9992,
  -33.0526,
  -33.1059,
  -33.158,
  -33.2105,
  -33.2622,
  -33.3131,
  -33.3631,
  -33.4122,
  -33.4605,
  -33.5084,
  -33.5558,
  -33.6025,
  -33.6486,
  -33.6936,
  -33.7378,
  -33.7809,
  -33.8235,
  -33.8654,
  -33.9065,
  -33.9464,
  -33.9841,
  -34.0217,
  -34.0582,
  -34.0936,
  -34.128,
  -34.1613,
  -34.1931,
  -34.2233,
  -34.2515,
  -34.2777,
  -34.3023,
  -34.3256,
  -34.3482,
  -34.3704,
  -34.3922,
  -34.4134,
  -34.4337,
  -34.4529,
  -34.4708,
  -34.4862,
  -34.5014,
  -34.5156,
  -34.5291,
  -34.5423,
  -34.5557,
  -34.5696,
  -34.5839,
  -34.5989,
  -34.6143,
  -34.6296,
  -34.6445,
  -34.6587,
  -34.672,
  -34.6847,
  -34.6973,
  -34.7102,
  -34.7239,
  -34.7389,
  -34.7549,
  -34.7723,
  -34.789,
  -34.8069,
  -34.8244,
  -34.8415,
  -34.8584,
  -34.8753,
  -34.8923,
  -34.9094,
  -34.9267,
  -34.9445,
  -34.9633,
  -34.983,
  -35.0047,
  -35.028,
  -35.0523,
  -35.0769,
  -35.1018,
  -35.1266,
  -35.1511,
  -35.1753,
  -35.1989,
  -35.2218,
  -35.2429,
  -35.2642,
  -35.2852,
  -35.3062,
  -35.3279,
  -35.3507,
  -35.3747,
  -35.3997,
  -35.4255,
  -35.4516,
  -35.4774,
  -35.5026,
  -35.5268,
  -35.5498,
  -35.5721,
  -35.5936,
  -35.6154,
  -35.638,
  -35.6615,
  -35.6858,
  -35.7108,
  -35.736,
  -35.7611,
  -35.7862,
  -35.81,
  -35.8352,
  -35.8611,
  -35.8882,
  -35.9169,
  -35.9476,
  -35.9811,
  -36.0181,
  -36.0591,
  -36.1046,
  -36.1542,
  -36.2071,
  -36.2626,
  -36.3197,
  -36.3776,
  -36.4354,
  -36.4928,
  -36.5484,
  -36.6017,
  -36.6521,
  -36.6992,
  -36.7434,
  -36.786,
  -36.8278,
  -36.8693,
  -36.9109,
  -36.9525,
  -36.9927,
  -37.0335,
  -37.0736,
  -37.113,
  -37.1514,
  -37.1882,
  -37.2234,
  -37.2571,
  -37.2888,
  -37.3182,
  -37.3451,
  -37.3689,
  -37.3899,
  -37.4085,
  -37.425,
  -37.4406,
  -37.456,
  -37.4721,
  -37.4893,
  -37.5078,
  -37.5271,
  -37.5466,
  -37.5654,
  -37.5828,
  -37.5985,
  -37.6125,
  -37.6249,
  -37.6361,
  -37.6463,
  -37.6559,
  -37.6651,
  -37.6744,
  -37.6825,
  -37.6911,
  -37.6986,
  -37.7047,
  -37.7089,
  -37.7114,
  -37.7127,
  -37.7133,
  -37.714,
  -37.7154,
  -37.7178,
  -37.7212,
  -37.7251,
  -37.7296,
  -37.7339,
  -37.7379,
  -37.7411,
  -37.7433,
  -37.7438,
  -37.7427,
  -37.7403,
  -37.7374,
  -37.7346,
  -37.7327,
  -37.7316,
  -37.7313,
  -37.7317,
  -37.7321,
  -37.7322,
  -37.7314,
  -37.7295,
  -37.7263,
  -37.7214,
  -37.7146,
  -37.7057,
  -37.6947,
  -37.682,
  -37.668,
  -37.6528,
  -37.6366,
  -37.6181,
  -37.5988,
  -37.5773,
  -37.5531,
  -37.526,
  -37.4958,
  -37.4618,
  -37.4236,
  -37.3805,
  -37.3325,
  -37.2802,
  -37.2249,
  -37.1681,
  -37.1115,
  -37.0569,
  -37.0058,
  -36.9595,
  -29.3467,
  -29.3903,
  -29.4351,
  -29.4809,
  -29.5276,
  -29.5746,
  -29.6211,
  -29.6665,
  -29.7107,
  -29.754,
  -29.7969,
  -29.8404,
  -29.8849,
  -29.9293,
  -29.9756,
  -30.0223,
  -30.0689,
  -30.115,
  -30.1602,
  -30.2044,
  -30.2478,
  -30.2906,
  -30.3332,
  -30.3759,
  -30.4193,
  -30.4636,
  -30.5093,
  -30.5562,
  -30.6034,
  -30.6524,
  -30.7017,
  -30.7514,
  -30.8013,
  -30.851,
  -30.9003,
  -30.9483,
  -30.9949,
  -31.0399,
  -31.0838,
  -31.1269,
  -31.17,
  -31.2137,
  -31.2584,
  -31.3033,
  -31.3506,
  -31.3993,
  -31.449,
  -31.4994,
  -31.5499,
  -31.5997,
  -31.6484,
  -31.695,
  -31.7396,
  -31.7824,
  -31.824,
  -31.8654,
  -31.9075,
  -31.9512,
  -31.9967,
  -32.0429,
  -32.0912,
  -32.1399,
  -32.1884,
  -32.2365,
  -32.2839,
  -32.3311,
  -32.3782,
  -32.426,
  -32.4743,
  -32.5232,
  -32.5726,
  -32.622,
  -32.6715,
  -32.7214,
  -32.7715,
  -32.8222,
  -32.8725,
  -32.9245,
  -32.9771,
  -33.0302,
  -33.0837,
  -33.1373,
  -33.1905,
  -33.2432,
  -33.295,
  -33.3458,
  -33.3956,
  -33.4446,
  -33.4929,
  -33.5407,
  -33.5878,
  -33.634,
  -33.6792,
  -33.7224,
  -33.7657,
  -33.8084,
  -33.8505,
  -33.8918,
  -33.932,
  -33.971,
  -34.0089,
  -34.0458,
  -34.0817,
  -34.1166,
  -34.1503,
  -34.1823,
  -34.2123,
  -34.2398,
  -34.265,
  -34.2882,
  -34.31,
  -34.3313,
  -34.3512,
  -34.3719,
  -34.3922,
  -34.4118,
  -34.4303,
  -34.4475,
  -34.4631,
  -34.4774,
  -34.4904,
  -34.5026,
  -34.5145,
  -34.5264,
  -34.5387,
  -34.5518,
  -34.5656,
  -34.58,
  -34.5943,
  -34.6081,
  -34.6209,
  -34.6328,
  -34.643,
  -34.6539,
  -34.665,
  -34.6769,
  -34.6901,
  -34.7047,
  -34.7212,
  -34.7384,
  -34.7558,
  -34.7732,
  -34.7901,
  -34.8067,
  -34.8233,
  -34.8399,
  -34.8565,
  -34.8733,
  -34.8904,
  -34.9087,
  -34.9285,
  -34.95,
  -34.9731,
  -34.9971,
  -35.0206,
  -35.0451,
  -35.0698,
  -35.0944,
  -35.1187,
  -35.1425,
  -35.1656,
  -35.1876,
  -35.209,
  -35.23,
  -35.2511,
  -35.2729,
  -35.2958,
  -35.3201,
  -35.3456,
  -35.3719,
  -35.3985,
  -35.4248,
  -35.4504,
  -35.4748,
  -35.4982,
  -35.5208,
  -35.5431,
  -35.5647,
  -35.5881,
  -35.6125,
  -35.6378,
  -35.6637,
  -35.6899,
  -35.7161,
  -35.7422,
  -35.7682,
  -35.7943,
  -35.8213,
  -35.8495,
  -35.8794,
  -35.9115,
  -35.9464,
  -35.9846,
  -36.0267,
  -36.0731,
  -36.1234,
  -36.177,
  -36.2327,
  -36.2899,
  -36.3478,
  -36.4056,
  -36.4626,
  -36.5179,
  -36.5696,
  -36.6191,
  -36.6655,
  -36.7091,
  -36.7507,
  -36.7915,
  -36.8321,
  -36.873,
  -36.914,
  -36.9548,
  -36.9953,
  -37.0353,
  -37.0744,
  -37.1124,
  -37.1491,
  -37.1843,
  -37.2181,
  -37.2503,
  -37.2806,
  -37.3083,
  -37.333,
  -37.3547,
  -37.3737,
  -37.3906,
  -37.4063,
  -37.4216,
  -37.4371,
  -37.4534,
  -37.4707,
  -37.489,
  -37.5075,
  -37.5244,
  -37.5411,
  -37.5561,
  -37.5693,
  -37.581,
  -37.5915,
  -37.6009,
  -37.6097,
  -37.6181,
  -37.6266,
  -37.635,
  -37.6431,
  -37.6501,
  -37.6557,
  -37.6598,
  -37.6625,
  -37.664,
  -37.6651,
  -37.6664,
  -37.6686,
  -37.6719,
  -37.6762,
  -37.681,
  -37.686,
  -37.6903,
  -37.6936,
  -37.696,
  -37.6968,
  -37.696,
  -37.6937,
  -37.6904,
  -37.6867,
  -37.6834,
  -37.6811,
  -37.6797,
  -37.6793,
  -37.6795,
  -37.6792,
  -37.6797,
  -37.6799,
  -37.6792,
  -37.6775,
  -37.6743,
  -37.6691,
  -37.6617,
  -37.6519,
  -37.6402,
  -37.6267,
  -37.6118,
  -37.5955,
  -37.5778,
  -37.5586,
  -37.5376,
  -37.5145,
  -37.4891,
  -37.4611,
  -37.4298,
  -37.3945,
  -37.3548,
  -37.3103,
  -37.2617,
  -37.2101,
  -37.1568,
  -37.1032,
  -37.0507,
  -37.0008,
  -36.9545,
  -29.3393,
  -29.3826,
  -29.4268,
  -29.4722,
  -29.5185,
  -29.565,
  -29.6113,
  -29.6563,
  -29.699,
  -29.7417,
  -29.784,
  -29.8266,
  -29.87,
  -29.9145,
  -29.9598,
  -30.0057,
  -30.0517,
  -30.0974,
  -30.1424,
  -30.1865,
  -30.2301,
  -30.2731,
  -30.3161,
  -30.3585,
  -30.4026,
  -30.4479,
  -30.4946,
  -30.5427,
  -30.5916,
  -30.6411,
  -30.6908,
  -30.7404,
  -30.7898,
  -30.8388,
  -30.8874,
  -30.9349,
  -30.9808,
  -31.0256,
  -31.0684,
  -31.1117,
  -31.1551,
  -31.199,
  -31.2439,
  -31.29,
  -31.3372,
  -31.3856,
  -31.435,
  -31.4849,
  -31.535,
  -31.5845,
  -31.6329,
  -31.6795,
  -31.724,
  -31.7667,
  -31.8071,
  -31.848,
  -31.8895,
  -31.9324,
  -31.9771,
  -32.0235,
  -32.0712,
  -32.1195,
  -32.1679,
  -32.216,
  -32.2635,
  -32.3109,
  -32.3584,
  -32.4061,
  -32.4545,
  -32.5034,
  -32.5517,
  -32.6012,
  -32.6509,
  -32.7011,
  -32.7513,
  -32.8019,
  -32.8529,
  -32.9046,
  -32.9568,
  -33.0094,
  -33.0631,
  -33.1172,
  -33.1713,
  -33.2249,
  -33.2776,
  -33.3292,
  -33.3797,
  -33.4292,
  -33.4771,
  -33.5252,
  -33.5726,
  -33.6191,
  -33.6645,
  -33.7089,
  -33.7524,
  -33.7953,
  -33.8376,
  -33.8791,
  -33.9196,
  -33.9589,
  -33.9972,
  -34.0345,
  -34.071,
  -34.1065,
  -34.1406,
  -34.1728,
  -34.2016,
  -34.2285,
  -34.2527,
  -34.2747,
  -34.2952,
  -34.3152,
  -34.3348,
  -34.3542,
  -34.3734,
  -34.392,
  -34.4097,
  -34.426,
  -34.4407,
  -34.4541,
  -34.466,
  -34.477,
  -34.4875,
  -34.4979,
  -34.5088,
  -34.5204,
  -34.5318,
  -34.5448,
  -34.5577,
  -34.57,
  -34.5814,
  -34.5919,
  -34.6016,
  -34.611,
  -34.6206,
  -34.6309,
  -34.6425,
  -34.6561,
  -34.6717,
  -34.6883,
  -34.7054,
  -34.7223,
  -34.7388,
  -34.755,
  -34.771,
  -34.7869,
  -34.8029,
  -34.8181,
  -34.8349,
  -34.8531,
  -34.8728,
  -34.8944,
  -34.9174,
  -34.9413,
  -34.9654,
  -34.9897,
  -35.0143,
  -35.0389,
  -35.0633,
  -35.0873,
  -35.1103,
  -35.1324,
  -35.1537,
  -35.1745,
  -35.1956,
  -35.2174,
  -35.2406,
  -35.2652,
  -35.2911,
  -35.3178,
  -35.3438,
  -35.3705,
  -35.3963,
  -35.4211,
  -35.4448,
  -35.4679,
  -35.4909,
  -35.5147,
  -35.5393,
  -35.5648,
  -35.5911,
  -35.6179,
  -35.645,
  -35.6721,
  -35.699,
  -35.726,
  -35.7533,
  -35.7813,
  -35.8107,
  -35.8418,
  -35.8753,
  -35.9115,
  -35.9511,
  -35.9944,
  -36.0418,
  -36.0919,
  -36.146,
  -36.2021,
  -36.2595,
  -36.3174,
  -36.375,
  -36.4316,
  -36.4862,
  -36.5381,
  -36.587,
  -36.6328,
  -36.6757,
  -36.7167,
  -36.7565,
  -36.7961,
  -36.8361,
  -36.8763,
  -36.9166,
  -36.9569,
  -36.9967,
  -37.0355,
  -37.0731,
  -37.1095,
  -37.1446,
  -37.1785,
  -37.211,
  -37.2417,
  -37.27,
  -37.2952,
  -37.3166,
  -37.3362,
  -37.3537,
  -37.37,
  -37.3854,
  -37.4006,
  -37.4161,
  -37.4323,
  -37.4493,
  -37.4666,
  -37.4835,
  -37.4994,
  -37.5137,
  -37.5263,
  -37.5374,
  -37.5472,
  -37.556,
  -37.5641,
  -37.5718,
  -37.5795,
  -37.5871,
  -37.5945,
  -37.6008,
  -37.6062,
  -37.6102,
  -37.6129,
  -37.6147,
  -37.6163,
  -37.6183,
  -37.6213,
  -37.6255,
  -37.6307,
  -37.6363,
  -37.6415,
  -37.6446,
  -37.6473,
  -37.6484,
  -37.6477,
  -37.6455,
  -37.6419,
  -37.6375,
  -37.6332,
  -37.6295,
  -37.6266,
  -37.6248,
  -37.6239,
  -37.6239,
  -37.6245,
  -37.6255,
  -37.6265,
  -37.6272,
  -37.6271,
  -37.6257,
  -37.6225,
  -37.6169,
  -37.6088,
  -37.5983,
  -37.5856,
  -37.5709,
  -37.5546,
  -37.5367,
  -37.5175,
  -37.4969,
  -37.475,
  -37.4513,
  -37.4253,
  -37.3965,
  -37.3641,
  -37.3273,
  -37.2861,
  -37.2409,
  -37.1927,
  -37.1425,
  -37.0915,
  -37.041,
  -36.9918,
  -36.9451,
  -29.3323,
  -29.3749,
  -29.4183,
  -29.4629,
  -29.5074,
  -29.5534,
  -29.5991,
  -29.6439,
  -29.6875,
  -29.7301,
  -29.7722,
  -29.8146,
  -29.8577,
  -29.9013,
  -29.9459,
  -29.9911,
  -30.0366,
  -30.0818,
  -30.1257,
  -30.1698,
  -30.2136,
  -30.257,
  -30.3005,
  -30.3446,
  -30.3894,
  -30.4354,
  -30.4829,
  -30.5314,
  -30.5809,
  -30.6306,
  -30.6801,
  -30.7295,
  -30.7783,
  -30.8258,
  -30.8736,
  -30.9205,
  -30.9664,
  -31.0114,
  -31.0553,
  -31.0991,
  -31.1428,
  -31.187,
  -31.2322,
  -31.2783,
  -31.3254,
  -31.3734,
  -31.422,
  -31.4711,
  -31.5204,
  -31.5684,
  -31.6165,
  -31.6632,
  -31.708,
  -31.7509,
  -31.7925,
  -31.8333,
  -31.8744,
  -31.9165,
  -31.9602,
  -32.0056,
  -32.0525,
  -32.1001,
  -32.148,
  -32.196,
  -32.2436,
  -32.2903,
  -32.338,
  -32.3858,
  -32.4345,
  -32.4835,
  -32.5327,
  -32.5823,
  -32.6322,
  -32.6824,
  -32.7326,
  -32.7834,
  -32.8341,
  -32.8853,
  -32.937,
  -32.9899,
  -33.0436,
  -33.0982,
  -33.152,
  -33.2064,
  -33.2599,
  -33.3122,
  -33.363,
  -33.413,
  -33.4623,
  -33.511,
  -33.559,
  -33.6058,
  -33.6517,
  -33.6965,
  -33.7405,
  -33.7835,
  -33.8259,
  -33.8675,
  -33.9081,
  -33.9477,
  -33.9852,
  -34.0231,
  -34.06,
  -34.096,
  -34.1306,
  -34.163,
  -34.1924,
  -34.2187,
  -34.2423,
  -34.2635,
  -34.2832,
  -34.3021,
  -34.3204,
  -34.3386,
  -34.3566,
  -34.3741,
  -34.3906,
  -34.4057,
  -34.4195,
  -34.4307,
  -34.4416,
  -34.4513,
  -34.4605,
  -34.4695,
  -34.479,
  -34.4892,
  -34.4999,
  -34.5111,
  -34.5223,
  -34.5328,
  -34.5426,
  -34.5517,
  -34.5601,
  -34.5682,
  -34.5765,
  -34.5855,
  -34.5961,
  -34.6089,
  -34.6235,
  -34.6395,
  -34.655,
  -34.6713,
  -34.6871,
  -34.7024,
  -34.7175,
  -34.7326,
  -34.7479,
  -34.7637,
  -34.7806,
  -34.799,
  -34.819,
  -34.8408,
  -34.8637,
  -34.8873,
  -34.9111,
  -34.9352,
  -34.9593,
  -34.9838,
  -35.0082,
  -35.0322,
  -35.0552,
  -35.0771,
  -35.0972,
  -35.1179,
  -35.1389,
  -35.161,
  -35.1844,
  -35.2094,
  -35.2356,
  -35.2627,
  -35.2899,
  -35.317,
  -35.343,
  -35.3678,
  -35.3917,
  -35.4154,
  -35.4396,
  -35.4646,
  -35.4906,
  -35.5174,
  -35.5447,
  -35.5724,
  -35.6001,
  -35.6278,
  -35.6555,
  -35.6834,
  -35.7116,
  -35.7399,
  -35.7704,
  -35.803,
  -35.8379,
  -35.8755,
  -35.9165,
  -35.9612,
  -36.0096,
  -36.0614,
  -36.1161,
  -36.1727,
  -36.2302,
  -36.288,
  -36.3453,
  -36.4012,
  -36.4552,
  -36.5066,
  -36.5549,
  -36.6001,
  -36.6427,
  -36.6832,
  -36.7222,
  -36.7608,
  -36.7995,
  -36.839,
  -36.8788,
  -36.9184,
  -36.9569,
  -36.9954,
  -37.0327,
  -37.0687,
  -37.1036,
  -37.1374,
  -37.1698,
  -37.2005,
  -37.2289,
  -37.2546,
  -37.2775,
  -37.298,
  -37.3166,
  -37.3337,
  -37.3495,
  -37.3646,
  -37.3795,
  -37.3947,
  -37.4103,
  -37.4262,
  -37.442,
  -37.4569,
  -37.4704,
  -37.4825,
  -37.493,
  -37.5023,
  -37.5105,
  -37.518,
  -37.5252,
  -37.5322,
  -37.539,
  -37.5455,
  -37.5503,
  -37.5551,
  -37.559,
  -37.5617,
  -37.564,
  -37.5662,
  -37.5689,
  -37.5726,
  -37.5776,
  -37.5834,
  -37.5894,
  -37.5945,
  -37.5982,
  -37.5999,
  -37.5996,
  -37.5974,
  -37.5938,
  -37.589,
  -37.5839,
  -37.579,
  -37.5747,
  -37.5712,
  -37.5689,
  -37.5675,
  -37.5672,
  -37.5677,
  -37.569,
  -37.5709,
  -37.5728,
  -37.5744,
  -37.575,
  -37.5738,
  -37.5702,
  -37.564,
  -37.5548,
  -37.543,
  -37.5288,
  -37.5125,
  -37.4947,
  -37.4755,
  -37.4555,
  -37.4338,
  -37.4119,
  -37.3882,
  -37.3618,
  -37.332,
  -37.2979,
  -37.2595,
  -37.2174,
  -37.1723,
  -37.125,
  -37.0763,
  -37.0272,
  -36.9786,
  -36.9315,
  -29.3244,
  -29.366,
  -29.4087,
  -29.4523,
  -29.4969,
  -29.5422,
  -29.5874,
  -29.6319,
  -29.6755,
  -29.7182,
  -29.7605,
  -29.8028,
  -29.8456,
  -29.8892,
  -29.9322,
  -29.977,
  -30.0223,
  -30.0674,
  -30.1122,
  -30.1566,
  -30.2005,
  -30.2441,
  -30.2881,
  -30.3326,
  -30.3782,
  -30.4249,
  -30.473,
  -30.5221,
  -30.5716,
  -30.6204,
  -30.6696,
  -30.7184,
  -30.7666,
  -30.8142,
  -30.8613,
  -30.9076,
  -30.9534,
  -30.9987,
  -31.0435,
  -31.088,
  -31.1325,
  -31.1774,
  -31.2228,
  -31.2688,
  -31.3143,
  -31.3614,
  -31.4091,
  -31.4571,
  -31.5056,
  -31.5541,
  -31.6021,
  -31.649,
  -31.6941,
  -31.7376,
  -31.7795,
  -31.8204,
  -31.8612,
  -31.9027,
  -31.9455,
  -31.9897,
  -32.0345,
  -32.0812,
  -32.1286,
  -32.1763,
  -32.2241,
  -32.2719,
  -32.3199,
  -32.368,
  -32.4166,
  -32.4656,
  -32.5147,
  -32.564,
  -32.6136,
  -32.6635,
  -32.7137,
  -32.7645,
  -32.8153,
  -32.866,
  -32.9176,
  -32.9705,
  -33.0246,
  -33.0795,
  -33.1349,
  -33.1899,
  -33.2439,
  -33.2965,
  -33.3477,
  -33.3983,
  -33.4481,
  -33.4975,
  -33.546,
  -33.5935,
  -33.6399,
  -33.6853,
  -33.7287,
  -33.7721,
  -33.8146,
  -33.8561,
  -33.8967,
  -33.9363,
  -33.9751,
  -34.0132,
  -34.0506,
  -34.087,
  -34.1219,
  -34.1542,
  -34.1835,
  -34.2097,
  -34.2327,
  -34.2534,
  -34.2726,
  -34.2906,
  -34.3081,
  -34.3242,
  -34.341,
  -34.3572,
  -34.3724,
  -34.3863,
  -34.3987,
  -34.4097,
  -34.4192,
  -34.4276,
  -34.4355,
  -34.4432,
  -34.4513,
  -34.4598,
  -34.4688,
  -34.4781,
  -34.4872,
  -34.496,
  -34.5041,
  -34.5117,
  -34.5188,
  -34.5248,
  -34.5321,
  -34.5404,
  -34.5504,
  -34.5625,
  -34.5764,
  -34.5914,
  -34.607,
  -34.6222,
  -34.6369,
  -34.6511,
  -34.6652,
  -34.6794,
  -34.6941,
  -34.7099,
  -34.727,
  -34.7459,
  -34.7663,
  -34.7883,
  -34.8111,
  -34.8344,
  -34.8579,
  -34.8805,
  -34.9045,
  -34.9288,
  -34.953,
  -34.9767,
  -34.9995,
  -35.0211,
  -35.0418,
  -35.0624,
  -35.0835,
  -35.1057,
  -35.1294,
  -35.1547,
  -35.1813,
  -35.2087,
  -35.2362,
  -35.2634,
  -35.2896,
  -35.3145,
  -35.3387,
  -35.3629,
  -35.3881,
  -35.4143,
  -35.4417,
  -35.4688,
  -35.4973,
  -35.5258,
  -35.5542,
  -35.5825,
  -35.6107,
  -35.6393,
  -35.6685,
  -35.6988,
  -35.7307,
  -35.7647,
  -35.801,
  -35.8403,
  -35.8829,
  -35.9289,
  -35.9783,
  -36.0309,
  -36.086,
  -36.1427,
  -36.2002,
  -36.2578,
  -36.3147,
  -36.3702,
  -36.4235,
  -36.4743,
  -36.5223,
  -36.5663,
  -36.6087,
  -36.6487,
  -36.6872,
  -36.7251,
  -36.7631,
  -36.8018,
  -36.8409,
  -36.8802,
  -36.9189,
  -36.9569,
  -36.9937,
  -37.0293,
  -37.0636,
  -37.097,
  -37.1291,
  -37.1595,
  -37.1878,
  -37.2137,
  -37.2374,
  -37.2588,
  -37.2786,
  -37.2966,
  -37.3131,
  -37.3283,
  -37.3427,
  -37.3569,
  -37.3712,
  -37.3856,
  -37.3999,
  -37.4136,
  -37.4253,
  -37.4367,
  -37.4467,
  -37.4556,
  -37.4634,
  -37.4705,
  -37.4771,
  -37.4834,
  -37.4896,
  -37.4953,
  -37.5005,
  -37.505,
  -37.5086,
  -37.5116,
  -37.5142,
  -37.5171,
  -37.5204,
  -37.5248,
  -37.5303,
  -37.5363,
  -37.5422,
  -37.5469,
  -37.5498,
  -37.5505,
  -37.5488,
  -37.5451,
  -37.5403,
  -37.5347,
  -37.5289,
  -37.5233,
  -37.5184,
  -37.5145,
  -37.5117,
  -37.5099,
  -37.5094,
  -37.5101,
  -37.5118,
  -37.5133,
  -37.5163,
  -37.5193,
  -37.5216,
  -37.5223,
  -37.5205,
  -37.5159,
  -37.5081,
  -37.4974,
  -37.484,
  -37.4683,
  -37.4509,
  -37.4325,
  -37.4134,
  -37.3941,
  -37.3739,
  -37.3523,
  -37.3282,
  -37.3006,
  -37.269,
  -37.2332,
  -37.1938,
  -37.1514,
  -37.1065,
  -37.0599,
  -37.0119,
  -36.9639,
  -36.9165,
  -29.3176,
  -29.3583,
  -29.4,
  -29.4426,
  -29.4863,
  -29.5307,
  -29.5754,
  -29.6198,
  -29.6634,
  -29.7055,
  -29.7481,
  -29.7907,
  -29.8335,
  -29.8768,
  -29.9207,
  -29.9654,
  -30.0105,
  -30.0557,
  -30.1007,
  -30.1451,
  -30.1893,
  -30.2334,
  -30.2779,
  -30.3229,
  -30.3681,
  -30.4154,
  -30.4638,
  -30.5132,
  -30.5627,
  -30.6122,
  -30.6612,
  -30.7094,
  -30.7569,
  -30.8038,
  -30.85,
  -30.8959,
  -30.9416,
  -30.9874,
  -31.0332,
  -31.0779,
  -31.1235,
  -31.1692,
  -31.2148,
  -31.2605,
  -31.3063,
  -31.3522,
  -31.3985,
  -31.4453,
  -31.4928,
  -31.5408,
  -31.5887,
  -31.6359,
  -31.6817,
  -31.7257,
  -31.7681,
  -31.8083,
  -31.8491,
  -31.8901,
  -31.932,
  -31.9751,
  -32.0196,
  -32.0654,
  -32.112,
  -32.1595,
  -32.2072,
  -32.2552,
  -32.3034,
  -32.3516,
  -32.4001,
  -32.4488,
  -32.4976,
  -32.5455,
  -32.5947,
  -32.6443,
  -32.6945,
  -32.7453,
  -32.7967,
  -32.8485,
  -32.9012,
  -32.9545,
  -33.0086,
  -33.0637,
  -33.1192,
  -33.1746,
  -33.2287,
  -33.2815,
  -33.3332,
  -33.384,
  -33.4346,
  -33.4836,
  -33.5329,
  -33.5812,
  -33.6283,
  -33.6744,
  -33.7193,
  -33.7629,
  -33.8054,
  -33.8468,
  -33.8872,
  -33.9267,
  -33.9656,
  -34.0038,
  -34.0415,
  -34.0782,
  -34.113,
  -34.1454,
  -34.1747,
  -34.1996,
  -34.2224,
  -34.243,
  -34.2619,
  -34.2796,
  -34.2963,
  -34.3125,
  -34.3282,
  -34.3432,
  -34.3571,
  -34.3696,
  -34.3806,
  -34.3899,
  -34.398,
  -34.4049,
  -34.4114,
  -34.4179,
  -34.4246,
  -34.4316,
  -34.4388,
  -34.4451,
  -34.4522,
  -34.459,
  -34.4654,
  -34.4715,
  -34.4773,
  -34.4832,
  -34.4897,
  -34.4974,
  -34.507,
  -34.5186,
  -34.5317,
  -34.5457,
  -34.5599,
  -34.5738,
  -34.5873,
  -34.6003,
  -34.6133,
  -34.6267,
  -34.6411,
  -34.657,
  -34.6736,
  -34.6929,
  -34.714,
  -34.7359,
  -34.7585,
  -34.7814,
  -34.8045,
  -34.8279,
  -34.8517,
  -34.8757,
  -34.8997,
  -34.923,
  -34.9452,
  -34.9663,
  -34.9867,
  -35.0071,
  -35.0282,
  -35.0506,
  -35.0746,
  -35.1003,
  -35.1271,
  -35.1548,
  -35.1827,
  -35.209,
  -35.2353,
  -35.2603,
  -35.2847,
  -35.3095,
  -35.3353,
  -35.3627,
  -35.3915,
  -35.4209,
  -35.4506,
  -35.48,
  -35.5091,
  -35.5379,
  -35.5668,
  -35.5961,
  -35.6263,
  -35.6578,
  -35.691,
  -35.7264,
  -35.7644,
  -35.8053,
  -35.8495,
  -35.8968,
  -35.9472,
  -36.0004,
  -36.0545,
  -36.111,
  -36.1683,
  -36.2255,
  -36.282,
  -36.337,
  -36.39,
  -36.4405,
  -36.4883,
  -36.5333,
  -36.5756,
  -36.6154,
  -36.6536,
  -36.6909,
  -36.7285,
  -36.7666,
  -36.8053,
  -36.8438,
  -36.8818,
  -36.9188,
  -36.955,
  -36.9898,
  -37.0236,
  -37.0564,
  -37.0879,
  -37.1178,
  -37.1458,
  -37.1719,
  -37.1962,
  -37.2177,
  -37.2386,
  -37.2577,
  -37.2748,
  -37.2903,
  -37.3044,
  -37.3178,
  -37.3307,
  -37.3436,
  -37.3563,
  -37.3686,
  -37.3802,
  -37.3909,
  -37.4005,
  -37.4091,
  -37.4167,
  -37.4235,
  -37.4297,
  -37.4356,
  -37.4412,
  -37.4464,
  -37.4512,
  -37.4552,
  -37.4587,
  -37.4618,
  -37.4647,
  -37.4682,
  -37.4724,
  -37.4775,
  -37.4829,
  -37.4887,
  -37.4938,
  -37.4977,
  -37.4995,
  -37.4989,
  -37.4952,
  -37.4904,
  -37.4847,
  -37.4783,
  -37.4719,
  -37.4658,
  -37.4603,
  -37.4558,
  -37.4527,
  -37.4508,
  -37.4505,
  -37.4512,
  -37.4532,
  -37.4563,
  -37.4601,
  -37.4642,
  -37.4677,
  -37.4699,
  -37.4697,
  -37.4665,
  -37.4601,
  -37.4505,
  -37.4383,
  -37.4239,
  -37.4078,
  -37.3906,
  -37.3728,
  -37.3549,
  -37.3365,
  -37.3168,
  -37.2947,
  -37.2692,
  -37.2398,
  -37.2064,
  -37.1695,
  -37.1295,
  -37.0867,
  -37.0416,
  -36.9949,
  -36.9474,
  -36.8998,
  -29.3109,
  -29.3506,
  -29.3913,
  -29.4331,
  -29.4761,
  -29.5188,
  -29.563,
  -29.6071,
  -29.6508,
  -29.694,
  -29.7369,
  -29.7797,
  -29.8227,
  -29.8661,
  -29.9101,
  -29.9548,
  -30,
  -30.0453,
  -30.0903,
  -30.134,
  -30.1784,
  -30.223,
  -30.268,
  -30.3139,
  -30.3608,
  -30.4088,
  -30.4577,
  -30.5071,
  -30.5568,
  -30.606,
  -30.6544,
  -30.7019,
  -30.7485,
  -30.7945,
  -30.839,
  -30.8846,
  -30.9305,
  -30.9769,
  -31.0238,
  -31.0709,
  -31.1178,
  -31.1642,
  -31.2101,
  -31.2553,
  -31.3001,
  -31.3446,
  -31.3894,
  -31.4349,
  -31.4814,
  -31.529,
  -31.5759,
  -31.6235,
  -31.6699,
  -31.7146,
  -31.7576,
  -31.7992,
  -31.84,
  -31.8807,
  -31.9217,
  -31.9638,
  -32.0072,
  -32.052,
  -32.098,
  -32.145,
  -32.1926,
  -32.2405,
  -32.2878,
  -32.336,
  -32.3842,
  -32.4324,
  -32.4806,
  -32.529,
  -32.5777,
  -32.627,
  -32.6772,
  -32.7284,
  -32.7804,
  -32.833,
  -32.8865,
  -32.9405,
  -32.9951,
  -33.0503,
  -33.106,
  -33.1605,
  -33.2148,
  -33.2679,
  -33.3197,
  -33.3708,
  -33.4215,
  -33.4719,
  -33.5219,
  -33.5709,
  -33.6187,
  -33.6653,
  -33.7104,
  -33.7542,
  -33.7966,
  -33.8378,
  -33.8781,
  -33.9176,
  -33.9564,
  -33.9937,
  -34.0316,
  -34.0683,
  -34.1032,
  -34.1357,
  -34.1648,
  -34.1906,
  -34.2134,
  -34.234,
  -34.2527,
  -34.27,
  -34.2863,
  -34.3017,
  -34.3164,
  -34.3303,
  -34.343,
  -34.3542,
  -34.3637,
  -34.3715,
  -34.378,
  -34.3825,
  -34.3876,
  -34.3927,
  -34.3981,
  -34.4036,
  -34.4092,
  -34.4146,
  -34.4197,
  -34.4246,
  -34.4291,
  -34.4334,
  -34.4378,
  -34.4426,
  -34.4482,
  -34.4554,
  -34.4646,
  -34.4756,
  -34.4879,
  -34.5008,
  -34.5137,
  -34.5252,
  -34.5373,
  -34.5493,
  -34.5614,
  -34.5742,
  -34.5883,
  -34.6043,
  -34.6222,
  -34.642,
  -34.6633,
  -34.6852,
  -34.7076,
  -34.7301,
  -34.7529,
  -34.7761,
  -34.7997,
  -34.8235,
  -34.8471,
  -34.8699,
  -34.8915,
  -34.9122,
  -34.9322,
  -34.9515,
  -34.9726,
  -34.995,
  -35.0192,
  -35.045,
  -35.0721,
  -35.1,
  -35.1281,
  -35.1558,
  -35.1822,
  -35.2075,
  -35.2321,
  -35.2572,
  -35.2837,
  -35.312,
  -35.3417,
  -35.3724,
  -35.4032,
  -35.4336,
  -35.4635,
  -35.4932,
  -35.5229,
  -35.5531,
  -35.5844,
  -35.6172,
  -35.6508,
  -35.6877,
  -35.7273,
  -35.7698,
  -35.8154,
  -35.864,
  -35.9153,
  -35.9687,
  -36.0238,
  -36.0799,
  -36.1366,
  -36.1933,
  -36.2493,
  -36.304,
  -36.3567,
  -36.407,
  -36.4548,
  -36.4998,
  -36.542,
  -36.5817,
  -36.6197,
  -36.657,
  -36.6944,
  -36.7324,
  -36.7706,
  -36.8086,
  -36.8459,
  -36.882,
  -36.916,
  -36.9498,
  -36.9827,
  -37.0147,
  -37.0455,
  -37.075,
  -37.1028,
  -37.1291,
  -37.1538,
  -37.1772,
  -37.1989,
  -37.2188,
  -37.2367,
  -37.2524,
  -37.2665,
  -37.2792,
  -37.291,
  -37.3024,
  -37.3135,
  -37.3242,
  -37.3344,
  -37.3442,
  -37.3532,
  -37.3615,
  -37.3691,
  -37.3758,
  -37.382,
  -37.3877,
  -37.393,
  -37.3978,
  -37.402,
  -37.4057,
  -37.4079,
  -37.411,
  -37.4145,
  -37.4186,
  -37.4233,
  -37.4287,
  -37.4343,
  -37.4397,
  -37.4442,
  -37.4469,
  -37.4476,
  -37.4461,
  -37.4421,
  -37.4364,
  -37.4297,
  -37.4227,
  -37.4158,
  -37.4093,
  -37.4034,
  -37.3987,
  -37.3952,
  -37.3934,
  -37.3931,
  -37.394,
  -37.3963,
  -37.3998,
  -37.404,
  -37.4087,
  -37.413,
  -37.4161,
  -37.4171,
  -37.4152,
  -37.4101,
  -37.4021,
  -37.3915,
  -37.3789,
  -37.3646,
  -37.3491,
  -37.3331,
  -37.3167,
  -37.2998,
  -37.2817,
  -37.2603,
  -37.2366,
  -37.2092,
  -37.178,
  -37.1433,
  -37.1053,
  -37.0644,
  -37.0208,
  -36.9752,
  -36.9282,
  -36.8807,
  -29.3035,
  -29.3423,
  -29.3824,
  -29.4235,
  -29.4659,
  -29.5091,
  -29.5527,
  -29.5964,
  -29.64,
  -29.6833,
  -29.7263,
  -29.7693,
  -29.8125,
  -29.8561,
  -29.9004,
  -29.9444,
  -29.9898,
  -30.0352,
  -30.0804,
  -30.1252,
  -30.17,
  -30.2151,
  -30.2609,
  -30.3075,
  -30.3552,
  -30.4037,
  -30.4531,
  -30.5028,
  -30.5524,
  -30.6003,
  -30.6483,
  -30.6951,
  -30.741,
  -30.7863,
  -30.8313,
  -30.8766,
  -30.9226,
  -30.9697,
  -31.0176,
  -31.066,
  -31.1141,
  -31.1612,
  -31.2071,
  -31.2518,
  -31.2955,
  -31.3377,
  -31.3811,
  -31.4255,
  -31.4712,
  -31.5182,
  -31.5662,
  -31.614,
  -31.661,
  -31.7063,
  -31.7497,
  -31.7917,
  -31.8325,
  -31.8729,
  -31.9133,
  -31.9545,
  -31.997,
  -32.0399,
  -32.0853,
  -32.1317,
  -32.1791,
  -32.2268,
  -32.2748,
  -32.3229,
  -32.3708,
  -32.4186,
  -32.4663,
  -32.5141,
  -32.5624,
  -32.6115,
  -32.6618,
  -32.7133,
  -32.7661,
  -32.8197,
  -32.8731,
  -32.9279,
  -32.983,
  -33.0385,
  -33.0943,
  -33.1498,
  -33.2043,
  -33.2574,
  -33.3093,
  -33.3605,
  -33.4112,
  -33.4619,
  -33.5122,
  -33.5618,
  -33.6101,
  -33.657,
  -33.7022,
  -33.7459,
  -33.7871,
  -33.828,
  -33.868,
  -33.9072,
  -33.946,
  -33.9844,
  -34.0223,
  -34.0592,
  -34.0942,
  -34.1265,
  -34.1556,
  -34.1813,
  -34.2042,
  -34.2246,
  -34.2433,
  -34.26,
  -34.2759,
  -34.2907,
  -34.3036,
  -34.3168,
  -34.3284,
  -34.3384,
  -34.3466,
  -34.353,
  -34.358,
  -34.3621,
  -34.3658,
  -34.3696,
  -34.3736,
  -34.3778,
  -34.3819,
  -34.3857,
  -34.3892,
  -34.3922,
  -34.3948,
  -34.3973,
  -34.4,
  -34.4032,
  -34.4068,
  -34.4132,
  -34.4218,
  -34.4321,
  -34.4436,
  -34.4554,
  -34.467,
  -34.4783,
  -34.4893,
  -34.5003,
  -34.5116,
  -34.524,
  -34.5379,
  -34.554,
  -34.5722,
  -34.5922,
  -34.6134,
  -34.6353,
  -34.6573,
  -34.6795,
  -34.702,
  -34.725,
  -34.7475,
  -34.7711,
  -34.7943,
  -34.8166,
  -34.8378,
  -34.8579,
  -34.8777,
  -34.8978,
  -34.9187,
  -34.9412,
  -34.9653,
  -34.9911,
  -35.0184,
  -35.0466,
  -35.075,
  -35.1029,
  -35.1296,
  -35.155,
  -35.1799,
  -35.2053,
  -35.2322,
  -35.261,
  -35.2914,
  -35.323,
  -35.3538,
  -35.3854,
  -35.4165,
  -35.4473,
  -35.4783,
  -35.5097,
  -35.5424,
  -35.5766,
  -35.6128,
  -35.6513,
  -35.6924,
  -35.7364,
  -35.7833,
  -35.8329,
  -35.8848,
  -35.9384,
  -35.9932,
  -36.0488,
  -36.1049,
  -36.1611,
  -36.2167,
  -36.271,
  -36.3234,
  -36.3736,
  -36.4212,
  -36.466,
  -36.508,
  -36.5466,
  -36.5844,
  -36.6218,
  -36.6595,
  -36.6975,
  -36.7356,
  -36.7731,
  -36.8095,
  -36.8446,
  -36.8784,
  -36.9109,
  -36.9425,
  -36.9735,
  -37.0036,
  -37.0327,
  -37.0604,
  -37.0868,
  -37.1118,
  -37.1357,
  -37.1581,
  -37.1786,
  -37.197,
  -37.2133,
  -37.2275,
  -37.2399,
  -37.2509,
  -37.2611,
  -37.2704,
  -37.2795,
  -37.2883,
  -37.2969,
  -37.3042,
  -37.3122,
  -37.3197,
  -37.3266,
  -37.3329,
  -37.3386,
  -37.3437,
  -37.3482,
  -37.3521,
  -37.3553,
  -37.3582,
  -37.3613,
  -37.3651,
  -37.3697,
  -37.3751,
  -37.3809,
  -37.3864,
  -37.3913,
  -37.3949,
  -37.3968,
  -37.3965,
  -37.3938,
  -37.389,
  -37.3826,
  -37.3752,
  -37.3676,
  -37.3603,
  -37.3535,
  -37.3476,
  -37.3427,
  -37.3391,
  -37.3373,
  -37.337,
  -37.3382,
  -37.3407,
  -37.3442,
  -37.3485,
  -37.3523,
  -37.357,
  -37.3607,
  -37.3625,
  -37.3616,
  -37.3579,
  -37.3516,
  -37.343,
  -37.3326,
  -37.3206,
  -37.3074,
  -37.2933,
  -37.2784,
  -37.2627,
  -37.2457,
  -37.2266,
  -37.2044,
  -37.1786,
  -37.1494,
  -37.1167,
  -37.0806,
  -37.0414,
  -36.9993,
  -36.9548,
  -36.9086,
  -36.8616,
  -29.2978,
  -29.336,
  -29.3756,
  -29.4166,
  -29.4586,
  -29.5013,
  -29.5444,
  -29.5876,
  -29.6308,
  -29.674,
  -29.7161,
  -29.7592,
  -29.8025,
  -29.8464,
  -29.8911,
  -29.9364,
  -29.982,
  -30.0276,
  -30.0729,
  -30.118,
  -30.1633,
  -30.2091,
  -30.2556,
  -30.303,
  -30.3513,
  -30.3994,
  -30.4492,
  -30.4991,
  -30.5487,
  -30.5975,
  -30.6449,
  -30.6912,
  -30.7366,
  -30.7813,
  -30.826,
  -30.8713,
  -30.9176,
  -30.9651,
  -31.0138,
  -31.063,
  -31.1108,
  -31.1583,
  -31.2043,
  -31.2485,
  -31.2914,
  -31.3335,
  -31.3758,
  -31.4191,
  -31.4643,
  -31.5108,
  -31.5586,
  -31.6067,
  -31.6538,
  -31.6995,
  -31.7433,
  -31.7854,
  -31.8251,
  -31.8652,
  -31.9052,
  -31.9459,
  -31.9877,
  -32.0309,
  -32.0755,
  -32.1215,
  -32.1684,
  -32.2159,
  -32.2637,
  -32.3113,
  -32.359,
  -32.4063,
  -32.4536,
  -32.501,
  -32.548,
  -32.597,
  -32.6475,
  -32.6994,
  -32.7531,
  -32.8075,
  -32.8629,
  -32.9186,
  -32.9742,
  -33.0301,
  -33.0859,
  -33.1413,
  -33.1959,
  -33.2489,
  -33.3009,
  -33.3519,
  -33.4027,
  -33.4534,
  -33.5028,
  -33.5526,
  -33.6013,
  -33.6482,
  -33.6934,
  -33.7366,
  -33.7784,
  -33.819,
  -33.8586,
  -33.8976,
  -33.9364,
  -33.9749,
  -34.0129,
  -34.0498,
  -34.0848,
  -34.1171,
  -34.146,
  -34.1716,
  -34.1933,
  -34.2136,
  -34.232,
  -34.2484,
  -34.2636,
  -34.2777,
  -34.2913,
  -34.3036,
  -34.3146,
  -34.3237,
  -34.3308,
  -34.3361,
  -34.3399,
  -34.3427,
  -34.3449,
  -34.3472,
  -34.35,
  -34.353,
  -34.3559,
  -34.3585,
  -34.3596,
  -34.361,
  -34.3618,
  -34.3622,
  -34.3629,
  -34.3644,
  -34.3675,
  -34.3728,
  -34.3804,
  -34.39,
  -34.4005,
  -34.4112,
  -34.4217,
  -34.4319,
  -34.4421,
  -34.4523,
  -34.4631,
  -34.4753,
  -34.4891,
  -34.5052,
  -34.5235,
  -34.5425,
  -34.5635,
  -34.585,
  -34.6067,
  -34.6285,
  -34.6508,
  -34.6737,
  -34.6971,
  -34.7204,
  -34.7432,
  -34.7652,
  -34.7859,
  -34.8058,
  -34.8254,
  -34.8452,
  -34.866,
  -34.8883,
  -34.9123,
  -34.9381,
  -34.9654,
  -34.9938,
  -35.0224,
  -35.0504,
  -35.0763,
  -35.1021,
  -35.1272,
  -35.1528,
  -35.1799,
  -35.2088,
  -35.2396,
  -35.2718,
  -35.3047,
  -35.3373,
  -35.37,
  -35.4023,
  -35.4349,
  -35.4681,
  -35.5024,
  -35.5383,
  -35.5761,
  -35.6162,
  -35.6587,
  -35.704,
  -35.7521,
  -35.8026,
  -35.855,
  -35.9088,
  -35.9633,
  -36.0184,
  -36.073,
  -36.1287,
  -36.1839,
  -36.238,
  -36.2902,
  -36.3401,
  -36.3872,
  -36.4313,
  -36.4729,
  -36.5121,
  -36.55,
  -36.5876,
  -36.6255,
  -36.6637,
  -36.7016,
  -36.7386,
  -36.7742,
  -36.8082,
  -36.8405,
  -36.8715,
  -36.9018,
  -36.9315,
  -36.9607,
  -36.9894,
  -37.0171,
  -37.0436,
  -37.0689,
  -37.093,
  -37.1156,
  -37.1355,
  -37.1544,
  -37.1711,
  -37.1857,
  -37.1983,
  -37.209,
  -37.2182,
  -37.2262,
  -37.2338,
  -37.241,
  -37.2483,
  -37.2558,
  -37.2633,
  -37.2709,
  -37.2779,
  -37.2844,
  -37.2902,
  -37.2952,
  -37.2994,
  -37.303,
  -37.3057,
  -37.3083,
  -37.3114,
  -37.3153,
  -37.3203,
  -37.3262,
  -37.3323,
  -37.3379,
  -37.3424,
  -37.3453,
  -37.3464,
  -37.3453,
  -37.3419,
  -37.3365,
  -37.3295,
  -37.3216,
  -37.3126,
  -37.305,
  -37.2982,
  -37.2924,
  -37.2876,
  -37.284,
  -37.2822,
  -37.2818,
  -37.283,
  -37.2854,
  -37.2888,
  -37.293,
  -37.2976,
  -37.3024,
  -37.3064,
  -37.3088,
  -37.309,
  -37.3067,
  -37.3021,
  -37.2956,
  -37.2874,
  -37.2777,
  -37.2666,
  -37.2543,
  -37.241,
  -37.2264,
  -37.2105,
  -37.1923,
  -37.1714,
  -37.147,
  -37.1194,
  -37.0885,
  -37.0543,
  -37.0169,
  -36.9764,
  -36.9332,
  -36.888,
  -36.8415,
  -29.2936,
  -29.3314,
  -29.371,
  -29.4121,
  -29.454,
  -29.4965,
  -29.5382,
  -29.5807,
  -29.6233,
  -29.666,
  -29.709,
  -29.7522,
  -29.7956,
  -29.8397,
  -29.8846,
  -29.9301,
  -29.976,
  -30.0219,
  -30.0676,
  -30.1131,
  -30.158,
  -30.2043,
  -30.2515,
  -30.2996,
  -30.3485,
  -30.3981,
  -30.4482,
  -30.4983,
  -30.5479,
  -30.5963,
  -30.6433,
  -30.6891,
  -30.7339,
  -30.7784,
  -30.8231,
  -30.8675,
  -30.9141,
  -30.9621,
  -31.0113,
  -31.0609,
  -31.1101,
  -31.1578,
  -31.2036,
  -31.2474,
  -31.2896,
  -31.3309,
  -31.3724,
  -31.4152,
  -31.4594,
  -31.5058,
  -31.5531,
  -31.5999,
  -31.6471,
  -31.693,
  -31.7369,
  -31.779,
  -31.8197,
  -31.8595,
  -31.8992,
  -31.9393,
  -31.9807,
  -32.0233,
  -32.0674,
  -32.1128,
  -32.1593,
  -32.2063,
  -32.2535,
  -32.2999,
  -32.3471,
  -32.3942,
  -32.4414,
  -32.4888,
  -32.5369,
  -32.586,
  -32.6366,
  -32.6891,
  -32.7433,
  -32.799,
  -32.8549,
  -32.911,
  -32.9671,
  -33.023,
  -33.0787,
  -33.134,
  -33.1875,
  -33.2407,
  -33.2927,
  -33.3436,
  -33.3943,
  -33.4449,
  -33.4954,
  -33.5454,
  -33.5942,
  -33.6411,
  -33.6861,
  -33.7288,
  -33.7702,
  -33.8103,
  -33.8494,
  -33.8882,
  -33.9269,
  -33.9653,
  -34.0023,
  -34.0391,
  -34.074,
  -34.1062,
  -34.1349,
  -34.1604,
  -34.1828,
  -34.2028,
  -34.2205,
  -34.2367,
  -34.2515,
  -34.2652,
  -34.2783,
  -34.2901,
  -34.3003,
  -34.3087,
  -34.3151,
  -34.3193,
  -34.3221,
  -34.3238,
  -34.3236,
  -34.3246,
  -34.3259,
  -34.3277,
  -34.3296,
  -34.3313,
  -34.3321,
  -34.3321,
  -34.3312,
  -34.3297,
  -34.3283,
  -34.3278,
  -34.3292,
  -34.3332,
  -34.3397,
  -34.3482,
  -34.3577,
  -34.3674,
  -34.377,
  -34.3863,
  -34.3948,
  -34.4046,
  -34.4151,
  -34.427,
  -34.4408,
  -34.4569,
  -34.475,
  -34.4948,
  -34.5154,
  -34.5364,
  -34.5577,
  -34.5793,
  -34.6014,
  -34.6243,
  -34.6476,
  -34.6706,
  -34.693,
  -34.7147,
  -34.7351,
  -34.7548,
  -34.7741,
  -34.7938,
  -34.8144,
  -34.8356,
  -34.8595,
  -34.8853,
  -34.9127,
  -34.941,
  -34.9695,
  -34.9975,
  -35.0245,
  -35.0503,
  -35.0757,
  -35.1016,
  -35.1288,
  -35.1579,
  -35.1889,
  -35.2216,
  -35.2552,
  -35.2891,
  -35.3234,
  -35.3577,
  -35.3922,
  -35.4272,
  -35.4633,
  -35.5009,
  -35.5404,
  -35.582,
  -35.625,
  -35.6715,
  -35.7206,
  -35.7719,
  -35.8248,
  -35.8787,
  -35.9332,
  -35.9881,
  -36.0433,
  -36.0986,
  -36.1535,
  -36.2073,
  -36.2591,
  -36.3084,
  -36.3549,
  -36.3984,
  -36.4392,
  -36.4781,
  -36.5161,
  -36.5538,
  -36.5918,
  -36.6298,
  -36.6673,
  -36.7037,
  -36.7384,
  -36.7712,
  -36.8021,
  -36.8316,
  -36.8593,
  -36.8876,
  -36.9158,
  -36.9439,
  -36.9715,
  -36.9981,
  -37.0234,
  -37.0474,
  -37.0699,
  -37.0911,
  -37.1102,
  -37.1274,
  -37.1425,
  -37.1555,
  -37.1662,
  -37.1749,
  -37.1822,
  -37.1886,
  -37.1946,
  -37.2007,
  -37.2073,
  -37.2144,
  -37.2218,
  -37.229,
  -37.2357,
  -37.2414,
  -37.2462,
  -37.25,
  -37.2533,
  -37.2556,
  -37.258,
  -37.2611,
  -37.2651,
  -37.2694,
  -37.2757,
  -37.282,
  -37.2877,
  -37.2922,
  -37.2948,
  -37.2955,
  -37.2939,
  -37.2899,
  -37.2839,
  -37.2763,
  -37.2679,
  -37.2595,
  -37.2519,
  -37.2454,
  -37.2398,
  -37.2353,
  -37.2319,
  -37.23,
  -37.2295,
  -37.2304,
  -37.2324,
  -37.2355,
  -37.2394,
  -37.244,
  -37.2487,
  -37.253,
  -37.2561,
  -37.2573,
  -37.2562,
  -37.2532,
  -37.2485,
  -37.2423,
  -37.2345,
  -37.2253,
  -37.2146,
  -37.2025,
  -37.1893,
  -37.1745,
  -37.1573,
  -37.1376,
  -37.1148,
  -37.0876,
  -37.0585,
  -37.026,
  -36.9902,
  -36.9515,
  -36.9098,
  -36.8657,
  -36.8197 ;
    } // group puerto_rico_virgin_islands_geoid18
  } // group puerto_rico_virgin_islands_geoid18
}

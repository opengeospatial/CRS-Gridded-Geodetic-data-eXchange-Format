netcdf nzgd2000-20180701 {

// global attributes:
		:Conventions = "GGXF-1.0, ACDD-1.3" ;
		:source_file = "nzgd2000-20180701.ggxf" ;
		:product_version = "20180701" ;
		:content = "deformationModel" ;
		:title = "New Zealand Deformation Model." ;
		:summary = "Defines the secular model (National Deformation Model)\nand patches for significant deformation events since 2000.\n" ;
		:institution = "Land Information New Zealand" ;
		:deliveryPoint = "Level 7, Radio New Zealand House\n155 The Terrace\nPO Box 5501\n" ;
		:city = "Wellington" ;
		:postalCode = "6145" ;
		:creator_email = "customersupport@linz.govt.nz" ;
		:publisher_url = "https://www.linz.govt.nz/nzgd2000" ;
		:date_issued = "2018-07-01" ;
		:extent_description = "New Zealand EEZ" ;
		:geospatial_lat_min = -55.94 ;
		:geospatial_lon_min = 160.62 ;
		:geospatial_lat_max = -25.89 ;
		:geospatial_lon_max = -171.23 ;
		:geospatial_bounds = "Polygon ((-32.42 168.65, -34.98 168.10, -37.58 170.07, -40.60 167.30,  -44.32 162.17, -51.17 160.62, -54.97 165.11, -55.94 168.78, -54.70 173.54, -53.26 174.64, -51.66 174.48, -53.04 178.46, -51.94 182.69, -50.45 183.84, -47.76 184.00, -46.81 187.31, -44.68 188.77, -42.93 188.53, -41.50 187.23, -40.26 182.07, -36.91 182.64, -34.59 180.22, -34.45 182.66, -33.12 184.50, -29.73 185.92, -27.47 185.34, -25.89 182.29, -27.22 179.01, -31.55 177.28, -34.32 179.37, -30.85 172.97, -30.88 171.22, -32.42 168.65))" ;
		:sourceCrsWkt = "GEOGCRS[\"NZGD2000\",DATUM[\"New Zealand Geodetic Datum 2000\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6167]],CS[ellipsoidal,3,ID[\"EPSG\",6423]],AXIS[\"Geodetic latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Geodetic longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],ID[\"EPSG\",4959]]" ;
		:targetCrsWkt = "GEOGCRS[\"ITRF96\", DYNAMIC[FRAMEEPOCH[1997.0]],DATUM[\"International Terrestrial Reference Frame 1996\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6654]],CS[ellipsoidal,3,ID[\"EPSG\",6423]],AXIS[\"Geodetic latitude (Lat)\",north,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Geodetic longitude (Lon)\",east,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]]],AXIS[\"Ellipsoidal height (h)\",up,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],ID[\"EPSG\",7907]]" ;
		:interpolationCrsWkt = "GEOGCRS[\"NZGD2000\",DATUM[\"New Zealand Geodetic Datum 2000\",ELLIPSOID[\"GRS 1980\",6378137,298.2572221,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]],ID[\"EPSG\",7019]],ID[\"EPSG\",6167]],CS[ellipsoidal,2,ID[\"EPSG\",6422]],AXIS[\"Geodetic latitude (Lat)\",north],AXIS[\"Geodetic longitude (Lon)\",east],ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9102]],ID[\"EPSG\",4167]]" ;
		:parameters.count = 3LL ;
		:parameters.0.parameterName = "displacementEast" ;
		:parameters.0.parameterSet = "displacement" ;
		:parameters.0.unitName = "metre" ;
		:parameters.0.unitSiRatio = 1. ;
		:parameters.0.sourceCrsAxis = 1LL ;
		:parameters.1.parameterName = "displacementNorth" ;
		:parameters.1.parameterSet = "displacement" ;
		:parameters.1.unitName = "metre" ;
		:parameters.1.unitSiRatio = 1. ;
		:parameters.1.sourceCrsAxis = 0LL ;
		:parameters.2.parameterName = "displacementUp" ;
		:parameters.2.parameterSet = "displacement" ;
		:parameters.2.unitName = "metre" ;
		:parameters.2.unitSiRatio = 1. ;
		:parameters.2.sourceCrsAxis = 2LL ;
		:operationAccuracy = 0.01 ;

group: nz_linz_nzgd2000-ndm-grid02 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Secular deformation model derived from NUVEL-1A rotation rates\nSecular deformation model derived from GNS model 2011 V4\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "velocity" ;
  		:timeFunctions.0.functionReferenceDate = "2000-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: ndm_grid_nuvel1a_eez {
    dimensions:
    	iNodeCount = 73 ;
    	jNodeCount = 67 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -25., 0., -0.5, 158., 0.5, 0. ;

    group: ndm_grid_igns2011_nz {
      dimensions:
      	iNodeCount = 141 ;
      	jNodeCount = 151 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -33., 0., -0.1, 165.5, 0.1, 0. ;
      } // group ndm_grid_igns2011_nz
    } // group ndm_grid_nuvel1a_eez
  } // group nz_linz_nzgd2000-ndm-grid02

group: nz_linz_nzgd2000-si20030821-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Secretary Island (Fiordland) earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2003-08-21T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2004-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_si_20030821_grid_si_l1 {
    dimensions:
    	iNodeCount = 44 ;
    	jNodeCount = 34 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -43.5, 0., -0.125, 165.85, 0.15, 0. ;

    group: patch_si_20030821_grid_si_l2 {
      dimensions:
      	iNodeCount = 47 ;
      	jNodeCount = 45 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -44.5, 0., -0.03125, 166.225, 0.0375, 0. ;

      group: patch_si_20030821_grid_si_l3 {
        dimensions:
        	iNodeCount = 93 ;
        	jNodeCount = 81 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -44.828125, 0., -0.0078125, 166.5625, 0.009375, 0. ;
        } // group patch_si_20030821_grid_si_l3
      } // group patch_si_20030821_grid_si_l2
    } // group patch_si_20030821_grid_si_l1
  } // group nz_linz_nzgd2000-si20030821-grid01

group: nz_linz_nzgd2000-mq20041223-grid011 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p0_l1 {
    dimensions:
    	iNodeCount = 10 ;
    	jNodeCount = 8 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -52.125, 0., -0.125, 168.4, 0.15, 0. ;
    } // group patch_mq_20041223_grid_mq_p0_l1
  } // group nz_linz_nzgd2000-mq20041223-grid011

group: nz_linz_nzgd2000-mq20041223-grid012 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p1_sl2 {
    dimensions:
    	iNodeCount = 105 ;
    	jNodeCount = 137 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -48.25, 0., -0.03125, 158.8, 0.0375, 0. ;
    } // group patch_mq_20041223_grid_mq_p1_sl2
  } // group nz_linz_nzgd2000-mq20041223-grid012

group: nz_linz_nzgd2000-mq20041223-grid013 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p2_l1 {
    dimensions:
    	iNodeCount = 11 ;
    	jNodeCount = 11 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -50.125, 0., -0.125, 165.4, 0.15, 0. ;
    } // group patch_mq_20041223_grid_mq_p2_l1
  } // group nz_linz_nzgd2000-mq20041223-grid013

group: nz_linz_nzgd2000-mq20041223-grid014 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p3_l1 {
    dimensions:
    	iNodeCount = 9 ;
    	jNodeCount = 8 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -49.25, 0., -0.125, 178.15, 0.15, 0. ;
    } // group patch_mq_20041223_grid_mq_p3_l1
  } // group nz_linz_nzgd2000-mq20041223-grid014

group: nz_linz_nzgd2000-mq20041223-grid015 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p4_l1 {
    dimensions:
    	iNodeCount = 70 ;
    	jNodeCount = 68 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.125, 0., -0.125, 165.85, 0.15, 0. ;
    } // group patch_mq_20041223_grid_mq_p4_l1
  } // group nz_linz_nzgd2000-mq20041223-grid015

group: nz_linz_nzgd2000-mq20041223-grid016 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Macquarie Plate earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2004-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2005-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_mq_20041223_grid_mq_p5_l1 {
    dimensions:
    	iNodeCount = 8 ;
    	jNodeCount = 7 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -47.375, 0., -0.125, 178.45, 0.15, 0. ;
    } // group patch_mq_20041223_grid_mq_p5_l1
  } // group nz_linz_nzgd2000-mq20041223-grid016

group: nz_linz_nzgd2000-gs20071016-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Fiordland (George Sound) earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2007-10-16T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2008-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_gs_20071016_grid_gs_l1 {
    dimensions:
    	iNodeCount = 37 ;
    	jNodeCount = 27 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -43.75, 0., -0.125, 165.85, 0.15, 0. ;

    group: patch_gs_20071016_grid_gs_l2 {
      dimensions:
      	iNodeCount = 45 ;
      	jNodeCount = 37 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -44.28125, 0., -0.03125, 166.6375, 0.0375, 0. ;

      group: patch_gs_20071016_grid_gs_l3 {
        dimensions:
        	iNodeCount = 54 ;
        	jNodeCount = 52 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -44.6171875, 0., -0.0078125, 167.0875, 0.009375, 0. ;
        } // group patch_gs_20071016_grid_gs_l3
      } // group patch_gs_20071016_grid_gs_l2
    } // group patch_gs_20071016_grid_gs_l1
  } // group nz_linz_nzgd2000-gs20071016-grid01

group: nz_linz_nzgd2000-ds20090715-grid011 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1.05 ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p0_l1 {
    dimensions:
    	iNodeCount = 11 ;
    	jNodeCount = 11 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -50.125, 0., -0.125, 165.4, 0.15, 0. ;
    } // group patch_ds_20090715_grid_ds_p0_l1
  } // group nz_linz_nzgd2000-ds20090715-grid011

group: nz_linz_nzgd2000-ds20090715-grid012 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1.05 ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p1_l1 {
    dimensions:
    	iNodeCount = 6 ;
    	jNodeCount = 7 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -49.25, 0., -0.125, 178.15, 0.15, 0. ;
    } // group patch_ds_20090715_grid_ds_p1_l1
  } // group nz_linz_nzgd2000-ds20090715-grid012

group: nz_linz_nzgd2000-ds20090715-grid013 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1.05 ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p2_l1 {
    dimensions:
    	iNodeCount = 85 ;
    	jNodeCount = 72 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39.625, 0., -0.125, 164.65, 0.15, 0. ;

    group: patch_ds_20090715_grid_ds_p2_l2 {
      dimensions:
      	iNodeCount = 67 ;
      	jNodeCount = 73 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -44.6875, 0., -0.03125, 165.2875, 0.0375, 0. ;

      group: patch_ds_20090715_grid_ds_p2_l3 {
        dimensions:
        	iNodeCount = 83 ;
        	jNodeCount = 138 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -45.28125, 0., -0.0078125, 166.075, 0.009375, 0. ;
        } // group patch_ds_20090715_grid_ds_p2_l3
      } // group patch_ds_20090715_grid_ds_p2_l2
    } // group patch_ds_20090715_grid_ds_p2_l1
  } // group nz_linz_nzgd2000-ds20090715-grid013

group: nz_linz_nzgd2000-ds20090715-grid014 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Dusky Sound (Fiordland) earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 2LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1.05 ;
  		:timeFunctions.1.functionType = "ramp" ;
  		:timeFunctions.1.startDate = "2009-07-15T00:00:00Z" ;
  		:timeFunctions.1.endDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.functionReferenceDate = "2011-09-01T00:00:00Z" ;
  		:timeFunctions.1.scaleFactor = 0.29 ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ds_20090715_grid_ds_p3_l1 {
    dimensions:
    	iNodeCount = 8 ;
    	jNodeCount = 7 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -47.375, 0., -0.125, 178.45, 0.15, 0. ;
    } // group patch_ds_20090715_grid_ds_p3_l1
  } // group nz_linz_nzgd2000-ds20090715-grid014

group: nz_linz_nzgd2000-c120100904-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Darfield earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2010-09-04T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2011-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c1_20100904_grid_c1_l1 {
    dimensions:
    	iNodeCount = 55 ;
    	jNodeCount = 52 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.375, 0., -0.125, 168.1, 0.15, 0. ;

    group: patch_c1_20100904_grid_c1_l2 {
      dimensions:
      	iNodeCount = 59 ;
      	jNodeCount = 50 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.8125, 0., -0.03125, 171.1, 0.0375, 0. ;

      group: patch_c1_20100904_grid_c1_l3 {
        dimensions:
        	iNodeCount = 118 ;
        	jNodeCount = 84 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.25, 0., -0.0078125, 171.625, 0.009375, 0. ;

        group: patch_c1_20100904_grid_c1_l4 {
          dimensions:
          	iNodeCount = 306 ;
          	jNodeCount = 141 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.423828125, 0., -0.001953125, 171.8125, 0.00234375, 0. ;
          } // group patch_c1_20100904_grid_c1_l4
        } // group patch_c1_20100904_grid_c1_l3
      } // group patch_c1_20100904_grid_c1_l2
    } // group patch_c1_20100904_grid_c1_l1
  } // group nz_linz_nzgd2000-c120100904-grid01

group: nz_linz_nzgd2000-c220110222-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Christchurch February earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2011-02-22T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2012-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c2_20110222_grid_c2_l1 {
    dimensions:
    	iNodeCount = 21 ;
    	jNodeCount = 18 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.375, 0., -0.125, 170.8, 0.15, 0. ;

    group: patch_c2_20110222_grid_c2_l2 {
      dimensions:
      	iNodeCount = 38 ;
      	jNodeCount = 34 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.03125, 0., -0.03125, 172., 0.0375, 0. ;

      group: patch_c2_20110222_grid_c2_l3 {
        dimensions:
        	iNodeCount = 62 ;
        	jNodeCount = 52 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.3515625, 0., -0.0078125, 172.4125, 0.009375, 0. ;

        group: patch_c2_20110222_grid_c2_l4 {
          dimensions:
          	iNodeCount = 118 ;
          	jNodeCount = 81 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.474609375, 0., -0.001953125, 172.56015625, 0.00234375, 0. ;
          } // group patch_c2_20110222_grid_c2_l4
        } // group patch_c2_20110222_grid_c2_l3
      } // group patch_c2_20110222_grid_c2_l2
    } // group patch_c2_20110222_grid_c2_l1
  } // group nz_linz_nzgd2000-c220110222-grid01

group: nz_linz_nzgd2000-c320110613-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Christchurch June earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2011-06-13T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2012-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c3_20110613_grid_c3_l1 {
    dimensions:
    	iNodeCount = 16 ;
    	jNodeCount = 15 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.625, 0., -0.125, 171.4, 0.15, 0. ;

    group: patch_c3_20110613_grid_c3_l2 {
      dimensions:
      	iNodeCount = 33 ;
      	jNodeCount = 31 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.09375, 0., -0.03125, 172.15, 0.0375, 0. ;

      group: patch_c3_20110613_grid_c3_l3 {
        dimensions:
        	iNodeCount = 51 ;
        	jNodeCount = 48 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.375, 0., -0.0078125, 172.515625, 0.009375, 0. ;

        group: patch_c3_20110613_grid_c3_l4 {
          dimensions:
          	iNodeCount = 88 ;
          	jNodeCount = 84 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.484375, 0., -0.001953125, 172.65390625, 0.00234375, 0. ;
          } // group patch_c3_20110613_grid_c3_l4
        } // group patch_c3_20110613_grid_c3_l3
      } // group patch_c3_20110613_grid_c3_l2
    } // group patch_c3_20110613_grid_c3_l1
  } // group nz_linz_nzgd2000-c320110613-grid01

group: nz_linz_nzgd2000-c420111223-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Christchurch earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2011-12-23T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2012-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_c4_20111223_grid_c4_l1 {
    dimensions:
    	iNodeCount = 15 ;
    	jNodeCount = 13 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.75, 0., -0.125, 171.55, 0.15, 0. ;

    group: patch_c4_20111223_grid_c4_l2 {
      dimensions:
      	iNodeCount = 32 ;
      	jNodeCount = 30 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.03125, 0., -0.03125, 172.1875, 0.0375, 0. ;

      group: patch_c4_20111223_grid_c4_l3 {
        dimensions:
        	iNodeCount = 52 ;
        	jNodeCount = 44 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.3125, 0., -0.0078125, 172.553125, 0.009375, 0. ;

        group: patch_c4_20111223_grid_c4_l4 {
          dimensions:
          	iNodeCount = 87 ;
          	jNodeCount = 61 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.421875, 0., -0.001953125, 172.67734375, 0.00234375, 0. ;
          } // group patch_c4_20111223_grid_c4_l4
        } // group patch_c4_20111223_grid_c4_l3
      } // group patch_c4_20111223_grid_c4_l2
    } // group patch_c4_20111223_grid_c4_l1
  } // group nz_linz_nzgd2000-c420111223-grid01

group: nz_linz_nzgd2000-cs20130721-grid02 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Mw 6.6 Cook Strait earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2013-07-21T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2014-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_cs_20130721_grid_cs_20130721_l1 {
    dimensions:
    	iNodeCount = 34 ;
    	jNodeCount = 32 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39.5, 0., -0.125, 171.55, 0.15, 0. ;

    group: patch_cs_20130721_grid_cs_20130721_l2 {
      dimensions:
      	iNodeCount = 43 ;
      	jNodeCount = 37 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.03125, 0., -0.03125, 173.5375, 0.0375, 0. ;

      group: patch_cs_20130721_grid_cs_20130721_l3 {
        dimensions:
        	iNodeCount = 73 ;
        	jNodeCount = 57 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.3828125, 0., -0.0078125, 173.9875, 0.009375, 0. ;

        group: patch_cs_20130721_grid_cs_20130721_l4 {
          dimensions:
          	iNodeCount = 90 ;
          	jNodeCount = 68 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.537109375, 0., -0.001953125, 174.28984375, 0.00234375, 0. ;
          } // group patch_cs_20130721_grid_cs_20130721_l4
        } // group patch_cs_20130721_grid_cs_20130721_l3
      } // group patch_cs_20130721_grid_cs_20130721_l2
    } // group patch_cs_20130721_grid_cs_20130721_l1
  } // group nz_linz_nzgd2000-cs20130721-grid02

group: nz_linz_nzgd2000-lg20130816-grid02 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Mw 6.6 Lake Grassmere earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2013-08-16T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2014-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_lg_20130816_grid_lg_20130816_l1 {
    dimensions:
    	iNodeCount = 39 ;
    	jNodeCount = 39 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39.25, 0., -0.125, 170.95, 0.15, 0. ;

    group: patch_lg_20130816_grid_lg_20130816_l2 {
      dimensions:
      	iNodeCount = 44 ;
      	jNodeCount = 40 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.09375, 0., -0.03125, 173.3875, 0.0375, 0. ;

      group: patch_lg_20130816_grid_lg_20130816_l3 {
        dimensions:
        	iNodeCount = 79 ;
        	jNodeCount = 63 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.4609375, 0., -0.0078125, 173.809375, 0.009375, 0. ;

        group: patch_lg_20130816_grid_lg_20130816_l4 {
          dimensions:
          	iNodeCount = 134 ;
          	jNodeCount = 104 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.60546875, 0., -0.001953125, 174.034375, 0.00234375, 0. ;
          } // group patch_lg_20130816_grid_lg_20130816_l4
        } // group patch_lg_20130816_grid_lg_20130816_l3
      } // group patch_lg_20130816_grid_lg_20130816_l2
    } // group patch_lg_20130816_grid_lg_20130816_l1
  } // group nz_linz_nzgd2000-lg20130816-grid02

group: nz_linz_nzgd2000-ch20160214-grid01 {
  dimensions:
  	displacementCount = 3 ;

  // group attributes:
  		:comment = "Christchurch Valentines Day earthquake" ;
  		string :gridParameters = "displacementEast", "displacementNorth", "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-02-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ch_20160214_grid_ch_20160214_l1 {
    dimensions:
    	iNodeCount = 14 ;
    	jNodeCount = 11 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -42.875, 0., -0.125, 171.7, 0.15, 0. ;

    group: patch_ch_20160214_grid_ch_20160214_l2 {
      dimensions:
      	iNodeCount = 29 ;
      	jNodeCount = 27 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -43.0625, 0., -0.03125, 172.225, 0.0375, 0. ;

      group: patch_ch_20160214_grid_ch_20160214_l3 {
        dimensions:
        	iNodeCount = 46 ;
        	jNodeCount = 38 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -43.3203125, 0., -0.0078125, 172.553125, 0.009375, 0. ;

        group: patch_ch_20160214_grid_ch_20160214_l4 {
          dimensions:
          	iNodeCount = 79 ;
          	jNodeCount = 61 ;
          variables:
          	float displacement(iNodeCount, jNodeCount, displacementCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -43.408203125, 0., -0.001953125, 172.67265625, 0.00234375, 0. ;
          } // group patch_ch_20160214_grid_ch_20160214_l4
        } // group patch_ch_20160214_grid_ch_20160214_l3
      } // group patch_ch_20160214_grid_ch_20160214_l2
    } // group patch_ch_20160214_grid_ch_20160214_l1
  } // group nz_linz_nzgd2000-ch20160214-grid01

group: nz_linz_nzgd2000-ka20161114-grid01 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-11-14T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114co_h_l1_f {
    dimensions:
    	iNodeCount = 89 ;
    	jNodeCount = 110 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -34., 0., -0.125, 165.85, 0.15, 0. ;

    group: patch_ka_20161114_grid_ka_20161114co_h_l2_f {
      dimensions:
      	iNodeCount = 95 ;
      	jNodeCount = 82 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -40.8125, 0., -0.03125, 171.925, 0.0375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114co_h_l2_f
    } // group patch_ka_20161114_grid_ka_20161114co_h_l1_f
  } // group nz_linz_nzgd2000-ka20161114-grid01

group: nz_linz_nzgd2000-ka20161114-grid02 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114co_h_l2_r {
    dimensions:
    	iNodeCount = 65 ;
    	jNodeCount = 53 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -41.28125, 0., -0.03125, 172.525, 0.0375, 0. ;

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_00 {
      dimensions:
      	iNodeCount = 115 ;
      	jNodeCount = 94 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.1484375, 0., -0.0078125, 172.571875, 0.009375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_00 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 107 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 172.7828125, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_00

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_01 {
        dimensions:
        	iNodeCount = 11 ;
        	jNodeCount = 26 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.435546875, 0., -0.001953125, 173.00546875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_01

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_02 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.02890625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_02

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_03 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 51 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.38671875, 0., -0.001953125, 173.02890625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_03

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_04 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 88 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.275, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_04

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_05 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.275, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_05

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_060 {
        dimensions:
        	iNodeCount = 21 ;
        	jNodeCount = 63 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.47421875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_060

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_080 {
        dimensions:
        	iNodeCount = 52 ;
        	jNodeCount = 30 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_080

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_090 {
        dimensions:
        	iNodeCount = 52 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_090

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_100 {
        dimensions:
        	iNodeCount = 52 ;
        	jNodeCount = 63 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_100
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_00

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_01 {
      dimensions:
      	iNodeCount = 53 ;
      	jNodeCount = 89 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.4609375, 0., -0.0078125, 173.153125, 0.009375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_061 {
        dimensions:
        	iNodeCount = 21 ;
        	jNodeCount = 49 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.47421875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_061

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_07 {
        dimensions:
        	iNodeCount = 9 ;
        	jNodeCount = 6 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.044921875, 0., -0.001953125, 173.50234375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_07

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_101 {
        dimensions:
        	iNodeCount = 52 ;
        	jNodeCount = 49 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_101

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_110 {
        dimensions:
        	iNodeCount = 52 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 173.52109375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_110
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_01

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_02 {
      dimensions:
      	iNodeCount = 73 ;
      	jNodeCount = 63 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.1484375, 0., -0.0078125, 173.640625, 0.009375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_081 {
        dimensions:
        	iNodeCount = 28 ;
        	jNodeCount = 30 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.484375, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_081

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_091 {
        dimensions:
        	iNodeCount = 55 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_091

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_102 {
        dimensions:
        	iNodeCount = 55 ;
        	jNodeCount = 63 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_102

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_13 {
        dimensions:
        	iNodeCount = 87 ;
        	jNodeCount = 95 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.26953125, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_13

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_140 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 63 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_140

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_170 {
        dimensions:
        	iNodeCount = 62 ;
        	jNodeCount = 41 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1484375, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_170
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_02

    group: patch_ka_20161114_grid_ka_20161114co_h_l3_r_03 {
      dimensions:
      	iNodeCount = 114 ;
      	jNodeCount = 94 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.421875, 0., -0.0078125, 173.640625, 0.009375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_103 {
        dimensions:
        	iNodeCount = 55 ;
        	jNodeCount = 49 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_103

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_111 {
        dimensions:
        	iNodeCount = 55 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 173.640625, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_111

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_12 {
        dimensions:
        	iNodeCount = 15 ;
        	jNodeCount = 10 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.822265625, 0., -0.001953125, 173.734375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_12

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_141 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 49 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_141

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_15 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_15

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_16 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 41 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.76171875, 0., -0.001953125, 173.7671875, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_16

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_171 {
        dimensions:
        	iNodeCount = 62 ;
        	jNodeCount = 49 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_171

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_18 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 111 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_18

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_19 {
        dimensions:
        	iNodeCount = 106 ;
        	jNodeCount = 93 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.66015625, 0., -0.001953125, 174.01328125, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_19

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_20 {
        dimensions:
        	iNodeCount = 59 ;
        	jNodeCount = 35 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.83984375, 0., -0.001953125, 174.259375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_20

      group: patch_ka_20161114_grid_ka_20161114co_h_l4_r_21 {
        dimensions:
        	iNodeCount = 104 ;
        	jNodeCount = 110 ;
        variables:
        	float displacement(iNodeCount, jNodeCount, displacementCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.626953125, 0., -0.001953125, 174.259375, 0.00234375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114co_h_l4_r_21
      } // group patch_ka_20161114_grid_ka_20161114co_h_l3_r_03
    } // group patch_ka_20161114_grid_ka_20161114co_h_l2_r
  } // group nz_linz_nzgd2000-ka20161114-grid02

group: nz_linz_nzgd2000-ka20161114-grid03 {

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		:gridParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114co_v_l1 {
    dimensions:
    	iNodeCount = 86 ;
    	jNodeCount = 108 ;
    variables:
    	float displacement(iNodeCount, jNodeCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -34.25, 0., -0.125, 166.3, 0.15, 0. ;

    group: patch_ka_20161114_grid_ka_20161114co_v_l2 {
      dimensions:
      	iNodeCount = 74 ;
      	jNodeCount = 67 ;
      variables:
      	float displacement(iNodeCount, jNodeCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.0625, 0., -0.03125, 172.225, 0.0375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_00 {
        dimensions:
        	iNodeCount = 103 ;
        	jNodeCount = 89 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1171875, 0., -0.0078125, 172.65625, 0.009375, 0. ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_00 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 88 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.490234375, 0., -0.001953125, 172.79921875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_00

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_01 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 105 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.03828125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_01

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_02 {
          dimensions:
          	iNodeCount = 89 ;
          	jNodeCount = 52 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.353515625, 0., -0.001953125, 173.07109375, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_02

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_03 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 100 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.27734375, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_03

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_04 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 89 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.28125, 0., -0.001953125, 173.27734375, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_04

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_050 {
          dimensions:
          	iNodeCount = 21 ;
          	jNodeCount = 67 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.46953125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_050

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_060 {
          dimensions:
          	iNodeCount = 42 ;
          	jNodeCount = 34 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_060

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_070 {
          dimensions:
          	iNodeCount = 42 ;
          	jNodeCount = 107 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.24609375, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_070

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_080 {
          dimensions:
          	iNodeCount = 42 ;
          	jNodeCount = 67 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_080
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_00

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_01 {
        dimensions:
        	iNodeCount = 44 ;
        	jNodeCount = 70 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.578125, 0., -0.0078125, 173.209375, 0.009375, 0. ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_051 {
          dimensions:
          	iNodeCount = 21 ;
          	jNodeCount = 33 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0546875, 0., -0.001953125, 173.46953125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_051

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_081 {
          dimensions:
          	iNodeCount = 42 ;
          	jNodeCount = 41 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.51640625, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_081

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_090 {
          dimensions:
          	iNodeCount = 12 ;
          	jNodeCount = 66 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.912109375, 0., -0.001953125, 173.58671875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_090
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_01

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_02 {
        dimensions:
        	iNodeCount = 79 ;
        	jNodeCount = 60 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.1171875, 0., -0.0078125, 173.6125, 0.009375, 0. ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_061 {
          dimensions:
          	iNodeCount = 62 ;
          	jNodeCount = 34 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_061

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_071 {
          dimensions:
          	iNodeCount = 62 ;
          	jNodeCount = 107 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.24609375, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_071

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_082 {
          dimensions:
          	iNodeCount = 62 ;
          	jNodeCount = 67 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_082

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_10 {
          dimensions:
          	iNodeCount = 7 ;
          	jNodeCount = 4 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.453125, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_10

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_11 {
          dimensions:
          	iNodeCount = 93 ;
          	jNodeCount = 107 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.24609375, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_11

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_120 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 67 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_120

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_140 {
          dimensions:
          	iNodeCount = 40 ;
          	jNodeCount = 59 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.1171875, 0., -0.001953125, 173.99453125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_140
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_02

      group: patch_ka_20161114_grid_ka_20161114co_v_l3_03 {
        dimensions:
        	iNodeCount = 103 ;
        	jNodeCount = 88 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.4375, 0., -0.0078125, 173.6125, 0.009375, 0. ;

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_083 {
          dimensions:
          	iNodeCount = 62 ;
          	jNodeCount = 41 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_083

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_091 {
          dimensions:
          	iNodeCount = 62 ;
          	jNodeCount = 66 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.912109375, 0., -0.001953125, 173.6125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_091

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_121 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 41 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_121

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_13 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 93 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.859375, 0., -0.001953125, 173.75546875, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_13

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_141 {
          dimensions:
          	iNodeCount = 40 ;
          	jNodeCount = 41 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -42.0390625, 0., -0.001953125, 173.99453125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_141

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_15 {
          dimensions:
          	iNodeCount = 103 ;
          	jNodeCount = 107 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.83203125, 0., -0.001953125, 173.99453125, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_15

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_16 {
          dimensions:
          	iNodeCount = 64 ;
          	jNodeCount = 78 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.681640625, 0., -0.001953125, 174.0859375, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_16

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_17 {
          dimensions:
          	iNodeCount = 56 ;
          	jNodeCount = 45 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.83203125, 0., -0.001953125, 174.23359375, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_17

        group: patch_ka_20161114_grid_ka_20161114co_v_l4_18 {
          dimensions:
          	iNodeCount = 101 ;
          	jNodeCount = 106 ;
          variables:
          	float displacement(iNodeCount, jNodeCount) ;
          		displacement:_Storage = "contiguous" ;
          		displacement:_Endianness = "little" ;

          // group attributes:
          		:affineCoeffs = -41.626953125, 0., -0.001953125, 174.23359375, 0.00234375, 0. ;
          } // group patch_ka_20161114_grid_ka_20161114co_v_l4_18
        } // group patch_ka_20161114_grid_ka_20161114co_v_l3_03
      } // group patch_ka_20161114_grid_ka_20161114co_v_l2
    } // group patch_ka_20161114_grid_ka_20161114co_v_l1
  } // group nz_linz_nzgd2000-ka20161114-grid03

group: nz_linz_nzgd2000-ka20161114-grid04 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake postearthquake month 0-1,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe1_h_l1_f {
    dimensions:
    	iNodeCount = 46 ;
    	jNodeCount = 39 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -39., 0., -0.125, 169.6, 0.15, 0. ;

    group: patch_ka_20161114_grid_ka_20161114pe1_h_l2_f {
      dimensions:
      	iNodeCount = 74 ;
      	jNodeCount = 59 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.125, 0., -0.03125, 172.6375, 0.0375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114pe1_h_l2_f
    } // group patch_ka_20161114_grid_ka_20161114pe1_h_l1_f
  } // group nz_linz_nzgd2000-ka20161114-grid04

group: nz_linz_nzgd2000-ka20161114-grid05 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake postearthquake month 0-1,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe1_h_l2_r {
    dimensions:
    	iNodeCount = 67 ;
    	jNodeCount = 56 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -41.28125, 0., -0.03125, 172.45, 0.0375, 0. ;

    group: patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_00 {
      dimensions:
      	iNodeCount = 93 ;
      	jNodeCount = 83 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42.0546875, 0., -0.0078125, 172.834375, 0.009375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_00

    group: patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_01 {
      dimensions:
      	iNodeCount = 92 ;
      	jNodeCount = 125 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.5703125, 0., -0.0078125, 173.696875, 0.009375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114pe1_h_l3_r_01
    } // group patch_ka_20161114_grid_ka_20161114pe1_h_l2_r
  } // group nz_linz_nzgd2000-ka20161114-grid05

group: nz_linz_nzgd2000-ka20161114-grid06 {

  // group attributes:
  		:comment = "Event: Kaikoura earthquake postearthquake month 0-1,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		:gridParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe1_v_l1 {
    dimensions:
    	iNodeCount = 29 ;
    	jNodeCount = 27 ;
    variables:
    	float displacement(iNodeCount, jNodeCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.5, 0., -0.125, 171.85, 0.15, 0. ;

    group: patch_ka_20161114_grid_ka_20161114pe1_v_l2 {
      dimensions:
      	iNodeCount = 72 ;
      	jNodeCount = 74 ;
      variables:
      	float displacement(iNodeCount, jNodeCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -40.75, 0., -0.03125, 172.675, 0.0375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114pe1_v_l3_00 {
        dimensions:
        	iNodeCount = 92 ;
        	jNodeCount = 82 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0546875, 0., -0.0078125, 172.84375, 0.009375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114pe1_v_l3_00

      group: patch_ka_20161114_grid_ka_20161114pe1_v_l3_01 {
        dimensions:
        	iNodeCount = 91 ;
        	jNodeCount = 119 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.609375, 0., -0.0078125, 173.696875, 0.009375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114pe1_v_l3_01
      } // group patch_ka_20161114_grid_ka_20161114pe1_v_l2
    } // group patch_ka_20161114_grid_ka_20161114pe1_v_l1
  } // group nz_linz_nzgd2000-ka20161114-grid06

group: nz_linz_nzgd2000-ka20161114-grid10 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake,  14 November 2016\nRefinement for horizontal difference between observations and model\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-11-14T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_hor_refinement {
    dimensions:
    	iNodeCount = 43 ;
    	jNodeCount = 40 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -38.625, 0., -0.125, 171.1, 0.15, 0. ;
    } // group patch_ka_20161114_grid_hor_refinement
  } // group nz_linz_nzgd2000-ka20161114-grid10

group: nz_linz_nzgd2000-ka20161114-grid11 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Kaikoura earthquake second refinement grid - horizontal" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_hor_refinement2 {
    dimensions:
    	iNodeCount = 214 ;
    	jNodeCount = 192 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.56, 0., -0.015, 171.5, 0.02, 0. ;
    } // group patch_ka_20161114_grid_hor_refinement2
  } // group nz_linz_nzgd2000-ka20161114-grid11

group: nz_linz_nzgd2000-ka20161114-grid12 {

  // group attributes:
  		:comment = "Kaikoura earthquake second refinement grid -vertical" ;
  		:gridParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "step" ;
  		:timeFunctions.0.eventDate = "2016-11-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-01-01T00:00:00Z" ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_vrt_refinement2 {
    dimensions:
    	iNodeCount = 216 ;
    	jNodeCount = 199 ;
    variables:
    	float displacement(iNodeCount, jNodeCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.395, 0., -0.015, 171.9, 0.02, 0. ;
    } // group patch_ka_20161114_grid_vrt_refinement2
  } // group nz_linz_nzgd2000-ka20161114-grid12

group: nz_linz_nzgd2000-ka20161114-grid07 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake months1-3 post-earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe3_h_l1_f {
    dimensions:
    	iNodeCount = 46 ;
    	jNodeCount = 40 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -38.875, 0., -0.125, 169.6, 0.15, 0. ;

    group: patch_ka_20161114_grid_ka_20161114pe3_h_l2_f {
      dimensions:
      	iNodeCount = 66 ;
      	jNodeCount = 60 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.0625, 0., -0.03125, 172.525, 0.0375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114pe3_h_l2_f
    } // group patch_ka_20161114_grid_ka_20161114pe3_h_l1_f
  } // group nz_linz_nzgd2000-ka20161114-grid07

group: nz_linz_nzgd2000-ka20161114-grid08 {
  dimensions:
  	displacementCount = 2 ;

  // group attributes:
  		:comment = "Event: Kaikoura earthquake months1-3 post-earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		string :gridParameters = "displacementEast", "displacementNorth" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe3_h_l2_r {
    dimensions:
    	iNodeCount = 67 ;
    	jNodeCount = 56 ;
    variables:
    	float displacement(iNodeCount, jNodeCount, displacementCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -41.28125, 0., -0.03125, 172.45, 0.0375, 0. ;

    group: patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_00 {
      dimensions:
      	iNodeCount = 88 ;
      	jNodeCount = 91 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -42., 0., -0.0078125, 172.91875, 0.009375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_00

    group: patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_01 {
      dimensions:
      	iNodeCount = 88 ;
      	jNodeCount = 122 ;
      variables:
      	float displacement(iNodeCount, jNodeCount, displacementCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -41.5546875, 0., -0.0078125, 173.734375, 0.009375, 0. ;
      } // group patch_ka_20161114_grid_ka_20161114pe3_h_l3_r_01
    } // group patch_ka_20161114_grid_ka_20161114pe3_h_l2_r
  } // group nz_linz_nzgd2000-ka20161114-grid08

group: nz_linz_nzgd2000-ka20161114-grid09 {

  // group attributes:
  		:comment = "Event: Kaikoura earthquake months1-3 post-earthquake,  14 November 2016\n Source model: Geodetic source model, based on GPS, InSAR, and LiDAR data; elastic half-space assumption; \n Version: Model 002, 23 June 2017\n" ;
  		:gridParameters = "displacementUp" ;
  		:timeFunctions.count = 1LL ;
  		:timeFunctions.0.functionType = "ramp" ;
  		:timeFunctions.0.startDate = "2016-12-14T00:00:00Z" ;
  		:timeFunctions.0.endDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.0.functionReferenceDate = "2017-02-14T00:00:00Z" ;
  		:timeFunctions.0.scaleFactor = 1. ;
  		:interpolationMethod = "bilinear" ;

  group: patch_ka_20161114_grid_ka_20161114pe3_v_l1 {
    dimensions:
    	iNodeCount = 31 ;
    	jNodeCount = 28 ;
    variables:
    	float displacement(iNodeCount, jNodeCount) ;
    		displacement:_Storage = "contiguous" ;
    		displacement:_Endianness = "little" ;

    // group attributes:
    		:affineCoeffs = -40.25, 0., -0.125, 171.4, 0.15, 0. ;

    group: patch_ka_20161114_grid_ka_20161114pe3_v_l2 {
      dimensions:
      	iNodeCount = 82 ;
      	jNodeCount = 76 ;
      variables:
      	float displacement(iNodeCount, jNodeCount) ;
      		displacement:_Storage = "contiguous" ;
      		displacement:_Endianness = "little" ;

      // group attributes:
      		:affineCoeffs = -40.65625, 0., -0.03125, 172.1875, 0.0375, 0. ;

      group: patch_ka_20161114_grid_ka_20161114pe3_v_l3_00 {
        dimensions:
        	iNodeCount = 92 ;
        	jNodeCount = 80 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -42.0703125, 0., -0.0078125, 172.825, 0.009375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114pe3_v_l3_00

      group: patch_ka_20161114_grid_ka_20161114pe3_v_l3_01 {
        dimensions:
        	iNodeCount = 92 ;
        	jNodeCount = 121 ;
        variables:
        	float displacement(iNodeCount, jNodeCount) ;
        		displacement:_Storage = "contiguous" ;
        		displacement:_Endianness = "little" ;

        // group attributes:
        		:affineCoeffs = -41.5859375, 0., -0.0078125, 173.678125, 0.009375, 0. ;
        } // group patch_ka_20161114_grid_ka_20161114pe3_v_l3_01
      } // group patch_ka_20161114_grid_ka_20161114pe3_v_l2
    } // group patch_ka_20161114_grid_ka_20161114pe3_v_l1
  } // group nz_linz_nzgd2000-ka20161114-grid09
}
